magic
tech sky130B
magscale 1 2
timestamp 1680599221
<< viali >>
rect 4905 33541 4939 33575
rect 7849 33541 7883 33575
rect 10793 33541 10827 33575
rect 14473 33541 14507 33575
rect 17049 33541 17083 33575
rect 19717 33541 19751 33575
rect 22661 33541 22695 33575
rect 25605 33541 25639 33575
rect 28549 33541 28583 33575
rect 31493 33541 31527 33575
rect 34253 33541 34287 33575
rect 8033 33337 8067 33371
rect 10977 33337 11011 33371
rect 14289 33337 14323 33371
rect 16865 33337 16899 33371
rect 19533 33337 19567 33371
rect 22477 33337 22511 33371
rect 25421 33337 25455 33371
rect 31309 33337 31343 33371
rect 34069 33337 34103 33371
rect 4997 33269 5031 33303
rect 28457 33269 28491 33303
rect 16589 32929 16623 32963
rect 20637 32929 20671 32963
rect 10241 32861 10275 32895
rect 16313 32861 16347 32895
rect 16497 32861 16531 32895
rect 20545 32861 20579 32895
rect 22477 32861 22511 32895
rect 15853 32793 15887 32827
rect 10149 32725 10183 32759
rect 20913 32725 20947 32759
rect 22385 32725 22419 32759
rect 12265 32521 12299 32555
rect 13461 32521 13495 32555
rect 17325 32521 17359 32555
rect 18061 32521 18095 32555
rect 20729 32521 20763 32555
rect 12081 32453 12115 32487
rect 13277 32453 13311 32487
rect 21189 32453 21223 32487
rect 22109 32453 22143 32487
rect 9873 32385 9907 32419
rect 10425 32385 10459 32419
rect 10517 32385 10551 32419
rect 17233 32385 17267 32419
rect 18061 32385 18095 32419
rect 18245 32385 18279 32419
rect 21097 32385 21131 32419
rect 22017 32385 22051 32419
rect 22201 32385 22235 32419
rect 23029 32385 23063 32419
rect 23213 32385 23247 32419
rect 24501 32385 24535 32419
rect 24685 32385 24719 32419
rect 27721 32385 27755 32419
rect 28089 32385 28123 32419
rect 30481 32385 30515 32419
rect 33333 32385 33367 32419
rect 10701 32317 10735 32351
rect 12357 32317 12391 32351
rect 13553 32317 13587 32351
rect 17417 32317 17451 32351
rect 21281 32317 21315 32351
rect 16865 32249 16899 32283
rect 22937 32249 22971 32283
rect 27169 32249 27203 32283
rect 9873 32181 9907 32215
rect 10609 32181 10643 32215
rect 11805 32181 11839 32215
rect 13001 32181 13035 32215
rect 24593 32181 24627 32215
rect 30297 32181 30331 32215
rect 33149 32181 33183 32215
rect 15761 31977 15795 32011
rect 18061 31977 18095 32011
rect 21281 31977 21315 32011
rect 23673 31977 23707 32011
rect 9321 31909 9355 31943
rect 11161 31909 11195 31943
rect 15945 31909 15979 31943
rect 18337 31909 18371 31943
rect 24593 31909 24627 31943
rect 8493 31841 8527 31875
rect 9781 31841 9815 31875
rect 9873 31841 9907 31875
rect 12633 31841 12667 31875
rect 13553 31841 13587 31875
rect 14381 31841 14415 31875
rect 16405 31841 16439 31875
rect 17141 31841 17175 31875
rect 19441 31841 19475 31875
rect 22017 31841 22051 31875
rect 22569 31841 22603 31875
rect 23029 31841 23063 31875
rect 25053 31841 25087 31875
rect 25145 31841 25179 31875
rect 8401 31773 8435 31807
rect 8585 31773 8619 31807
rect 9689 31773 9723 31807
rect 11437 31773 11471 31807
rect 11713 31773 11747 31807
rect 13461 31773 13495 31807
rect 14289 31773 14323 31807
rect 14473 31773 14507 31807
rect 17233 31773 17267 31807
rect 17325 31773 17359 31807
rect 18337 31773 18371 31807
rect 18521 31773 18555 31807
rect 20269 31773 20303 31807
rect 20453 31773 20487 31807
rect 21005 31773 21039 31807
rect 21281 31773 21315 31807
rect 22845 31773 22879 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 26433 31773 26467 31807
rect 26617 31773 26651 31807
rect 15577 31705 15611 31739
rect 16865 31705 16899 31739
rect 21097 31705 21131 31739
rect 11621 31637 11655 31671
rect 15777 31637 15811 31671
rect 23489 31637 23523 31671
rect 24961 31637 24995 31671
rect 9505 31433 9539 31467
rect 13553 31433 13587 31467
rect 16129 31433 16163 31467
rect 17049 31433 17083 31467
rect 17601 31433 17635 31467
rect 20846 31433 20880 31467
rect 24777 31433 24811 31467
rect 25881 31433 25915 31467
rect 28641 31433 28675 31467
rect 10701 31365 10735 31399
rect 16865 31365 16899 31399
rect 22201 31365 22235 31399
rect 27169 31365 27203 31399
rect 9137 31297 9171 31331
rect 10241 31297 10275 31331
rect 10333 31297 10367 31331
rect 13185 31297 13219 31331
rect 14105 31297 14139 31331
rect 14841 31297 14875 31331
rect 14933 31297 14967 31331
rect 16129 31297 16163 31331
rect 16313 31297 16347 31331
rect 17141 31297 17175 31331
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 20637 31297 20671 31331
rect 21097 31297 21131 31331
rect 22661 31297 22695 31331
rect 22753 31297 22787 31331
rect 23029 31297 23063 31331
rect 23305 31297 23339 31331
rect 23489 31297 23523 31331
rect 24225 31297 24259 31331
rect 24593 31297 24627 31331
rect 25237 31297 25271 31331
rect 25421 31297 25455 31331
rect 25605 31297 25639 31331
rect 25697 31297 25731 31331
rect 27353 31297 27387 31331
rect 27905 31297 27939 31331
rect 28579 31297 28613 31331
rect 9229 31229 9263 31263
rect 10425 31229 10459 31263
rect 13277 31229 13311 31263
rect 20545 31229 20579 31263
rect 29101 31229 29135 31263
rect 10885 31161 10919 31195
rect 25513 31161 25547 31195
rect 14289 31093 14323 31127
rect 16865 31093 16899 31127
rect 24593 31093 24627 31127
rect 28457 31093 28491 31127
rect 29009 31093 29043 31127
rect 9413 30889 9447 30923
rect 10057 30889 10091 30923
rect 10701 30889 10735 30923
rect 13553 30889 13587 30923
rect 17049 30889 17083 30923
rect 21005 30889 21039 30923
rect 22753 30889 22787 30923
rect 23121 30821 23155 30855
rect 27537 30821 27571 30855
rect 13461 30753 13495 30787
rect 15761 30753 15795 30787
rect 9321 30685 9355 30719
rect 9505 30685 9539 30719
rect 9965 30685 9999 30719
rect 10149 30685 10183 30719
rect 10609 30685 10643 30719
rect 10793 30685 10827 30719
rect 13645 30685 13679 30719
rect 13737 30685 13771 30719
rect 14565 30685 14599 30719
rect 14933 30685 14967 30719
rect 15485 30685 15519 30719
rect 15945 30685 15979 30719
rect 16129 30685 16163 30719
rect 16865 30685 16899 30719
rect 17049 30685 17083 30719
rect 20729 30685 20763 30719
rect 20821 30685 20855 30719
rect 22937 30685 22971 30719
rect 23213 30685 23247 30719
rect 25053 30685 25087 30719
rect 25605 30685 25639 30719
rect 26065 30685 26099 30719
rect 26249 30685 26283 30719
rect 27721 30685 27755 30719
rect 28089 30685 28123 30719
rect 28457 30685 28491 30719
rect 28917 30685 28951 30719
rect 26157 30617 26191 30651
rect 29745 30345 29779 30379
rect 28089 30277 28123 30311
rect 28549 30277 28583 30311
rect 14289 30209 14323 30243
rect 14933 30209 14967 30243
rect 19717 30209 19751 30243
rect 20269 30209 20303 30243
rect 21005 30209 21039 30243
rect 24685 30209 24719 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 25605 30209 25639 30243
rect 25881 30209 25915 30243
rect 26065 30209 26099 30243
rect 27353 30209 27387 30243
rect 27629 30209 27663 30243
rect 28733 30209 28767 30243
rect 29009 30209 29043 30243
rect 29193 30209 29227 30243
rect 29653 30209 29687 30243
rect 29837 30209 29871 30243
rect 27445 30141 27479 30175
rect 13461 30005 13495 30039
rect 20913 30005 20947 30039
rect 14841 29801 14875 29835
rect 25053 29801 25087 29835
rect 10425 29733 10459 29767
rect 27353 29733 27387 29767
rect 30021 29733 30055 29767
rect 20453 29665 20487 29699
rect 21557 29665 21591 29699
rect 27721 29665 27755 29699
rect 28825 29665 28859 29699
rect 9689 29597 9723 29631
rect 9965 29597 9999 29631
rect 10425 29597 10459 29631
rect 10517 29597 10551 29631
rect 13001 29597 13035 29631
rect 13185 29597 13219 29631
rect 14933 29597 14967 29631
rect 19625 29597 19659 29631
rect 20177 29597 20211 29631
rect 21005 29597 21039 29631
rect 21373 29597 21407 29631
rect 24777 29597 24811 29631
rect 24869 29597 24903 29631
rect 27537 29597 27571 29631
rect 27629 29597 27663 29631
rect 27813 29597 27847 29631
rect 28365 29597 28399 29631
rect 28549 29597 28583 29631
rect 28917 29597 28951 29631
rect 29745 29597 29779 29631
rect 29929 29597 29963 29631
rect 10701 29529 10735 29563
rect 15117 29529 15151 29563
rect 9505 29461 9539 29495
rect 9873 29461 9907 29495
rect 12817 29461 12851 29495
rect 19533 29461 19567 29495
rect 21373 29461 21407 29495
rect 14565 29257 14599 29291
rect 20177 29257 20211 29291
rect 22109 29257 22143 29291
rect 27905 29257 27939 29291
rect 28933 29257 28967 29291
rect 29101 29257 29135 29291
rect 15393 29189 15427 29223
rect 17693 29189 17727 29223
rect 25237 29189 25271 29223
rect 27261 29189 27295 29223
rect 28733 29189 28767 29223
rect 9045 29121 9079 29155
rect 9321 29121 9355 29155
rect 9505 29121 9539 29155
rect 11805 29121 11839 29155
rect 12541 29121 12575 29155
rect 12633 29121 12667 29155
rect 12909 29121 12943 29155
rect 13185 29121 13219 29155
rect 14749 29121 14783 29155
rect 15577 29121 15611 29155
rect 15761 29121 15795 29155
rect 19165 29121 19199 29155
rect 19533 29121 19567 29155
rect 20361 29121 20395 29155
rect 20453 29121 20487 29155
rect 20637 29121 20671 29155
rect 20729 29121 20763 29155
rect 21189 29121 21223 29155
rect 21373 29121 21407 29155
rect 22293 29121 22327 29155
rect 22569 29121 22603 29155
rect 22753 29121 22787 29155
rect 25329 29121 25363 29155
rect 25605 29121 25639 29155
rect 27169 29121 27203 29155
rect 27353 29121 27387 29155
rect 28089 29121 28123 29155
rect 14933 29053 14967 29087
rect 28273 29053 28307 29087
rect 21281 28985 21315 29019
rect 22385 28985 22419 29019
rect 22477 28985 22511 29019
rect 9413 28917 9447 28951
rect 11805 28917 11839 28951
rect 28917 28917 28951 28951
rect 21189 28713 21223 28747
rect 28825 28713 28859 28747
rect 15209 28645 15243 28679
rect 10977 28577 11011 28611
rect 11621 28577 11655 28611
rect 13185 28577 13219 28611
rect 13370 28577 13404 28611
rect 20177 28577 20211 28611
rect 26249 28577 26283 28611
rect 9321 28509 9355 28543
rect 9597 28509 9631 28543
rect 11345 28509 11379 28543
rect 12081 28509 12115 28543
rect 12357 28509 12391 28543
rect 13093 28509 13127 28543
rect 13277 28509 13311 28543
rect 14565 28509 14599 28543
rect 14933 28509 14967 28543
rect 15393 28509 15427 28543
rect 16313 28509 16347 28543
rect 19809 28509 19843 28543
rect 19993 28509 20027 28543
rect 20627 28509 20661 28543
rect 20717 28509 20751 28543
rect 20913 28509 20947 28543
rect 21005 28509 21039 28543
rect 22845 28509 22879 28543
rect 23397 28509 23431 28543
rect 28733 28509 28767 28543
rect 16681 28441 16715 28475
rect 9137 28373 9171 28407
rect 9505 28373 9539 28407
rect 12909 28373 12943 28407
rect 27261 28373 27295 28407
rect 8125 28169 8159 28203
rect 15393 28169 15427 28203
rect 22293 28169 22327 28203
rect 23213 28169 23247 28203
rect 15945 28101 15979 28135
rect 20637 28101 20671 28135
rect 23673 28101 23707 28135
rect 30297 28101 30331 28135
rect 7941 28033 7975 28067
rect 8217 28033 8251 28067
rect 9045 28033 9079 28067
rect 9689 28033 9723 28067
rect 9873 28033 9907 28067
rect 12173 28033 12207 28067
rect 12541 28033 12575 28067
rect 12909 28033 12943 28067
rect 13369 28033 13403 28067
rect 13829 28033 13863 28067
rect 14013 28033 14047 28067
rect 14197 28033 14231 28067
rect 15393 28033 15427 28067
rect 19257 28033 19291 28067
rect 19441 28033 19475 28067
rect 20269 28033 20303 28067
rect 20545 28033 20579 28067
rect 25053 28033 25087 28067
rect 25697 28033 25731 28067
rect 27261 28033 27295 28067
rect 27537 28033 27571 28067
rect 30113 28033 30147 28067
rect 30389 28033 30423 28067
rect 8769 27965 8803 27999
rect 8861 27965 8895 27999
rect 8953 27965 8987 27999
rect 12449 27965 12483 27999
rect 15301 27965 15335 27999
rect 19349 27965 19383 27999
rect 22753 27965 22787 27999
rect 25789 27965 25823 27999
rect 27169 27965 27203 27999
rect 22477 27897 22511 27931
rect 23397 27897 23431 27931
rect 24869 27897 24903 27931
rect 7757 27829 7791 27863
rect 9229 27829 9263 27863
rect 9781 27829 9815 27863
rect 29929 27829 29963 27863
rect 16865 27557 16899 27591
rect 25237 27557 25271 27591
rect 27905 27557 27939 27591
rect 9229 27489 9263 27523
rect 12817 27489 12851 27523
rect 28457 27489 28491 27523
rect 9321 27421 9355 27455
rect 9689 27421 9723 27455
rect 13185 27421 13219 27455
rect 13369 27421 13403 27455
rect 14933 27421 14967 27455
rect 15945 27421 15979 27455
rect 16037 27421 16071 27455
rect 16221 27421 16255 27455
rect 18245 27421 18279 27455
rect 22017 27421 22051 27455
rect 22293 27421 22327 27455
rect 25421 27421 25455 27455
rect 25697 27421 25731 27455
rect 26065 27421 26099 27455
rect 26341 27421 26375 27455
rect 26709 27421 26743 27455
rect 27445 27421 27479 27455
rect 27721 27421 27755 27455
rect 28365 27421 28399 27455
rect 28549 27421 28583 27455
rect 29837 27421 29871 27455
rect 10149 27353 10183 27387
rect 14381 27353 14415 27387
rect 16405 27353 16439 27387
rect 17978 27353 18012 27387
rect 30104 27353 30138 27387
rect 22109 27285 22143 27319
rect 22477 27285 22511 27319
rect 27537 27285 27571 27319
rect 31217 27285 31251 27319
rect 12081 27081 12115 27115
rect 19533 27081 19567 27115
rect 21189 27081 21223 27115
rect 31125 27081 31159 27115
rect 8309 27013 8343 27047
rect 15485 27013 15519 27047
rect 22661 27013 22695 27047
rect 27537 27013 27571 27047
rect 8217 26945 8251 26979
rect 8493 26945 8527 26979
rect 9229 26945 9263 26979
rect 11897 26945 11931 26979
rect 12173 26945 12207 26979
rect 13737 26945 13771 26979
rect 15669 26945 15703 26979
rect 15761 26945 15795 26979
rect 18245 26945 18279 26979
rect 21005 26945 21039 26979
rect 21281 26945 21315 26979
rect 22109 26945 22143 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 25881 26945 25915 26979
rect 27261 26945 27295 26979
rect 27445 26945 27479 26979
rect 30021 26945 30055 26979
rect 9045 26877 9079 26911
rect 9137 26877 9171 26911
rect 9321 26877 9355 26911
rect 26433 26877 26467 26911
rect 29745 26877 29779 26911
rect 8493 26809 8527 26843
rect 9505 26741 9539 26775
rect 11713 26741 11747 26775
rect 13645 26741 13679 26775
rect 20821 26741 20855 26775
rect 12357 26537 12391 26571
rect 13461 26537 13495 26571
rect 16681 26537 16715 26571
rect 25237 26537 25271 26571
rect 27077 26537 27111 26571
rect 32229 26537 32263 26571
rect 9413 26469 9447 26503
rect 13277 26469 13311 26503
rect 31309 26469 31343 26503
rect 11161 26401 11195 26435
rect 11713 26401 11747 26435
rect 12725 26401 12759 26435
rect 18061 26401 18095 26435
rect 25513 26401 25547 26435
rect 27721 26401 27755 26435
rect 11345 26333 11379 26367
rect 12633 26333 12667 26367
rect 19625 26333 19659 26367
rect 19809 26333 19843 26367
rect 19901 26333 19935 26367
rect 25421 26333 25455 26367
rect 25605 26333 25639 26367
rect 25697 26333 25731 26367
rect 25881 26333 25915 26367
rect 26525 26333 26559 26367
rect 26617 26333 26651 26367
rect 26801 26333 26835 26367
rect 26893 26333 26927 26367
rect 27537 26333 27571 26367
rect 32413 26333 32447 26367
rect 32689 26333 32723 26367
rect 9137 26265 9171 26299
rect 11621 26265 11655 26299
rect 13429 26265 13463 26299
rect 13645 26265 13679 26299
rect 17794 26265 17828 26299
rect 19441 26265 19475 26299
rect 22569 26265 22603 26299
rect 30021 26265 30055 26299
rect 32597 26265 32631 26299
rect 9597 26197 9631 26231
rect 21097 26197 21131 26231
rect 12265 25993 12299 26027
rect 16865 25993 16899 26027
rect 25605 25993 25639 26027
rect 27169 25993 27203 26027
rect 29929 25993 29963 26027
rect 10517 25925 10551 25959
rect 12357 25925 12391 25959
rect 12449 25925 12483 25959
rect 13093 25925 13127 25959
rect 13369 25925 13403 25959
rect 17233 25925 17267 25959
rect 21373 25925 21407 25959
rect 24593 25925 24627 25959
rect 25145 25925 25179 25959
rect 28641 25925 28675 25959
rect 32689 25925 32723 25959
rect 9505 25857 9539 25891
rect 9781 25857 9815 25891
rect 10425 25857 10459 25891
rect 10701 25857 10735 25891
rect 13277 25857 13311 25891
rect 13466 25857 13500 25891
rect 17049 25857 17083 25891
rect 17325 25857 17359 25891
rect 19625 25857 19659 25891
rect 20821 25857 20855 25891
rect 22017 25857 22051 25891
rect 22293 25857 22327 25891
rect 24501 25857 24535 25891
rect 24685 25857 24719 25891
rect 26525 25857 26559 25891
rect 27629 25857 27663 25891
rect 32505 25857 32539 25891
rect 32781 25857 32815 25891
rect 9597 25789 9631 25823
rect 12081 25789 12115 25823
rect 23489 25789 23523 25823
rect 26617 25789 26651 25823
rect 27353 25789 27387 25823
rect 27445 25789 27479 25823
rect 27537 25789 27571 25823
rect 9965 25721 9999 25755
rect 25421 25721 25455 25755
rect 10701 25653 10735 25687
rect 12633 25653 12667 25687
rect 13093 25653 13127 25687
rect 18337 25653 18371 25687
rect 32321 25653 32355 25687
rect 15393 25449 15427 25483
rect 19809 25449 19843 25483
rect 26065 25449 26099 25483
rect 26249 25449 26283 25483
rect 28273 25449 28307 25483
rect 16313 25381 16347 25415
rect 21189 25313 21223 25347
rect 26617 25313 26651 25347
rect 3433 25245 3467 25279
rect 4077 25245 4111 25279
rect 4261 25245 4295 25279
rect 6745 25245 6779 25279
rect 6929 25245 6963 25279
rect 12265 25245 12299 25279
rect 12541 25245 12575 25279
rect 12725 25245 12759 25279
rect 16037 25245 16071 25279
rect 16313 25245 16347 25279
rect 20922 25245 20956 25279
rect 24593 25245 24627 25279
rect 24869 25245 24903 25279
rect 27352 25245 27386 25279
rect 27445 25245 27479 25279
rect 28365 25245 28399 25279
rect 30113 25245 30147 25279
rect 3985 25177 4019 25211
rect 15377 25177 15411 25211
rect 15577 25177 15611 25211
rect 21649 25177 21683 25211
rect 26249 25177 26283 25211
rect 30380 25177 30414 25211
rect 3341 25109 3375 25143
rect 6745 25109 6779 25143
rect 12081 25109 12115 25143
rect 15209 25109 15243 25143
rect 16129 25109 16163 25143
rect 22937 25109 22971 25143
rect 27077 25109 27111 25143
rect 31493 25109 31527 25143
rect 31493 24905 31527 24939
rect 5273 24837 5307 24871
rect 21097 24837 21131 24871
rect 21465 24837 21499 24871
rect 23673 24837 23707 24871
rect 28641 24837 28675 24871
rect 28825 24837 28859 24871
rect 2329 24769 2363 24803
rect 6929 24769 6963 24803
rect 14841 24769 14875 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 15945 24769 15979 24803
rect 16129 24769 16163 24803
rect 18153 24769 18187 24803
rect 21005 24769 21039 24803
rect 21281 24769 21315 24803
rect 25237 24769 25271 24803
rect 25329 24769 25363 24803
rect 26157 24769 26191 24803
rect 29101 24769 29135 24803
rect 30380 24769 30414 24803
rect 2605 24701 2639 24735
rect 4721 24701 4755 24735
rect 7941 24701 7975 24735
rect 15301 24701 15335 24735
rect 17877 24701 17911 24735
rect 19349 24701 19383 24735
rect 22017 24701 22051 24735
rect 22293 24701 22327 24735
rect 26433 24701 26467 24735
rect 30113 24701 30147 24735
rect 3893 24633 3927 24667
rect 25145 24633 25179 24667
rect 16129 24565 16163 24599
rect 25973 24565 26007 24599
rect 26341 24565 26375 24599
rect 28825 24565 28859 24599
rect 2789 24361 2823 24395
rect 6837 24361 6871 24395
rect 30573 24361 30607 24395
rect 2329 24293 2363 24327
rect 5273 24293 5307 24327
rect 22845 24293 22879 24327
rect 4169 24225 4203 24259
rect 4353 24225 4387 24259
rect 5181 24225 5215 24259
rect 21005 24225 21039 24259
rect 2053 24157 2087 24191
rect 2973 24157 3007 24191
rect 3065 24157 3099 24191
rect 4445 24157 4479 24191
rect 4537 24157 4571 24191
rect 4629 24157 4663 24191
rect 5549 24157 5583 24191
rect 5733 24157 5767 24191
rect 7573 24157 7607 24191
rect 8493 24157 8527 24191
rect 11897 24157 11931 24191
rect 12081 24157 12115 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 14749 24157 14783 24191
rect 14841 24157 14875 24191
rect 15669 24157 15703 24191
rect 15853 24157 15887 24191
rect 17049 24157 17083 24191
rect 17233 24157 17267 24191
rect 17923 24157 17957 24191
rect 18153 24157 18187 24191
rect 20729 24157 20763 24191
rect 20821 24157 20855 24191
rect 21465 24157 21499 24191
rect 23489 24157 23523 24191
rect 23765 24157 23799 24191
rect 25237 24157 25271 24191
rect 25421 24157 25455 24191
rect 30757 24157 30791 24191
rect 31033 24157 31067 24191
rect 2329 24089 2363 24123
rect 3341 24089 3375 24123
rect 3433 24089 3467 24123
rect 18061 24089 18095 24123
rect 21732 24089 21766 24123
rect 23305 24089 23339 24123
rect 2145 24021 2179 24055
rect 12081 24021 12115 24055
rect 14289 24021 14323 24055
rect 15485 24021 15519 24055
rect 17141 24021 17175 24055
rect 17693 24021 17727 24055
rect 23673 24021 23707 24055
rect 25329 24021 25363 24055
rect 30941 24021 30975 24055
rect 5089 23817 5123 23851
rect 14933 23817 14967 23851
rect 15117 23817 15151 23851
rect 15945 23817 15979 23851
rect 30113 23817 30147 23851
rect 10241 23749 10275 23783
rect 19993 23749 20027 23783
rect 22293 23749 22327 23783
rect 28641 23749 28675 23783
rect 2973 23681 3007 23715
rect 3709 23681 3743 23715
rect 5365 23681 5399 23715
rect 5549 23681 5583 23715
rect 9229 23681 9263 23715
rect 9873 23681 9907 23715
rect 10057 23681 10091 23715
rect 12909 23681 12943 23715
rect 13277 23681 13311 23715
rect 14381 23681 14415 23715
rect 16129 23681 16163 23715
rect 16313 23681 16347 23715
rect 20453 23681 20487 23715
rect 20637 23681 20671 23715
rect 22661 23681 22695 23715
rect 25513 23681 25547 23715
rect 4629 23613 4663 23647
rect 5273 23613 5307 23647
rect 5457 23613 5491 23647
rect 6837 23613 6871 23647
rect 7113 23613 7147 23647
rect 9045 23613 9079 23647
rect 9413 23613 9447 23647
rect 12265 23613 12299 23647
rect 13001 23613 13035 23647
rect 13185 23613 13219 23647
rect 14841 23613 14875 23647
rect 15209 23613 15243 23647
rect 15301 23613 15335 23647
rect 20821 23613 20855 23647
rect 14289 23545 14323 23579
rect 18705 23545 18739 23579
rect 8401 23477 8435 23511
rect 15485 23477 15519 23511
rect 25421 23477 25455 23511
rect 3249 23273 3283 23307
rect 3341 23273 3375 23307
rect 4169 23273 4203 23307
rect 6929 23273 6963 23307
rect 18705 23273 18739 23307
rect 21925 23273 21959 23307
rect 9137 23205 9171 23239
rect 15577 23205 15611 23239
rect 16129 23205 16163 23239
rect 19717 23205 19751 23239
rect 3433 23137 3467 23171
rect 8309 23137 8343 23171
rect 8585 23137 8619 23171
rect 15209 23137 15243 23171
rect 15301 23137 15335 23171
rect 16497 23137 16531 23171
rect 17325 23137 17359 23171
rect 24961 23137 24995 23171
rect 25329 23137 25363 23171
rect 32689 23137 32723 23171
rect 33149 23137 33183 23171
rect 3157 23069 3191 23103
rect 7113 23069 7147 23103
rect 7415 23069 7449 23103
rect 7573 23069 7607 23103
rect 8125 23069 8159 23103
rect 8217 23069 8251 23103
rect 8401 23069 8435 23103
rect 9321 23069 9355 23103
rect 9413 23069 9447 23103
rect 12081 23069 12115 23103
rect 12541 23069 12575 23103
rect 15117 23069 15151 23103
rect 15393 23069 15427 23103
rect 17592 23069 17626 23103
rect 19441 23069 19475 23103
rect 19717 23069 19751 23103
rect 20637 23069 20671 23103
rect 24869 23069 24903 23103
rect 27537 23069 27571 23103
rect 27997 23069 28031 23103
rect 28273 23069 28307 23103
rect 31769 23069 31803 23103
rect 32045 23069 32079 23103
rect 32781 23069 32815 23103
rect 33609 23069 33643 23103
rect 33793 23069 33827 23103
rect 4353 23001 4387 23035
rect 7205 23001 7239 23035
rect 7297 23001 7331 23035
rect 9137 23001 9171 23035
rect 11805 23001 11839 23035
rect 13277 23001 13311 23035
rect 27813 23001 27847 23035
rect 3985 22933 4019 22967
rect 4153 22933 4187 22967
rect 10333 22933 10367 22967
rect 16037 22933 16071 22967
rect 24685 22933 24719 22967
rect 25053 22933 25087 22967
rect 25237 22933 25271 22967
rect 31033 22933 31067 22967
rect 33701 22933 33735 22967
rect 7205 22729 7239 22763
rect 32413 22729 32447 22763
rect 8125 22661 8159 22695
rect 8309 22661 8343 22695
rect 8493 22661 8527 22695
rect 9689 22661 9723 22695
rect 12541 22661 12575 22695
rect 14381 22661 14415 22695
rect 23765 22661 23799 22695
rect 25237 22661 25271 22695
rect 33057 22661 33091 22695
rect 33517 22661 33551 22695
rect 4445 22593 4479 22627
rect 7389 22593 7423 22627
rect 7573 22593 7607 22627
rect 7665 22593 7699 22627
rect 9413 22593 9447 22627
rect 9597 22593 9631 22627
rect 10333 22593 10367 22627
rect 11713 22593 11747 22627
rect 11897 22593 11931 22627
rect 12909 22593 12943 22627
rect 13277 22593 13311 22627
rect 13369 22593 13403 22627
rect 13645 22593 13679 22627
rect 13921 22593 13955 22627
rect 14657 22593 14691 22627
rect 15301 22593 15335 22627
rect 15485 22593 15519 22627
rect 15577 22593 15611 22627
rect 17325 22593 17359 22627
rect 17509 22593 17543 22627
rect 18153 22593 18187 22627
rect 18613 22593 18647 22627
rect 19993 22593 20027 22627
rect 20158 22593 20192 22627
rect 20269 22593 20303 22627
rect 20361 22593 20395 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 23673 22593 23707 22627
rect 24869 22593 24903 22627
rect 27997 22593 28031 22627
rect 28365 22593 28399 22627
rect 29929 22593 29963 22627
rect 31033 22593 31067 22627
rect 31218 22593 31252 22627
rect 32689 22593 32723 22627
rect 33701 22593 33735 22627
rect 4997 22525 5031 22559
rect 10977 22525 11011 22559
rect 14381 22525 14415 22559
rect 18245 22525 18279 22559
rect 24777 22525 24811 22559
rect 25145 22525 25179 22559
rect 29745 22525 29779 22559
rect 31125 22525 31159 22559
rect 31310 22525 31344 22559
rect 32551 22525 32585 22559
rect 32965 22525 32999 22559
rect 17417 22457 17451 22491
rect 22017 22457 22051 22491
rect 30113 22457 30147 22491
rect 11805 22389 11839 22423
rect 14565 22389 14599 22423
rect 15117 22389 15151 22423
rect 17969 22389 18003 22423
rect 19809 22389 19843 22423
rect 24593 22389 24627 22423
rect 27353 22389 27387 22423
rect 30849 22389 30883 22423
rect 33793 22389 33827 22423
rect 10241 22185 10275 22219
rect 11725 22185 11759 22219
rect 23029 22185 23063 22219
rect 23213 22185 23247 22219
rect 33517 22185 33551 22219
rect 12821 22117 12855 22151
rect 11989 22049 12023 22083
rect 17785 22049 17819 22083
rect 24777 22049 24811 22083
rect 24869 22049 24903 22083
rect 25053 22049 25087 22083
rect 26985 22049 27019 22083
rect 30205 22049 30239 22083
rect 33149 22049 33183 22083
rect 7205 21981 7239 22015
rect 8585 21981 8619 22015
rect 12725 21981 12759 22015
rect 12909 21981 12943 22015
rect 13001 21981 13035 22015
rect 17969 21981 18003 22015
rect 18337 21981 18371 22015
rect 19809 21981 19843 22015
rect 20821 21981 20855 22015
rect 23213 21981 23247 22015
rect 23397 21981 23431 22015
rect 24961 21981 24995 22015
rect 26065 21981 26099 22015
rect 26249 21981 26283 22015
rect 27077 21981 27111 22015
rect 27813 21981 27847 22015
rect 28641 21981 28675 22015
rect 30113 21981 30147 22015
rect 31033 21981 31067 22015
rect 31401 21981 31435 22015
rect 31585 21981 31619 22015
rect 32045 21981 32079 22015
rect 32413 21981 32447 22015
rect 32597 21981 32631 22015
rect 33333 21981 33367 22015
rect 20177 21913 20211 21947
rect 26157 21913 26191 21947
rect 28273 21913 28307 21947
rect 28457 21913 28491 21947
rect 31125 21913 31159 21947
rect 32137 21913 32171 21947
rect 7205 21845 7239 21879
rect 8493 21845 8527 21879
rect 12541 21845 12575 21879
rect 18245 21845 18279 21879
rect 22293 21845 22327 21879
rect 25237 21845 25271 21879
rect 27721 21845 27755 21879
rect 29745 21845 29779 21879
rect 27169 21641 27203 21675
rect 30297 21641 30331 21675
rect 31677 21641 31711 21675
rect 11713 21573 11747 21607
rect 30481 21573 30515 21607
rect 2881 21505 2915 21539
rect 3801 21505 3835 21539
rect 4077 21505 4111 21539
rect 11805 21505 11839 21539
rect 12081 21505 12115 21539
rect 14473 21505 14507 21539
rect 14565 21505 14599 21539
rect 15301 21505 15335 21539
rect 15485 21505 15519 21539
rect 19441 21505 19475 21539
rect 19809 21505 19843 21539
rect 20545 21505 20579 21539
rect 20637 21505 20671 21539
rect 22017 21505 22051 21539
rect 22293 21505 22327 21539
rect 27537 21505 27571 21539
rect 28181 21505 28215 21539
rect 28365 21505 28399 21539
rect 30205 21505 30239 21539
rect 31493 21505 31527 21539
rect 31677 21505 31711 21539
rect 2973 21437 3007 21471
rect 3157 21437 3191 21471
rect 19533 21437 19567 21471
rect 22385 21437 22419 21471
rect 23213 21437 23247 21471
rect 23489 21437 23523 21471
rect 27629 21437 27663 21471
rect 3893 21369 3927 21403
rect 3985 21369 4019 21403
rect 24777 21369 24811 21403
rect 3065 21301 3099 21335
rect 3617 21301 3651 21335
rect 15485 21301 15519 21335
rect 28365 21301 28399 21335
rect 30481 21301 30515 21335
rect 13461 21097 13495 21131
rect 14657 21097 14691 21131
rect 16129 21097 16163 21131
rect 21281 21097 21315 21131
rect 23581 21097 23615 21131
rect 32413 21097 32447 21131
rect 19533 21029 19567 21063
rect 33149 21029 33183 21063
rect 7389 20961 7423 20995
rect 19717 20961 19751 20995
rect 20085 20961 20119 20995
rect 20177 20961 20211 20995
rect 31309 20961 31343 20995
rect 3249 20893 3283 20927
rect 3433 20893 3467 20927
rect 7573 20893 7607 20927
rect 7665 20893 7699 20927
rect 10425 20893 10459 20927
rect 10701 20893 10735 20927
rect 13553 20893 13587 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 17417 20893 17451 20927
rect 19809 20893 19843 20927
rect 22569 20893 22603 20927
rect 23765 20893 23799 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 24796 20893 24830 20927
rect 25053 20893 25087 20927
rect 31584 20893 31618 20927
rect 31677 20893 31711 20927
rect 32229 20893 32263 20927
rect 32505 20893 32539 20927
rect 32965 20893 32999 20927
rect 33149 20893 33183 20927
rect 24593 20825 24627 20859
rect 3341 20757 3375 20791
rect 7389 20757 7423 20791
rect 10241 20757 10275 20791
rect 10609 20757 10643 20791
rect 14381 20757 14415 20791
rect 24961 20757 24995 20791
rect 7849 20553 7883 20587
rect 8401 20553 8435 20587
rect 19165 20553 19199 20587
rect 21097 20553 21131 20587
rect 31585 20553 31619 20587
rect 32597 20553 32631 20587
rect 3617 20485 3651 20519
rect 7481 20485 7515 20519
rect 20821 20485 20855 20519
rect 23213 20485 23247 20519
rect 3157 20417 3191 20451
rect 3249 20417 3283 20451
rect 4445 20417 4479 20451
rect 7389 20417 7423 20451
rect 7665 20417 7699 20451
rect 8309 20417 8343 20451
rect 8493 20417 8527 20451
rect 8585 20417 8619 20451
rect 11069 20417 11103 20451
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 15117 20417 15151 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 18337 20417 18371 20451
rect 18521 20417 18555 20451
rect 18613 20417 18647 20451
rect 19073 20417 19107 20451
rect 19349 20417 19383 20451
rect 20545 20417 20579 20451
rect 20729 20417 20763 20451
rect 20959 20417 20993 20451
rect 27997 20417 28031 20451
rect 31585 20417 31619 20451
rect 31769 20417 31803 20451
rect 32781 20417 32815 20451
rect 33057 20417 33091 20451
rect 3525 20349 3559 20383
rect 4077 20349 4111 20383
rect 4353 20349 4387 20383
rect 10333 20349 10367 20383
rect 12817 20349 12851 20383
rect 14657 20349 14691 20383
rect 27905 20349 27939 20383
rect 27629 20281 27663 20315
rect 32965 20281 32999 20315
rect 2973 20213 3007 20247
rect 15853 20213 15887 20247
rect 18153 20213 18187 20247
rect 19533 20213 19567 20247
rect 24501 20213 24535 20247
rect 27997 20213 28031 20247
rect 3985 20009 4019 20043
rect 7573 20009 7607 20043
rect 14473 20009 14507 20043
rect 18797 20009 18831 20043
rect 20085 20009 20119 20043
rect 7113 19941 7147 19975
rect 7757 19941 7791 19975
rect 9137 19941 9171 19975
rect 13645 19941 13679 19975
rect 32321 19941 32355 19975
rect 2421 19873 2455 19907
rect 3249 19873 3283 19907
rect 5161 19873 5195 19907
rect 10517 19873 10551 19907
rect 11897 19873 11931 19907
rect 22569 19873 22603 19907
rect 1685 19805 1719 19839
rect 1869 19805 1903 19839
rect 3157 19805 3191 19839
rect 4169 19805 4203 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 5365 19805 5399 19839
rect 6837 19805 6871 19839
rect 6929 19805 6963 19839
rect 7113 19805 7147 19839
rect 8033 19805 8067 19839
rect 9413 19805 9447 19839
rect 10425 19805 10459 19839
rect 10793 19805 10827 19839
rect 11069 19805 11103 19839
rect 11713 19805 11747 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 14381 19805 14415 19839
rect 15117 19805 15151 19839
rect 16313 19805 16347 19839
rect 18521 19805 18555 19839
rect 19441 19805 19475 19839
rect 19534 19805 19568 19839
rect 19717 19805 19751 19839
rect 19906 19805 19940 19839
rect 31953 19805 31987 19839
rect 32137 19805 32171 19839
rect 32413 19805 32447 19839
rect 32597 19805 32631 19839
rect 1777 19737 1811 19771
rect 4261 19737 4295 19771
rect 4353 19737 4387 19771
rect 5089 19737 5123 19771
rect 5273 19737 5307 19771
rect 9137 19737 9171 19771
rect 9321 19737 9355 19771
rect 15669 19737 15703 19771
rect 16865 19737 16899 19771
rect 19809 19737 19843 19771
rect 20821 19737 20855 19771
rect 11529 19669 11563 19703
rect 4445 19465 4479 19499
rect 16313 19465 16347 19499
rect 17233 19465 17267 19499
rect 20361 19465 20395 19499
rect 32505 19465 32539 19499
rect 32689 19465 32723 19499
rect 32873 19465 32907 19499
rect 2780 19397 2814 19431
rect 24777 19397 24811 19431
rect 28365 19397 28399 19431
rect 32321 19397 32355 19431
rect 2513 19329 2547 19363
rect 4629 19329 4663 19363
rect 7113 19329 7147 19363
rect 7380 19329 7414 19363
rect 9045 19329 9079 19363
rect 9229 19329 9263 19363
rect 10793 19329 10827 19363
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 15200 19329 15234 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17325 19329 17359 19363
rect 18981 19329 19015 19363
rect 19237 19329 19271 19363
rect 23121 19329 23155 19363
rect 27261 19329 27295 19363
rect 27445 19329 27479 19363
rect 29009 19329 29043 19363
rect 29377 19329 29411 19363
rect 31217 19329 31251 19363
rect 31401 19329 31435 19363
rect 32597 19329 32631 19363
rect 4813 19261 4847 19295
rect 10517 19261 10551 19295
rect 14933 19261 14967 19295
rect 23397 19261 23431 19295
rect 28825 19261 28859 19295
rect 29285 19261 29319 19295
rect 31125 19261 31159 19295
rect 3893 19125 3927 19159
rect 8493 19125 8527 19159
rect 9137 19125 9171 19159
rect 10241 19125 10275 19159
rect 10701 19125 10735 19159
rect 27353 19125 27387 19159
rect 7665 18921 7699 18955
rect 14565 18921 14599 18955
rect 16681 18921 16715 18955
rect 18705 18921 18739 18955
rect 20821 18921 20855 18955
rect 25881 18921 25915 18955
rect 33149 18921 33183 18955
rect 3157 18853 3191 18887
rect 7849 18785 7883 18819
rect 7941 18785 7975 18819
rect 8217 18785 8251 18819
rect 12357 18785 12391 18819
rect 26065 18785 26099 18819
rect 26157 18785 26191 18819
rect 31861 18785 31895 18819
rect 3341 18717 3375 18751
rect 3433 18717 3467 18751
rect 8309 18717 8343 18751
rect 10425 18717 10459 18751
rect 10517 18717 10551 18751
rect 11989 18717 12023 18751
rect 12265 18717 12299 18751
rect 15301 18717 15335 18751
rect 19441 18717 19475 18751
rect 23765 18717 23799 18751
rect 24041 18717 24075 18751
rect 24777 18717 24811 18751
rect 25053 18717 25087 18751
rect 26249 18717 26283 18751
rect 26341 18717 26375 18751
rect 27721 18717 27755 18751
rect 27905 18717 27939 18751
rect 28549 18717 28583 18751
rect 28825 18717 28859 18751
rect 29009 18717 29043 18751
rect 29837 18717 29871 18751
rect 30113 18717 30147 18751
rect 32045 18717 32079 18751
rect 32229 18717 32263 18751
rect 32689 18717 32723 18751
rect 32781 18717 32815 18751
rect 32965 18717 32999 18751
rect 3157 18649 3191 18683
rect 14381 18649 14415 18683
rect 14565 18649 14599 18683
rect 15568 18649 15602 18683
rect 18889 18649 18923 18683
rect 19708 18649 19742 18683
rect 27353 18649 27387 18683
rect 29745 18649 29779 18683
rect 8033 18581 8067 18615
rect 14749 18581 14783 18615
rect 18521 18581 18555 18615
rect 18705 18581 18739 18615
rect 23581 18581 23615 18615
rect 23949 18581 23983 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 28365 18581 28399 18615
rect 8217 18377 8251 18411
rect 15761 18377 15795 18411
rect 16129 18377 16163 18411
rect 24777 18377 24811 18411
rect 25697 18377 25731 18411
rect 32781 18377 32815 18411
rect 6837 18309 6871 18343
rect 14749 18309 14783 18343
rect 19257 18309 19291 18343
rect 8033 18241 8067 18275
rect 8217 18241 8251 18275
rect 10333 18241 10367 18275
rect 12265 18241 12299 18275
rect 12449 18241 12483 18275
rect 13001 18241 13035 18275
rect 15945 18241 15979 18275
rect 16221 18241 16255 18275
rect 23489 18241 23523 18275
rect 25329 18241 25363 18275
rect 25513 18241 25547 18275
rect 27905 18241 27939 18275
rect 28825 18241 28859 18275
rect 29101 18241 29135 18275
rect 29377 18241 29411 18275
rect 29745 18241 29779 18275
rect 32505 18241 32539 18275
rect 6745 18173 6779 18207
rect 6929 18173 6963 18207
rect 12173 18173 12207 18207
rect 23213 18173 23247 18207
rect 27537 18173 27571 18207
rect 27997 18173 28031 18207
rect 32321 18173 32355 18207
rect 32873 18173 32907 18207
rect 34345 18173 34379 18207
rect 7297 18105 7331 18139
rect 28641 18105 28675 18139
rect 10241 18037 10275 18071
rect 20545 18037 20579 18071
rect 25329 18037 25363 18071
rect 6469 17833 6503 17867
rect 27997 17833 28031 17867
rect 32689 17833 32723 17867
rect 3433 17765 3467 17799
rect 21557 17765 21591 17799
rect 13093 17697 13127 17731
rect 27629 17697 27663 17731
rect 28457 17697 28491 17731
rect 33609 17697 33643 17731
rect 3249 17629 3283 17663
rect 6377 17629 6411 17663
rect 6561 17629 6595 17663
rect 15209 17629 15243 17663
rect 17601 17629 17635 17663
rect 17877 17629 17911 17663
rect 18429 17629 18463 17663
rect 18705 17629 18739 17663
rect 19441 17629 19475 17663
rect 21373 17629 21407 17663
rect 24777 17629 24811 17663
rect 25053 17629 25087 17663
rect 27537 17629 27571 17663
rect 27721 17629 27755 17663
rect 27813 17629 27847 17663
rect 28641 17629 28675 17663
rect 28917 17629 28951 17663
rect 30757 17629 30791 17663
rect 30941 17629 30975 17663
rect 31769 17629 31803 17663
rect 31953 17629 31987 17663
rect 32597 17629 32631 17663
rect 33241 17629 33275 17663
rect 33425 17629 33459 17663
rect 2881 17561 2915 17595
rect 12817 17561 12851 17595
rect 18889 17561 18923 17595
rect 19686 17561 19720 17595
rect 31125 17561 31159 17595
rect 31861 17561 31895 17595
rect 32413 17561 32447 17595
rect 3065 17493 3099 17527
rect 3157 17493 3191 17527
rect 11345 17493 11379 17527
rect 16497 17493 16531 17527
rect 17417 17493 17451 17527
rect 17785 17493 17819 17527
rect 18521 17493 18555 17527
rect 20821 17493 20855 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 28825 17493 28859 17527
rect 4445 17289 4479 17323
rect 19533 17289 19567 17323
rect 25697 17289 25731 17323
rect 28549 17289 28583 17323
rect 30757 17289 30791 17323
rect 30941 17289 30975 17323
rect 32521 17289 32555 17323
rect 32689 17289 32723 17323
rect 33241 17289 33275 17323
rect 2973 17221 3007 17255
rect 9597 17221 9631 17255
rect 13277 17221 13311 17255
rect 16865 17221 16899 17255
rect 18245 17221 18279 17255
rect 20821 17221 20855 17255
rect 23388 17221 23422 17255
rect 25421 17221 25455 17255
rect 28641 17221 28675 17255
rect 29837 17221 29871 17255
rect 30849 17221 30883 17255
rect 31493 17221 31527 17255
rect 32321 17221 32355 17255
rect 6745 17153 6779 17187
rect 7113 17153 7147 17187
rect 7573 17153 7607 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 9873 17153 9907 17187
rect 16221 17153 16255 17187
rect 17693 17153 17727 17187
rect 20637 17153 20671 17187
rect 20913 17153 20947 17187
rect 25053 17153 25087 17187
rect 25146 17153 25180 17187
rect 25329 17153 25363 17187
rect 25559 17153 25593 17187
rect 26157 17153 26191 17187
rect 28549 17153 28583 17187
rect 28825 17153 28859 17187
rect 29745 17153 29779 17187
rect 29929 17153 29963 17187
rect 30481 17153 30515 17187
rect 30625 17153 30659 17187
rect 31677 17153 31711 17187
rect 31769 17153 31803 17187
rect 33149 17153 33183 17187
rect 33333 17153 33367 17187
rect 2697 17085 2731 17119
rect 6653 17085 6687 17119
rect 9781 17085 9815 17119
rect 13553 17085 13587 17119
rect 15945 17085 15979 17119
rect 23121 17085 23155 17119
rect 26433 17085 26467 17119
rect 31493 17017 31527 17051
rect 8217 16949 8251 16983
rect 9689 16949 9723 16983
rect 10057 16949 10091 16983
rect 11805 16949 11839 16983
rect 20453 16949 20487 16983
rect 24501 16949 24535 16983
rect 32505 16949 32539 16983
rect 3249 16745 3283 16779
rect 4261 16745 4295 16779
rect 6837 16745 6871 16779
rect 12265 16745 12299 16779
rect 21373 16745 21407 16779
rect 31217 16745 31251 16779
rect 32229 16745 32263 16779
rect 3065 16677 3099 16711
rect 5917 16677 5951 16711
rect 7205 16677 7239 16711
rect 9781 16677 9815 16711
rect 14841 16677 14875 16711
rect 7113 16609 7147 16643
rect 7334 16609 7368 16643
rect 15301 16609 15335 16643
rect 17509 16609 17543 16643
rect 29745 16609 29779 16643
rect 32597 16609 32631 16643
rect 4077 16541 4111 16575
rect 4261 16541 4295 16575
rect 9689 16541 9723 16575
rect 9965 16541 9999 16575
rect 10057 16541 10091 16575
rect 12173 16541 12207 16575
rect 12357 16541 12391 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 15568 16541 15602 16575
rect 17233 16541 17267 16575
rect 19441 16541 19475 16575
rect 19708 16541 19742 16575
rect 21557 16541 21591 16575
rect 24593 16541 24627 16575
rect 26433 16541 26467 16575
rect 29929 16541 29963 16575
rect 31217 16541 31251 16575
rect 31493 16541 31527 16575
rect 31621 16541 31655 16575
rect 32413 16541 32447 16575
rect 3433 16473 3467 16507
rect 5549 16473 5583 16507
rect 7481 16473 7515 16507
rect 24860 16473 24894 16507
rect 26709 16473 26743 16507
rect 30021 16473 30055 16507
rect 31401 16473 31435 16507
rect 3233 16405 3267 16439
rect 6009 16405 6043 16439
rect 10241 16405 10275 16439
rect 14473 16405 14507 16439
rect 16681 16405 16715 16439
rect 20821 16405 20855 16439
rect 25973 16405 26007 16439
rect 30113 16405 30147 16439
rect 30297 16405 30331 16439
rect 6745 16201 6779 16235
rect 10977 16201 11011 16235
rect 13461 16201 13495 16235
rect 19533 16201 19567 16235
rect 20453 16201 20487 16235
rect 22661 16201 22695 16235
rect 26065 16201 26099 16235
rect 33701 16201 33735 16235
rect 5733 16133 5767 16167
rect 8861 16133 8895 16167
rect 14289 16133 14323 16167
rect 15200 16133 15234 16167
rect 18245 16133 18279 16167
rect 20729 16133 20763 16167
rect 26433 16133 26467 16167
rect 28641 16133 28675 16167
rect 5457 16065 5491 16099
rect 5549 16065 5583 16099
rect 6561 16065 6595 16099
rect 6745 16065 6779 16099
rect 7389 16065 7423 16099
rect 8769 16065 8803 16099
rect 10425 16065 10459 16099
rect 10977 16065 11011 16099
rect 11161 16065 11195 16099
rect 13277 16065 13311 16099
rect 14013 16065 14047 16099
rect 17417 16065 17451 16099
rect 17693 16065 17727 16099
rect 20591 16065 20625 16099
rect 20821 16065 20855 16099
rect 20949 16065 20983 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 22110 16065 22144 16099
rect 22293 16065 22327 16099
rect 22385 16065 22419 16099
rect 22523 16065 22557 16099
rect 25145 16065 25179 16099
rect 26249 16065 26283 16099
rect 26525 16065 26559 16099
rect 28549 16065 28583 16099
rect 28733 16065 28767 16099
rect 28917 16065 28951 16099
rect 29561 16065 29595 16099
rect 32588 16065 32622 16099
rect 7665 15997 7699 16031
rect 14933 15997 14967 16031
rect 17785 15997 17819 16031
rect 32321 15997 32355 16031
rect 7941 15929 7975 15963
rect 7757 15861 7791 15895
rect 16313 15861 16347 15895
rect 23857 15861 23891 15895
rect 28365 15861 28399 15895
rect 29469 15861 29503 15895
rect 5273 15657 5307 15691
rect 10885 15657 10919 15691
rect 26433 15657 26467 15691
rect 31677 15657 31711 15691
rect 33885 15657 33919 15691
rect 2881 15589 2915 15623
rect 13645 15589 13679 15623
rect 27997 15589 28031 15623
rect 14933 15521 14967 15555
rect 16129 15521 16163 15555
rect 18245 15521 18279 15555
rect 22569 15521 22603 15555
rect 28181 15521 28215 15555
rect 28365 15521 28399 15555
rect 2697 15453 2731 15487
rect 2973 15453 3007 15487
rect 6101 15453 6135 15487
rect 6285 15453 6319 15487
rect 6745 15453 6779 15487
rect 12633 15453 12667 15487
rect 12725 15453 12759 15487
rect 13369 15453 13403 15487
rect 13645 15453 13679 15487
rect 15117 15453 15151 15487
rect 15301 15453 15335 15487
rect 16037 15453 16071 15487
rect 16313 15453 16347 15487
rect 17877 15453 17911 15487
rect 20821 15453 20855 15487
rect 23213 15453 23247 15487
rect 23489 15453 23523 15487
rect 28273 15453 28307 15487
rect 28457 15453 28491 15487
rect 33425 15453 33459 15487
rect 33701 15453 33735 15487
rect 5457 15385 5491 15419
rect 6193 15385 6227 15419
rect 12173 15385 12207 15419
rect 17693 15385 17727 15419
rect 23397 15385 23431 15419
rect 25145 15385 25179 15419
rect 32965 15385 32999 15419
rect 5089 15317 5123 15351
rect 5257 15317 5291 15351
rect 6837 15317 6871 15351
rect 23029 15317 23063 15351
rect 33517 15317 33551 15351
rect 5448 15113 5482 15147
rect 16037 15113 16071 15147
rect 22293 15113 22327 15147
rect 23489 15113 23523 15147
rect 33609 15113 33643 15147
rect 5825 15045 5859 15079
rect 9689 15045 9723 15079
rect 17417 15045 17451 15079
rect 23121 15045 23155 15079
rect 23305 15045 23339 15079
rect 29837 15045 29871 15079
rect 4169 14977 4203 15011
rect 9045 14977 9079 15011
rect 9229 14977 9263 15011
rect 10425 14977 10459 15011
rect 10517 14977 10551 15011
rect 10701 14977 10735 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 18245 14977 18279 15011
rect 20637 14977 20671 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 22385 14977 22419 15011
rect 25154 14977 25188 15011
rect 32321 14977 32355 15011
rect 1685 14909 1719 14943
rect 1961 14909 1995 14943
rect 4077 14909 4111 14943
rect 8953 14909 8987 14943
rect 11161 14909 11195 14943
rect 25421 14909 25455 14943
rect 3433 14841 3467 14875
rect 29653 14841 29687 14875
rect 5273 14773 5307 14807
rect 5457 14773 5491 14807
rect 19717 14773 19751 14807
rect 20453 14773 20487 14807
rect 23305 14773 23339 14807
rect 24041 14773 24075 14807
rect 6193 14569 6227 14603
rect 7205 14569 7239 14603
rect 19625 14569 19659 14603
rect 22109 14569 22143 14603
rect 25973 14569 26007 14603
rect 33241 14569 33275 14603
rect 7389 14501 7423 14535
rect 8493 14501 8527 14535
rect 9229 14501 9263 14535
rect 17325 14433 17359 14467
rect 24593 14433 24627 14467
rect 31401 14433 31435 14467
rect 31861 14433 31895 14467
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 6101 14365 6135 14399
rect 6377 14365 6411 14399
rect 7941 14365 7975 14399
rect 12817 14365 12851 14399
rect 12909 14365 12943 14399
rect 15577 14365 15611 14399
rect 17785 14365 17819 14399
rect 18245 14365 18279 14399
rect 18521 14365 18555 14399
rect 20729 14365 20763 14399
rect 20996 14365 21030 14399
rect 24860 14365 24894 14399
rect 26433 14365 26467 14399
rect 28273 14365 28307 14399
rect 28549 14365 28583 14399
rect 31125 14365 31159 14399
rect 32137 14365 32171 14399
rect 2973 14297 3007 14331
rect 7021 14297 7055 14331
rect 8033 14297 8067 14331
rect 8217 14297 8251 14331
rect 9505 14297 9539 14331
rect 9781 14297 9815 14331
rect 13093 14297 13127 14331
rect 19441 14297 19475 14331
rect 26700 14297 26734 14331
rect 28733 14297 28767 14331
rect 29745 14297 29779 14331
rect 6561 14229 6595 14263
rect 7231 14229 7265 14263
rect 9689 14229 9723 14263
rect 19625 14229 19659 14263
rect 19809 14229 19843 14263
rect 27813 14229 27847 14263
rect 28365 14229 28399 14263
rect 2605 14025 2639 14059
rect 5917 14025 5951 14059
rect 22017 14025 22051 14059
rect 29101 14025 29135 14059
rect 30113 14025 30147 14059
rect 31401 14025 31435 14059
rect 4445 13957 4479 13991
rect 6561 13957 6595 13991
rect 6745 13957 6779 13991
rect 12081 13957 12115 13991
rect 17601 13957 17635 13991
rect 19073 13957 19107 13991
rect 19984 13957 20018 13991
rect 22293 13957 22327 13991
rect 24685 13957 24719 13991
rect 27491 13957 27525 13991
rect 27629 13957 27663 13991
rect 28733 13957 28767 13991
rect 28917 13957 28951 13991
rect 29745 13957 29779 13991
rect 2697 13889 2731 13923
rect 7021 13889 7055 13923
rect 9597 13889 9631 13923
rect 9781 13889 9815 13923
rect 14197 13889 14231 13923
rect 14381 13889 14415 13923
rect 15393 13889 15427 13923
rect 16313 13889 16347 13923
rect 16865 13889 16899 13923
rect 17325 13889 17359 13923
rect 18797 13889 18831 13923
rect 19717 13889 19751 13923
rect 22201 13889 22235 13923
rect 22385 13889 22419 13923
rect 22569 13889 22603 13923
rect 24593 13889 24627 13923
rect 24869 13889 24903 13923
rect 27721 13889 27755 13923
rect 27813 13889 27847 13923
rect 29653 13889 29687 13923
rect 29929 13889 29963 13923
rect 31325 13879 31359 13913
rect 31585 13889 31619 13923
rect 31769 13889 31803 13923
rect 32597 13889 32631 13923
rect 4169 13821 4203 13855
rect 9873 13821 9907 13855
rect 11805 13821 11839 13855
rect 13553 13821 13587 13855
rect 14105 13821 14139 13855
rect 27353 13821 27387 13855
rect 27997 13821 28031 13855
rect 32321 13821 32355 13855
rect 33701 13821 33735 13855
rect 16037 13753 16071 13787
rect 21097 13753 21131 13787
rect 25053 13753 25087 13787
rect 6745 13685 6779 13719
rect 28917 13685 28951 13719
rect 3433 13481 3467 13515
rect 5549 13481 5583 13515
rect 15669 13481 15703 13515
rect 27353 13481 27387 13515
rect 31677 13481 31711 13515
rect 2973 13345 3007 13379
rect 9137 13345 9171 13379
rect 12081 13345 12115 13379
rect 13553 13345 13587 13379
rect 18521 13345 18555 13379
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 4629 13277 4663 13311
rect 5365 13277 5399 13311
rect 5641 13277 5675 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 11805 13277 11839 13311
rect 15117 13277 15151 13311
rect 15485 13277 15519 13311
rect 16405 13277 16439 13311
rect 18061 13277 18095 13311
rect 18337 13277 18371 13311
rect 20269 13277 20303 13311
rect 26065 13277 26099 13311
rect 32965 13277 32999 13311
rect 4261 13209 4295 13243
rect 8585 13209 8619 13243
rect 9413 13209 9447 13243
rect 16221 13209 16255 13243
rect 16773 13209 16807 13243
rect 2421 13141 2455 13175
rect 10885 13141 10919 13175
rect 21557 13141 21591 13175
rect 3893 12937 3927 12971
rect 4353 12937 4387 12971
rect 22937 12937 22971 12971
rect 27905 12937 27939 12971
rect 28733 12937 28767 12971
rect 32321 12937 32355 12971
rect 32689 12937 32723 12971
rect 2421 12869 2455 12903
rect 9413 12869 9447 12903
rect 13001 12869 13035 12903
rect 14749 12869 14783 12903
rect 19165 12869 19199 12903
rect 22661 12869 22695 12903
rect 27537 12869 27571 12903
rect 27629 12869 27663 12903
rect 2145 12801 2179 12835
rect 4353 12801 4387 12835
rect 4537 12801 4571 12835
rect 9689 12801 9723 12835
rect 15393 12801 15427 12835
rect 16037 12801 16071 12835
rect 17601 12801 17635 12835
rect 18061 12801 18095 12835
rect 18797 12801 18831 12835
rect 18981 12801 19015 12835
rect 19973 12801 20007 12835
rect 22293 12801 22327 12835
rect 22386 12801 22420 12835
rect 22569 12801 22603 12835
rect 22799 12801 22833 12835
rect 27261 12801 27295 12835
rect 27409 12801 27443 12835
rect 27767 12801 27801 12835
rect 28549 12801 28583 12835
rect 28825 12801 28859 12835
rect 29745 12801 29779 12835
rect 32505 12801 32539 12835
rect 32781 12801 32815 12835
rect 16129 12733 16163 12767
rect 18337 12733 18371 12767
rect 19717 12733 19751 12767
rect 29561 12733 29595 12767
rect 7941 12597 7975 12631
rect 21097 12597 21131 12631
rect 28365 12597 28399 12631
rect 3065 12393 3099 12427
rect 19901 12393 19935 12427
rect 22109 12393 22143 12427
rect 23029 12393 23063 12427
rect 16681 12257 16715 12291
rect 3065 12189 3099 12223
rect 3157 12189 3191 12223
rect 14565 12189 14599 12223
rect 15209 12189 15243 12223
rect 15945 12189 15979 12223
rect 16589 12189 16623 12223
rect 17509 12189 17543 12223
rect 17969 12189 18003 12223
rect 18245 12189 18279 12223
rect 19441 12189 19475 12223
rect 19533 12189 19567 12223
rect 19717 12189 19751 12223
rect 23213 12189 23247 12223
rect 23305 12189 23339 12223
rect 23489 12189 23523 12223
rect 23581 12189 23615 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 28135 12189 28169 12223
rect 28548 12189 28582 12223
rect 28641 12189 28675 12223
rect 15025 12121 15059 12155
rect 20821 12121 20855 12155
rect 28273 12121 28307 12155
rect 28365 12121 28399 12155
rect 24593 12053 24627 12087
rect 24961 12053 24995 12087
rect 27997 12053 28031 12087
rect 17141 11849 17175 11883
rect 22385 11849 22419 11883
rect 25237 11849 25271 11883
rect 31217 11849 31251 11883
rect 32689 11849 32723 11883
rect 15761 11781 15795 11815
rect 16313 11781 16347 11815
rect 22753 11781 22787 11815
rect 24124 11781 24158 11815
rect 25697 11781 25731 11815
rect 25881 11781 25915 11815
rect 27712 11781 27746 11815
rect 14197 11713 14231 11747
rect 14749 11713 14783 11747
rect 15945 11713 15979 11747
rect 16865 11713 16899 11747
rect 17049 11713 17083 11747
rect 17693 11713 17727 11747
rect 18153 11713 18187 11747
rect 20352 11713 20386 11747
rect 22569 11713 22603 11747
rect 22661 11713 22695 11747
rect 22937 11713 22971 11747
rect 31125 11713 31159 11747
rect 31401 11713 31435 11747
rect 32505 11713 32539 11747
rect 32781 11713 32815 11747
rect 18429 11645 18463 11679
rect 20085 11645 20119 11679
rect 23857 11645 23891 11679
rect 27445 11645 27479 11679
rect 14289 11577 14323 11611
rect 21465 11577 21499 11611
rect 28825 11577 28859 11611
rect 25881 11509 25915 11543
rect 26065 11509 26099 11543
rect 31585 11509 31619 11543
rect 32321 11509 32355 11543
rect 4169 11305 4203 11339
rect 20545 11305 20579 11339
rect 21005 11305 21039 11339
rect 31493 11305 31527 11339
rect 13645 11237 13679 11271
rect 18245 11169 18279 11203
rect 5549 11101 5583 11135
rect 10333 11101 10367 11135
rect 10600 11101 10634 11135
rect 12725 11101 12759 11135
rect 13093 11101 13127 11135
rect 16773 11101 16807 11135
rect 16957 11101 16991 11135
rect 17509 11101 17543 11135
rect 17969 11101 18003 11135
rect 19901 11101 19935 11135
rect 20049 11101 20083 11135
rect 20177 11101 20211 11135
rect 20366 11101 20400 11135
rect 21189 11101 21223 11135
rect 21373 11101 21407 11135
rect 21465 11101 21499 11135
rect 23765 11101 23799 11135
rect 23949 11101 23983 11135
rect 24041 11101 24075 11135
rect 26065 11101 26099 11135
rect 29929 11101 29963 11135
rect 30205 11101 30239 11135
rect 32873 11101 32907 11135
rect 3985 11033 4019 11067
rect 5816 11033 5850 11067
rect 12633 11033 12667 11067
rect 13461 11033 13495 11067
rect 16681 11033 16715 11067
rect 20269 11033 20303 11067
rect 23581 11033 23615 11067
rect 30113 11033 30147 11067
rect 32606 11033 32640 11067
rect 4185 10965 4219 10999
rect 4353 10965 4387 10999
rect 6929 10965 6963 10999
rect 11713 10965 11747 10999
rect 12357 10965 12391 10999
rect 27353 10965 27387 10999
rect 29745 10965 29779 10999
rect 7941 10761 7975 10795
rect 9965 10761 9999 10795
rect 13645 10761 13679 10795
rect 25605 10761 25639 10795
rect 28181 10761 28215 10795
rect 29929 10761 29963 10795
rect 33701 10761 33735 10795
rect 6837 10693 6871 10727
rect 7113 10693 7147 10727
rect 7205 10693 7239 10727
rect 7573 10693 7607 10727
rect 8861 10693 8895 10727
rect 9096 10693 9130 10727
rect 9229 10693 9263 10727
rect 9597 10693 9631 10727
rect 12541 10693 12575 10727
rect 12909 10693 12943 10727
rect 13277 10693 13311 10727
rect 18245 10693 18279 10727
rect 19993 10693 20027 10727
rect 25145 10693 25179 10727
rect 28641 10693 28675 10727
rect 30849 10693 30883 10727
rect 31033 10693 31067 10727
rect 32566 10693 32600 10727
rect 3249 10625 3283 10659
rect 3433 10625 3467 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 12817 10625 12851 10659
rect 25743 10625 25777 10659
rect 25881 10625 25915 10659
rect 25973 10625 26007 10659
rect 26156 10625 26190 10659
rect 26249 10625 26283 10659
rect 27537 10625 27571 10659
rect 27685 10625 27719 10659
rect 27813 10625 27847 10659
rect 27905 10625 27939 10659
rect 28043 10625 28077 10659
rect 3157 10557 3191 10591
rect 3341 10557 3375 10591
rect 32321 10557 32355 10591
rect 4077 10489 4111 10523
rect 2973 10421 3007 10455
rect 8125 10421 8159 10455
rect 10149 10421 10183 10455
rect 13829 10421 13863 10455
rect 23857 10421 23891 10455
rect 31033 10421 31067 10455
rect 31217 10421 31251 10455
rect 4169 10217 4203 10251
rect 6745 10217 6779 10251
rect 8585 10217 8619 10251
rect 12633 10217 12667 10251
rect 21281 10217 21315 10251
rect 25973 10217 26007 10251
rect 29745 10217 29779 10251
rect 31677 10217 31711 10251
rect 4353 10149 4387 10183
rect 27353 10149 27387 10183
rect 3249 10081 3283 10115
rect 5365 10081 5399 10115
rect 7205 10081 7239 10115
rect 11253 10081 11287 10115
rect 24593 10081 24627 10115
rect 28733 10081 28767 10115
rect 2237 10013 2271 10047
rect 2697 10013 2731 10047
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 3341 10013 3375 10047
rect 7472 10013 7506 10047
rect 17049 10013 17083 10047
rect 17325 10013 17359 10047
rect 20637 10013 20671 10047
rect 20730 10013 20764 10047
rect 20913 10013 20947 10047
rect 21102 10013 21136 10047
rect 24860 10013 24894 10047
rect 28477 10013 28511 10047
rect 29929 10013 29963 10047
rect 30113 10013 30147 10047
rect 30297 10013 30331 10047
rect 33425 10013 33459 10047
rect 33701 10013 33735 10047
rect 3985 9945 4019 9979
rect 4201 9945 4235 9979
rect 5632 9945 5666 9979
rect 11520 9945 11554 9979
rect 17233 9945 17267 9979
rect 21005 9945 21039 9979
rect 30021 9945 30055 9979
rect 32965 9945 32999 9979
rect 2145 9877 2179 9911
rect 3065 9877 3099 9911
rect 16865 9877 16899 9911
rect 33517 9877 33551 9911
rect 33885 9877 33919 9911
rect 4261 9673 4295 9707
rect 8585 9673 8619 9707
rect 27721 9673 27755 9707
rect 2329 9605 2363 9639
rect 3341 9605 3375 9639
rect 4077 9605 4111 9639
rect 7472 9605 7506 9639
rect 27353 9605 27387 9639
rect 27445 9605 27479 9639
rect 31401 9605 31435 9639
rect 32321 9605 32355 9639
rect 2145 9537 2179 9571
rect 2421 9537 2455 9571
rect 3249 9537 3283 9571
rect 4537 9537 4571 9571
rect 4997 9537 5031 9571
rect 7205 9537 7239 9571
rect 11969 9537 12003 9571
rect 17601 9537 17635 9571
rect 17785 9537 17819 9571
rect 17877 9537 17911 9571
rect 18337 9537 18371 9571
rect 18521 9537 18555 9571
rect 18613 9537 18647 9571
rect 18705 9537 18739 9571
rect 19441 9537 19475 9571
rect 19625 9537 19659 9571
rect 19717 9537 19751 9571
rect 19809 9537 19843 9571
rect 20637 9537 20671 9571
rect 20821 9537 20855 9571
rect 20913 9537 20947 9571
rect 27169 9537 27203 9571
rect 27537 9537 27571 9571
rect 31309 9537 31343 9571
rect 31585 9537 31619 9571
rect 3525 9469 3559 9503
rect 11713 9469 11747 9503
rect 5089 9401 5123 9435
rect 13093 9401 13127 9435
rect 18889 9401 18923 9435
rect 19993 9401 20027 9435
rect 1961 9333 1995 9367
rect 2881 9333 2915 9367
rect 4261 9333 4295 9367
rect 17417 9333 17451 9367
rect 20453 9333 20487 9367
rect 31769 9333 31803 9367
rect 33609 9333 33643 9367
rect 2973 9129 3007 9163
rect 12173 9129 12207 9163
rect 16405 9129 16439 9163
rect 21281 9129 21315 9163
rect 32321 9129 32355 9163
rect 2789 9061 2823 9095
rect 3985 8993 4019 9027
rect 10793 8993 10827 9027
rect 3341 8925 3375 8959
rect 4169 8925 4203 8959
rect 11060 8925 11094 8959
rect 15025 8925 15059 8959
rect 16865 8925 16899 8959
rect 19901 8925 19935 8959
rect 20168 8925 20202 8959
rect 22661 8925 22695 8959
rect 22845 8925 22879 8959
rect 22937 8925 22971 8959
rect 24593 8925 24627 8959
rect 24869 8925 24903 8959
rect 28733 8925 28767 8959
rect 28825 8925 28859 8959
rect 29009 8925 29043 8959
rect 29929 8925 29963 8959
rect 30205 8925 30239 8959
rect 33701 8925 33735 8959
rect 2927 8857 2961 8891
rect 15292 8857 15326 8891
rect 17132 8857 17166 8891
rect 24685 8857 24719 8891
rect 30113 8857 30147 8891
rect 33456 8857 33490 8891
rect 4353 8789 4387 8823
rect 18245 8789 18279 8823
rect 22477 8789 22511 8823
rect 25053 8789 25087 8823
rect 29193 8789 29227 8823
rect 29745 8789 29779 8823
rect 2697 8585 2731 8619
rect 3065 8585 3099 8619
rect 3617 8585 3651 8619
rect 14933 8585 14967 8619
rect 23673 8585 23707 8619
rect 25881 8585 25915 8619
rect 30021 8585 30055 8619
rect 33701 8585 33735 8619
rect 9597 8517 9631 8551
rect 16068 8517 16102 8551
rect 20637 8517 20671 8551
rect 20729 8517 20763 8551
rect 22753 8517 22787 8551
rect 22937 8517 22971 8551
rect 24808 8517 24842 8551
rect 30481 8517 30515 8551
rect 32566 8517 32600 8551
rect 2605 8449 2639 8483
rect 2881 8449 2915 8483
rect 3709 8449 3743 8483
rect 16313 8449 16347 8483
rect 17509 8449 17543 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 18245 8449 18279 8483
rect 20453 8449 20487 8483
rect 20821 8449 20855 8483
rect 25513 8449 25547 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 28641 8449 28675 8483
rect 28908 8449 28942 8483
rect 30665 8449 30699 8483
rect 30849 8449 30883 8483
rect 30941 8449 30975 8483
rect 32321 8449 32355 8483
rect 19993 8381 20027 8415
rect 25053 8381 25087 8415
rect 17325 8313 17359 8347
rect 21005 8313 21039 8347
rect 23121 8313 23155 8347
rect 8125 8245 8159 8279
rect 22937 8245 22971 8279
rect 22937 8041 22971 8075
rect 28273 8041 28307 8075
rect 32413 8041 32447 8075
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 9781 7837 9815 7871
rect 9965 7837 9999 7871
rect 19441 7837 19475 7871
rect 24593 7837 24627 7871
rect 28549 7837 28583 7871
rect 29745 7837 29779 7871
rect 33701 7837 33735 7871
rect 7389 7769 7423 7803
rect 10149 7769 10183 7803
rect 16313 7769 16347 7803
rect 21649 7769 21683 7803
rect 28089 7769 28123 7803
rect 28273 7769 28307 7803
rect 17601 7701 17635 7735
rect 20729 7701 20763 7735
rect 25881 7701 25915 7735
rect 31033 7701 31067 7735
rect 10701 7497 10735 7531
rect 12173 7497 12207 7531
rect 15945 7497 15979 7531
rect 17325 7497 17359 7531
rect 19533 7497 19567 7531
rect 20637 7497 20671 7531
rect 20821 7497 20855 7531
rect 22385 7497 22419 7531
rect 25973 7497 26007 7531
rect 29101 7497 29135 7531
rect 6837 7429 6871 7463
rect 15577 7429 15611 7463
rect 15761 7429 15795 7463
rect 18245 7429 18279 7463
rect 20453 7429 20487 7463
rect 23397 7429 23431 7463
rect 25053 7429 25087 7463
rect 2697 7361 2731 7395
rect 8953 7361 8987 7395
rect 14749 7361 14783 7395
rect 17509 7361 17543 7395
rect 17693 7361 17727 7395
rect 17785 7361 17819 7395
rect 22201 7361 22235 7395
rect 22477 7361 22511 7395
rect 25789 7361 25823 7395
rect 26065 7361 26099 7395
rect 30389 7361 30423 7395
rect 6561 7293 6595 7327
rect 9229 7293 9263 7327
rect 11897 7293 11931 7327
rect 12081 7293 12115 7327
rect 2605 7157 2639 7191
rect 8309 7157 8343 7191
rect 12541 7157 12575 7191
rect 13461 7157 13495 7191
rect 15761 7157 15795 7191
rect 20637 7157 20671 7191
rect 22017 7157 22051 7191
rect 25605 7157 25639 7191
rect 1856 6953 1890 6987
rect 13093 6953 13127 6987
rect 1593 6817 1627 6851
rect 3341 6817 3375 6851
rect 5457 6817 5491 6851
rect 7941 6817 7975 6851
rect 10149 6817 10183 6851
rect 10701 6817 10735 6851
rect 15577 6817 15611 6851
rect 21281 6817 21315 6851
rect 5724 6749 5758 6783
rect 10241 6749 10275 6783
rect 10563 6749 10597 6783
rect 11713 6749 11747 6783
rect 13553 6749 13587 6783
rect 13737 6749 13771 6783
rect 17601 6749 17635 6783
rect 17877 6749 17911 6783
rect 19441 6749 19475 6783
rect 19708 6749 19742 6783
rect 21548 6749 21582 6783
rect 23765 6749 23799 6783
rect 23949 6749 23983 6783
rect 24041 6749 24075 6783
rect 24593 6749 24627 6783
rect 28926 6749 28960 6783
rect 29193 6749 29227 6783
rect 30113 6749 30147 6783
rect 7757 6681 7791 6715
rect 11958 6681 11992 6715
rect 15844 6681 15878 6715
rect 17417 6681 17451 6715
rect 17785 6681 17819 6715
rect 24860 6681 24894 6715
rect 30358 6681 30392 6715
rect 6837 6613 6871 6647
rect 7297 6613 7331 6647
rect 7665 6613 7699 6647
rect 10977 6613 11011 6647
rect 13645 6613 13679 6647
rect 16957 6613 16991 6647
rect 20821 6613 20855 6647
rect 22661 6613 22695 6647
rect 23581 6613 23615 6647
rect 25973 6613 26007 6647
rect 27813 6613 27847 6647
rect 31493 6613 31527 6647
rect 6929 6409 6963 6443
rect 13001 6409 13035 6443
rect 21005 6409 21039 6443
rect 2789 6341 2823 6375
rect 3709 6341 3743 6375
rect 6837 6341 6871 6375
rect 12909 6341 12943 6375
rect 19892 6341 19926 6375
rect 24694 6341 24728 6375
rect 29570 6341 29604 6375
rect 2973 6273 3007 6307
rect 3157 6273 3191 6307
rect 6653 6205 6687 6239
rect 12725 6205 12759 6239
rect 19625 6205 19659 6239
rect 24961 6205 24995 6239
rect 29837 6205 29871 6239
rect 7297 6137 7331 6171
rect 23581 6137 23615 6171
rect 28457 6137 28491 6171
rect 3801 6069 3835 6103
rect 13369 6069 13403 6103
rect 25973 5865 26007 5899
rect 29193 5865 29227 5899
rect 3985 5729 4019 5763
rect 4353 5729 4387 5763
rect 24593 5661 24627 5695
rect 24860 5661 24894 5695
rect 28733 5661 28767 5695
rect 29009 5661 29043 5695
rect 28825 5593 28859 5627
rect 6101 5525 6135 5559
rect 5641 5321 5675 5355
rect 10517 5321 10551 5355
rect 19533 5321 19567 5355
rect 24685 5321 24719 5355
rect 4353 5253 4387 5287
rect 9505 5253 9539 5287
rect 18245 5253 18279 5287
rect 23397 5253 23431 5287
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 5733 5185 5767 5219
rect 9597 5185 9631 5219
rect 10425 5185 10459 5219
rect 10609 5185 10643 5219
rect 11969 5185 12003 5219
rect 13553 5185 13587 5219
rect 15209 5185 15243 5219
rect 25789 5185 25823 5219
rect 25973 5185 26007 5219
rect 9321 5117 9355 5151
rect 11713 5117 11747 5151
rect 13829 5117 13863 5151
rect 9965 4981 9999 5015
rect 13093 4981 13127 5015
rect 13645 4981 13679 5015
rect 13737 4981 13771 5015
rect 15117 4981 15151 5015
rect 25605 4981 25639 5015
rect 10885 4777 10919 4811
rect 11989 4777 12023 4811
rect 14565 4709 14599 4743
rect 24685 4709 24719 4743
rect 7205 4641 7239 4675
rect 9137 4641 9171 4675
rect 9413 4641 9447 4675
rect 16221 4641 16255 4675
rect 18705 4641 18739 4675
rect 20453 4641 20487 4675
rect 25053 4641 25087 4675
rect 7472 4573 7506 4607
rect 11897 4573 11931 4607
rect 12265 4573 12299 4607
rect 14289 4573 14323 4607
rect 14565 4573 14599 4607
rect 15945 4573 15979 4607
rect 17417 4573 17451 4607
rect 18429 4573 18463 4607
rect 20177 4573 20211 4607
rect 21649 4573 21683 4607
rect 22293 4573 22327 4607
rect 25881 4573 25915 4607
rect 26148 4505 26182 4539
rect 8585 4437 8619 4471
rect 12449 4437 12483 4471
rect 14381 4437 14415 4471
rect 15577 4437 15611 4471
rect 16037 4437 16071 4471
rect 17509 4437 17543 4471
rect 18061 4437 18095 4471
rect 18521 4437 18555 4471
rect 19809 4437 19843 4471
rect 20269 4437 20303 4471
rect 21557 4437 21591 4471
rect 22201 4437 22235 4471
rect 24593 4437 24627 4471
rect 27261 4437 27295 4471
rect 9321 4233 9355 4267
rect 9689 4233 9723 4267
rect 26157 4233 26191 4267
rect 7389 4165 7423 4199
rect 13369 4165 13403 4199
rect 15200 4165 15234 4199
rect 9781 4097 9815 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 10885 4097 10919 4131
rect 13461 4097 13495 4131
rect 14933 4097 14967 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 17960 4097 17994 4131
rect 21198 4097 21232 4131
rect 21465 4097 21499 4131
rect 22017 4097 22051 4131
rect 22284 4097 22318 4131
rect 24317 4097 24351 4131
rect 24584 4097 24618 4131
rect 26617 4097 26651 4131
rect 27169 4097 27203 4131
rect 27436 4097 27470 4131
rect 7113 4029 7147 4063
rect 8861 4029 8895 4063
rect 9965 4029 9999 4063
rect 13645 4029 13679 4063
rect 26249 3961 26283 3995
rect 13001 3893 13035 3927
rect 16313 3893 16347 3927
rect 16957 3893 16991 3927
rect 19073 3893 19107 3927
rect 20085 3893 20119 3927
rect 23397 3893 23431 3927
rect 25697 3893 25731 3927
rect 28549 3893 28583 3927
rect 7941 3689 7975 3723
rect 13737 3689 13771 3723
rect 20821 3689 20855 3723
rect 22109 3689 22143 3723
rect 24593 3689 24627 3723
rect 27077 3689 27111 3723
rect 27813 3689 27847 3723
rect 26801 3621 26835 3655
rect 26893 3621 26927 3655
rect 27905 3621 27939 3655
rect 16681 3553 16715 3587
rect 22753 3553 22787 3587
rect 26985 3553 27019 3587
rect 28273 3553 28307 3587
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 12357 3485 12391 3519
rect 12624 3485 12658 3519
rect 15669 3485 15703 3519
rect 19441 3485 19475 3519
rect 22477 3485 22511 3519
rect 22569 3485 22603 3519
rect 25706 3485 25740 3519
rect 25973 3485 26007 3519
rect 26433 3485 26467 3519
rect 15402 3417 15436 3451
rect 16948 3417 16982 3451
rect 19708 3417 19742 3451
rect 14289 3349 14323 3383
rect 18061 3349 18095 3383
rect 12541 3145 12575 3179
rect 14381 3145 14415 3179
rect 14749 3145 14783 3179
rect 15301 3145 15335 3179
rect 16957 3145 16991 3179
rect 17325 3145 17359 3179
rect 17417 3145 17451 3179
rect 19625 3145 19659 3179
rect 20729 3145 20763 3179
rect 29101 3145 29135 3179
rect 21097 3077 21131 3111
rect 30389 3077 30423 3111
rect 12633 3009 12667 3043
rect 15209 3009 15243 3043
rect 19717 3009 19751 3043
rect 20913 3009 20947 3043
rect 21189 3009 21223 3043
rect 25145 3009 25179 3043
rect 26065 3009 26099 3043
rect 14197 2941 14231 2975
rect 14289 2941 14323 2975
rect 17601 2941 17635 2975
rect 25513 2941 25547 2975
rect 25605 2873 25639 2907
rect 25697 2805 25731 2839
rect 2053 2397 2087 2431
rect 3065 2397 3099 2431
rect 4445 2397 4479 2431
rect 5641 2397 5675 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 11713 2397 11747 2431
rect 12909 2397 12943 2431
rect 14289 2397 14323 2431
rect 15485 2397 15519 2431
rect 16865 2397 16899 2431
rect 18061 2397 18095 2431
rect 19441 2397 19475 2431
rect 20637 2397 20671 2431
rect 22017 2397 22051 2431
rect 23213 2397 23247 2431
rect 25053 2397 25087 2431
rect 26249 2397 26283 2431
rect 27629 2397 27663 2431
rect 28365 2397 28399 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 32321 2397 32355 2431
rect 33517 2397 33551 2431
rect 1777 2329 1811 2363
rect 2789 2329 2823 2363
rect 4169 2329 4203 2363
rect 5365 2329 5399 2363
rect 14565 2329 14599 2363
rect 15761 2329 15795 2363
rect 17141 2329 17175 2363
rect 18337 2329 18371 2363
rect 19717 2329 19751 2363
rect 20913 2329 20947 2363
rect 22293 2329 22327 2363
rect 23489 2329 23523 2363
rect 24777 2329 24811 2363
rect 25973 2329 26007 2363
rect 27353 2329 27387 2363
rect 28641 2329 28675 2363
rect 34345 2261 34379 2295
<< metal1 >>
rect 1104 33754 35027 33776
rect 1104 33702 9390 33754
rect 9442 33702 9454 33754
rect 9506 33702 9518 33754
rect 9570 33702 9582 33754
rect 9634 33702 9646 33754
rect 9698 33702 17831 33754
rect 17883 33702 17895 33754
rect 17947 33702 17959 33754
rect 18011 33702 18023 33754
rect 18075 33702 18087 33754
rect 18139 33702 26272 33754
rect 26324 33702 26336 33754
rect 26388 33702 26400 33754
rect 26452 33702 26464 33754
rect 26516 33702 26528 33754
rect 26580 33702 34713 33754
rect 34765 33702 34777 33754
rect 34829 33702 34841 33754
rect 34893 33702 34905 33754
rect 34957 33702 34969 33754
rect 35021 33702 35027 33754
rect 1104 33680 35027 33702
rect 4890 33572 4896 33584
rect 4851 33544 4896 33572
rect 4890 33532 4896 33544
rect 4948 33532 4954 33584
rect 7834 33572 7840 33584
rect 7795 33544 7840 33572
rect 7834 33532 7840 33544
rect 7892 33532 7898 33584
rect 10594 33532 10600 33584
rect 10652 33572 10658 33584
rect 10781 33575 10839 33581
rect 10781 33572 10793 33575
rect 10652 33544 10793 33572
rect 10652 33532 10658 33544
rect 10781 33541 10793 33544
rect 10827 33541 10839 33575
rect 10781 33535 10839 33541
rect 13814 33532 13820 33584
rect 13872 33572 13878 33584
rect 14461 33575 14519 33581
rect 14461 33572 14473 33575
rect 13872 33544 14473 33572
rect 13872 33532 13878 33544
rect 14461 33541 14473 33544
rect 14507 33541 14519 33575
rect 14461 33535 14519 33541
rect 16574 33532 16580 33584
rect 16632 33572 16638 33584
rect 17037 33575 17095 33581
rect 17037 33572 17049 33575
rect 16632 33544 17049 33572
rect 16632 33532 16638 33544
rect 17037 33541 17049 33544
rect 17083 33541 17095 33575
rect 17037 33535 17095 33541
rect 19426 33532 19432 33584
rect 19484 33572 19490 33584
rect 19705 33575 19763 33581
rect 19705 33572 19717 33575
rect 19484 33544 19717 33572
rect 19484 33532 19490 33544
rect 19705 33541 19717 33544
rect 19751 33541 19763 33575
rect 22646 33572 22652 33584
rect 22607 33544 22652 33572
rect 19705 33535 19763 33541
rect 22646 33532 22652 33544
rect 22704 33532 22710 33584
rect 25590 33572 25596 33584
rect 25551 33544 25596 33572
rect 25590 33532 25596 33544
rect 25648 33532 25654 33584
rect 28534 33572 28540 33584
rect 28495 33544 28540 33572
rect 28534 33532 28540 33544
rect 28592 33532 28598 33584
rect 31478 33572 31484 33584
rect 31439 33544 31484 33572
rect 31478 33532 31484 33544
rect 31536 33532 31542 33584
rect 34238 33572 34244 33584
rect 34199 33544 34244 33572
rect 34238 33532 34244 33544
rect 34296 33532 34302 33584
rect 8018 33368 8024 33380
rect 7979 33340 8024 33368
rect 8018 33328 8024 33340
rect 8076 33328 8082 33380
rect 10965 33371 11023 33377
rect 10965 33337 10977 33371
rect 11011 33368 11023 33371
rect 12250 33368 12256 33380
rect 11011 33340 12256 33368
rect 11011 33337 11023 33340
rect 10965 33331 11023 33337
rect 12250 33328 12256 33340
rect 12308 33328 12314 33380
rect 14274 33368 14280 33380
rect 14235 33340 14280 33368
rect 14274 33328 14280 33340
rect 14332 33328 14338 33380
rect 16850 33368 16856 33380
rect 16811 33340 16856 33368
rect 16850 33328 16856 33340
rect 16908 33328 16914 33380
rect 19518 33368 19524 33380
rect 19479 33340 19524 33368
rect 19518 33328 19524 33340
rect 19576 33328 19582 33380
rect 20254 33328 20260 33380
rect 20312 33368 20318 33380
rect 22465 33371 22523 33377
rect 22465 33368 22477 33371
rect 20312 33340 22477 33368
rect 20312 33328 20318 33340
rect 22465 33337 22477 33340
rect 22511 33337 22523 33371
rect 25406 33368 25412 33380
rect 25367 33340 25412 33368
rect 22465 33331 22523 33337
rect 25406 33328 25412 33340
rect 25464 33328 25470 33380
rect 31294 33368 31300 33380
rect 31255 33340 31300 33368
rect 31294 33328 31300 33340
rect 31352 33328 31358 33380
rect 33318 33328 33324 33380
rect 33376 33368 33382 33380
rect 34057 33371 34115 33377
rect 34057 33368 34069 33371
rect 33376 33340 34069 33368
rect 33376 33328 33382 33340
rect 34057 33337 34069 33340
rect 34103 33337 34115 33371
rect 34057 33331 34115 33337
rect 4982 33300 4988 33312
rect 4943 33272 4988 33300
rect 4982 33260 4988 33272
rect 5040 33260 5046 33312
rect 20438 33260 20444 33312
rect 20496 33300 20502 33312
rect 28445 33303 28503 33309
rect 28445 33300 28457 33303
rect 20496 33272 28457 33300
rect 20496 33260 20502 33272
rect 28445 33269 28457 33272
rect 28491 33269 28503 33303
rect 28445 33263 28503 33269
rect 1104 33210 34868 33232
rect 1104 33158 5170 33210
rect 5222 33158 5234 33210
rect 5286 33158 5298 33210
rect 5350 33158 5362 33210
rect 5414 33158 5426 33210
rect 5478 33158 13611 33210
rect 13663 33158 13675 33210
rect 13727 33158 13739 33210
rect 13791 33158 13803 33210
rect 13855 33158 13867 33210
rect 13919 33158 22052 33210
rect 22104 33158 22116 33210
rect 22168 33158 22180 33210
rect 22232 33158 22244 33210
rect 22296 33158 22308 33210
rect 22360 33158 30493 33210
rect 30545 33158 30557 33210
rect 30609 33158 30621 33210
rect 30673 33158 30685 33210
rect 30737 33158 30749 33210
rect 30801 33158 34868 33210
rect 1104 33136 34868 33158
rect 12066 33056 12072 33108
rect 12124 33096 12130 33108
rect 12124 33068 16712 33096
rect 12124 33056 12130 33068
rect 16684 33028 16712 33068
rect 20254 33028 20260 33040
rect 16684 33000 20260 33028
rect 20254 32988 20260 33000
rect 20312 32988 20318 33040
rect 16577 32963 16635 32969
rect 16577 32929 16589 32963
rect 16623 32960 16635 32963
rect 20438 32960 20444 32972
rect 16623 32932 20444 32960
rect 16623 32929 16635 32932
rect 16577 32923 16635 32929
rect 20438 32920 20444 32932
rect 20496 32920 20502 32972
rect 20622 32960 20628 32972
rect 20583 32932 20628 32960
rect 20622 32920 20628 32932
rect 20680 32920 20686 32972
rect 24578 32960 24584 32972
rect 21928 32932 24584 32960
rect 10229 32895 10287 32901
rect 10229 32861 10241 32895
rect 10275 32892 10287 32895
rect 10502 32892 10508 32904
rect 10275 32864 10508 32892
rect 10275 32861 10287 32864
rect 10229 32855 10287 32861
rect 10502 32852 10508 32864
rect 10560 32852 10566 32904
rect 16301 32895 16359 32901
rect 16301 32861 16313 32895
rect 16347 32861 16359 32895
rect 16301 32855 16359 32861
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32892 16543 32895
rect 16850 32892 16856 32904
rect 16531 32864 16856 32892
rect 16531 32861 16543 32864
rect 16485 32855 16543 32861
rect 15841 32827 15899 32833
rect 15841 32793 15853 32827
rect 15887 32824 15899 32827
rect 16206 32824 16212 32836
rect 15887 32796 16212 32824
rect 15887 32793 15899 32796
rect 15841 32787 15899 32793
rect 16206 32784 16212 32796
rect 16264 32784 16270 32836
rect 16316 32824 16344 32855
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 19334 32852 19340 32904
rect 19392 32892 19398 32904
rect 20533 32895 20591 32901
rect 20533 32892 20545 32895
rect 19392 32864 20545 32892
rect 19392 32852 19398 32864
rect 20533 32861 20545 32864
rect 20579 32892 20591 32895
rect 21928 32892 21956 32932
rect 24578 32920 24584 32932
rect 24636 32920 24642 32972
rect 20579 32864 21956 32892
rect 22465 32895 22523 32901
rect 20579 32861 20591 32864
rect 20533 32855 20591 32861
rect 22465 32861 22477 32895
rect 22511 32892 22523 32895
rect 22830 32892 22836 32904
rect 22511 32864 22836 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 22830 32852 22836 32864
rect 22888 32852 22894 32904
rect 16758 32824 16764 32836
rect 16316 32796 16764 32824
rect 16758 32784 16764 32796
rect 16816 32784 16822 32836
rect 25406 32824 25412 32836
rect 20180 32796 25412 32824
rect 10134 32756 10140 32768
rect 10095 32728 10140 32756
rect 10134 32716 10140 32728
rect 10192 32716 10198 32768
rect 13262 32716 13268 32768
rect 13320 32756 13326 32768
rect 20180 32756 20208 32796
rect 25406 32784 25412 32796
rect 25464 32784 25470 32836
rect 13320 32728 20208 32756
rect 20901 32759 20959 32765
rect 13320 32716 13326 32728
rect 20901 32725 20913 32759
rect 20947 32756 20959 32759
rect 21266 32756 21272 32768
rect 20947 32728 21272 32756
rect 20947 32725 20959 32728
rect 20901 32719 20959 32725
rect 21266 32716 21272 32728
rect 21324 32716 21330 32768
rect 22002 32716 22008 32768
rect 22060 32756 22066 32768
rect 22373 32759 22431 32765
rect 22373 32756 22385 32759
rect 22060 32728 22385 32756
rect 22060 32716 22066 32728
rect 22373 32725 22385 32728
rect 22419 32725 22431 32759
rect 22373 32719 22431 32725
rect 1104 32666 35027 32688
rect 1104 32614 9390 32666
rect 9442 32614 9454 32666
rect 9506 32614 9518 32666
rect 9570 32614 9582 32666
rect 9634 32614 9646 32666
rect 9698 32614 17831 32666
rect 17883 32614 17895 32666
rect 17947 32614 17959 32666
rect 18011 32614 18023 32666
rect 18075 32614 18087 32666
rect 18139 32614 26272 32666
rect 26324 32614 26336 32666
rect 26388 32614 26400 32666
rect 26452 32614 26464 32666
rect 26516 32614 26528 32666
rect 26580 32614 34713 32666
rect 34765 32614 34777 32666
rect 34829 32614 34841 32666
rect 34893 32614 34905 32666
rect 34957 32614 34969 32666
rect 35021 32614 35027 32666
rect 1104 32592 35027 32614
rect 12250 32552 12256 32564
rect 12211 32524 12256 32552
rect 12250 32512 12256 32524
rect 12308 32512 12314 32564
rect 13449 32555 13507 32561
rect 13449 32521 13461 32555
rect 13495 32552 13507 32555
rect 14274 32552 14280 32564
rect 13495 32524 14280 32552
rect 13495 32521 13507 32524
rect 13449 32515 13507 32521
rect 14274 32512 14280 32524
rect 14332 32512 14338 32564
rect 17313 32555 17371 32561
rect 17313 32521 17325 32555
rect 17359 32552 17371 32555
rect 18049 32555 18107 32561
rect 18049 32552 18061 32555
rect 17359 32524 18061 32552
rect 17359 32521 17371 32524
rect 17313 32515 17371 32521
rect 18049 32521 18061 32524
rect 18095 32521 18107 32555
rect 18049 32515 18107 32521
rect 20717 32555 20775 32561
rect 20717 32521 20729 32555
rect 20763 32521 20775 32555
rect 20717 32515 20775 32521
rect 12066 32484 12072 32496
rect 12027 32456 12072 32484
rect 12066 32444 12072 32456
rect 12124 32444 12130 32496
rect 13262 32484 13268 32496
rect 13223 32456 13268 32484
rect 13262 32444 13268 32456
rect 13320 32444 13326 32496
rect 19518 32484 19524 32496
rect 16546 32456 19524 32484
rect 9861 32419 9919 32425
rect 9861 32385 9873 32419
rect 9907 32416 9919 32419
rect 10318 32416 10324 32428
rect 9907 32388 10324 32416
rect 9907 32385 9919 32388
rect 9861 32379 9919 32385
rect 10318 32376 10324 32388
rect 10376 32416 10382 32428
rect 10413 32419 10471 32425
rect 10413 32416 10425 32419
rect 10376 32388 10425 32416
rect 10376 32376 10382 32388
rect 10413 32385 10425 32388
rect 10459 32385 10471 32419
rect 10413 32379 10471 32385
rect 10502 32376 10508 32428
rect 10560 32416 10566 32428
rect 10560 32388 10605 32416
rect 10560 32376 10566 32388
rect 11422 32376 11428 32428
rect 11480 32416 11486 32428
rect 16546 32416 16574 32456
rect 19518 32444 19524 32456
rect 19576 32444 19582 32496
rect 11480 32388 16574 32416
rect 17221 32419 17279 32425
rect 11480 32376 11486 32388
rect 17221 32385 17233 32419
rect 17267 32416 17279 32419
rect 17862 32416 17868 32428
rect 17267 32388 17868 32416
rect 17267 32385 17279 32388
rect 17221 32379 17279 32385
rect 17862 32376 17868 32388
rect 17920 32416 17926 32428
rect 18049 32419 18107 32425
rect 18049 32416 18061 32419
rect 17920 32388 18061 32416
rect 17920 32376 17926 32388
rect 18049 32385 18061 32388
rect 18095 32385 18107 32419
rect 18049 32379 18107 32385
rect 18230 32376 18236 32428
rect 18288 32416 18294 32428
rect 20732 32416 20760 32515
rect 21177 32487 21235 32493
rect 21177 32453 21189 32487
rect 21223 32484 21235 32487
rect 22097 32487 22155 32493
rect 22097 32484 22109 32487
rect 21223 32456 22109 32484
rect 21223 32453 21235 32456
rect 21177 32447 21235 32453
rect 22097 32453 22109 32456
rect 22143 32453 22155 32487
rect 22097 32447 22155 32453
rect 18288 32388 20760 32416
rect 21085 32419 21143 32425
rect 18288 32376 18294 32388
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 22002 32416 22008 32428
rect 21131 32388 22008 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 22462 32416 22468 32428
rect 22235 32388 22468 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 22462 32376 22468 32388
rect 22520 32376 22526 32428
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32385 23075 32419
rect 23198 32416 23204 32428
rect 23159 32388 23204 32416
rect 23017 32379 23075 32385
rect 10689 32351 10747 32357
rect 10689 32317 10701 32351
rect 10735 32317 10747 32351
rect 12342 32348 12348 32360
rect 12255 32320 12348 32348
rect 10689 32311 10747 32317
rect 8570 32240 8576 32292
rect 8628 32280 8634 32292
rect 10704 32280 10732 32311
rect 12342 32308 12348 32320
rect 12400 32348 12406 32360
rect 13541 32351 13599 32357
rect 13541 32348 13553 32351
rect 12400 32320 13553 32348
rect 12400 32308 12406 32320
rect 13541 32317 13553 32320
rect 13587 32348 13599 32351
rect 16758 32348 16764 32360
rect 13587 32320 16764 32348
rect 13587 32317 13599 32320
rect 13541 32311 13599 32317
rect 16758 32308 16764 32320
rect 16816 32308 16822 32360
rect 17402 32348 17408 32360
rect 17363 32320 17408 32348
rect 17402 32308 17408 32320
rect 17460 32308 17466 32360
rect 21266 32348 21272 32360
rect 21227 32320 21272 32348
rect 21266 32308 21272 32320
rect 21324 32308 21330 32360
rect 23032 32348 23060 32379
rect 23198 32376 23204 32388
rect 23256 32376 23262 32428
rect 24486 32416 24492 32428
rect 24447 32388 24492 32416
rect 24486 32376 24492 32388
rect 24544 32376 24550 32428
rect 24578 32376 24584 32428
rect 24636 32416 24642 32428
rect 24673 32419 24731 32425
rect 24673 32416 24685 32419
rect 24636 32388 24685 32416
rect 24636 32376 24642 32388
rect 24673 32385 24685 32388
rect 24719 32385 24731 32419
rect 27706 32416 27712 32428
rect 27667 32388 27712 32416
rect 24673 32379 24731 32385
rect 27706 32376 27712 32388
rect 27764 32376 27770 32428
rect 28074 32416 28080 32428
rect 28035 32388 28080 32416
rect 28074 32376 28080 32388
rect 28132 32376 28138 32428
rect 30469 32419 30527 32425
rect 30469 32385 30481 32419
rect 30515 32416 30527 32419
rect 31294 32416 31300 32428
rect 30515 32388 31300 32416
rect 30515 32385 30527 32388
rect 30469 32379 30527 32385
rect 31294 32376 31300 32388
rect 31352 32376 31358 32428
rect 33318 32416 33324 32428
rect 33279 32388 33324 32416
rect 33318 32376 33324 32388
rect 33376 32376 33382 32428
rect 23382 32348 23388 32360
rect 23032 32320 23388 32348
rect 23382 32308 23388 32320
rect 23440 32308 23446 32360
rect 16853 32283 16911 32289
rect 16853 32280 16865 32283
rect 8628 32252 16865 32280
rect 8628 32240 8634 32252
rect 16853 32249 16865 32252
rect 16899 32249 16911 32283
rect 16853 32243 16911 32249
rect 21082 32240 21088 32292
rect 21140 32280 21146 32292
rect 22925 32283 22983 32289
rect 22925 32280 22937 32283
rect 21140 32252 22937 32280
rect 21140 32240 21146 32252
rect 22925 32249 22937 32252
rect 22971 32249 22983 32283
rect 27157 32283 27215 32289
rect 27157 32280 27169 32283
rect 22925 32243 22983 32249
rect 23032 32252 27169 32280
rect 9861 32215 9919 32221
rect 9861 32181 9873 32215
rect 9907 32212 9919 32215
rect 10042 32212 10048 32224
rect 9907 32184 10048 32212
rect 9907 32181 9919 32184
rect 9861 32175 9919 32181
rect 10042 32172 10048 32184
rect 10100 32172 10106 32224
rect 10594 32172 10600 32224
rect 10652 32212 10658 32224
rect 11793 32215 11851 32221
rect 10652 32184 10697 32212
rect 10652 32172 10658 32184
rect 11793 32181 11805 32215
rect 11839 32212 11851 32215
rect 11882 32212 11888 32224
rect 11839 32184 11888 32212
rect 11839 32181 11851 32184
rect 11793 32175 11851 32181
rect 11882 32172 11888 32184
rect 11940 32172 11946 32224
rect 12989 32215 13047 32221
rect 12989 32181 13001 32215
rect 13035 32212 13047 32215
rect 13170 32212 13176 32224
rect 13035 32184 13176 32212
rect 13035 32181 13047 32184
rect 12989 32175 13047 32181
rect 13170 32172 13176 32184
rect 13228 32172 13234 32224
rect 22830 32172 22836 32224
rect 22888 32212 22894 32224
rect 23032 32212 23060 32252
rect 27157 32249 27169 32252
rect 27203 32249 27215 32283
rect 27157 32243 27215 32249
rect 22888 32184 23060 32212
rect 24581 32215 24639 32221
rect 22888 32172 22894 32184
rect 24581 32181 24593 32215
rect 24627 32212 24639 32215
rect 25038 32212 25044 32224
rect 24627 32184 25044 32212
rect 24627 32181 24639 32184
rect 24581 32175 24639 32181
rect 25038 32172 25044 32184
rect 25096 32172 25102 32224
rect 30190 32172 30196 32224
rect 30248 32212 30254 32224
rect 30285 32215 30343 32221
rect 30285 32212 30297 32215
rect 30248 32184 30297 32212
rect 30248 32172 30254 32184
rect 30285 32181 30297 32184
rect 30331 32181 30343 32215
rect 33134 32212 33140 32224
rect 33095 32184 33140 32212
rect 30285 32175 30343 32181
rect 33134 32172 33140 32184
rect 33192 32172 33198 32224
rect 1104 32122 34868 32144
rect 1104 32070 5170 32122
rect 5222 32070 5234 32122
rect 5286 32070 5298 32122
rect 5350 32070 5362 32122
rect 5414 32070 5426 32122
rect 5478 32070 13611 32122
rect 13663 32070 13675 32122
rect 13727 32070 13739 32122
rect 13791 32070 13803 32122
rect 13855 32070 13867 32122
rect 13919 32070 22052 32122
rect 22104 32070 22116 32122
rect 22168 32070 22180 32122
rect 22232 32070 22244 32122
rect 22296 32070 22308 32122
rect 22360 32070 30493 32122
rect 30545 32070 30557 32122
rect 30609 32070 30621 32122
rect 30673 32070 30685 32122
rect 30737 32070 30749 32122
rect 30801 32070 34868 32122
rect 1104 32048 34868 32070
rect 15749 32011 15807 32017
rect 15749 31977 15761 32011
rect 15795 32008 15807 32011
rect 16114 32008 16120 32020
rect 15795 31980 16120 32008
rect 15795 31977 15807 31980
rect 15749 31971 15807 31977
rect 16114 31968 16120 31980
rect 16172 31968 16178 32020
rect 18049 32011 18107 32017
rect 18049 31977 18061 32011
rect 18095 32008 18107 32011
rect 18230 32008 18236 32020
rect 18095 31980 18236 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18230 31968 18236 31980
rect 18288 31968 18294 32020
rect 20622 31968 20628 32020
rect 20680 32008 20686 32020
rect 21269 32011 21327 32017
rect 21269 32008 21281 32011
rect 20680 31980 21281 32008
rect 20680 31968 20686 31980
rect 21269 31977 21281 31980
rect 21315 31977 21327 32011
rect 21269 31971 21327 31977
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 23661 32011 23719 32017
rect 23661 32008 23673 32011
rect 23256 31980 23673 32008
rect 23256 31968 23262 31980
rect 23661 31977 23673 31980
rect 23707 31977 23719 32011
rect 23661 31971 23719 31977
rect 8754 31900 8760 31952
rect 8812 31940 8818 31952
rect 9309 31943 9367 31949
rect 9309 31940 9321 31943
rect 8812 31912 9321 31940
rect 8812 31900 8818 31912
rect 9309 31909 9321 31912
rect 9355 31909 9367 31943
rect 9309 31903 9367 31909
rect 11149 31943 11207 31949
rect 11149 31909 11161 31943
rect 11195 31940 11207 31943
rect 11698 31940 11704 31952
rect 11195 31912 11704 31940
rect 11195 31909 11207 31912
rect 11149 31903 11207 31909
rect 11698 31900 11704 31912
rect 11756 31900 11762 31952
rect 15933 31943 15991 31949
rect 15933 31909 15945 31943
rect 15979 31940 15991 31943
rect 16850 31940 16856 31952
rect 15979 31912 16856 31940
rect 15979 31909 15991 31912
rect 15933 31903 15991 31909
rect 16850 31900 16856 31912
rect 16908 31900 16914 31952
rect 18325 31943 18383 31949
rect 18325 31909 18337 31943
rect 18371 31909 18383 31943
rect 18325 31903 18383 31909
rect 8481 31875 8539 31881
rect 8481 31841 8493 31875
rect 8527 31872 8539 31875
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 8527 31844 9781 31872
rect 8527 31841 8539 31844
rect 8481 31835 8539 31841
rect 9769 31841 9781 31844
rect 9815 31841 9827 31875
rect 9769 31835 9827 31841
rect 9858 31832 9864 31884
rect 9916 31872 9922 31884
rect 9916 31844 9961 31872
rect 9916 31832 9922 31844
rect 10502 31832 10508 31884
rect 10560 31872 10566 31884
rect 12621 31875 12679 31881
rect 12621 31872 12633 31875
rect 10560 31844 12633 31872
rect 10560 31832 10566 31844
rect 12621 31841 12633 31844
rect 12667 31841 12679 31875
rect 12621 31835 12679 31841
rect 13541 31875 13599 31881
rect 13541 31841 13553 31875
rect 13587 31872 13599 31875
rect 14369 31875 14427 31881
rect 14369 31872 14381 31875
rect 13587 31844 14381 31872
rect 13587 31841 13599 31844
rect 13541 31835 13599 31841
rect 14369 31841 14381 31844
rect 14415 31841 14427 31875
rect 16393 31875 16451 31881
rect 16393 31872 16405 31875
rect 14369 31835 14427 31841
rect 14660 31844 16405 31872
rect 14660 31816 14688 31844
rect 16393 31841 16405 31844
rect 16439 31841 16451 31875
rect 17126 31872 17132 31884
rect 17087 31844 17132 31872
rect 16393 31835 16451 31841
rect 17126 31832 17132 31844
rect 17184 31832 17190 31884
rect 18340 31872 18368 31903
rect 20530 31900 20536 31952
rect 20588 31940 20594 31952
rect 22462 31940 22468 31952
rect 20588 31912 22048 31940
rect 22375 31912 22468 31940
rect 20588 31900 20594 31912
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 17512 31844 18368 31872
rect 18432 31844 19441 31872
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31804 8447 31807
rect 8435 31776 8524 31804
rect 8435 31773 8447 31776
rect 8389 31767 8447 31773
rect 8496 31736 8524 31776
rect 8570 31764 8576 31816
rect 8628 31804 8634 31816
rect 9677 31807 9735 31813
rect 9677 31804 9689 31807
rect 8628 31776 8673 31804
rect 8772 31776 9689 31804
rect 8628 31764 8634 31776
rect 8772 31736 8800 31776
rect 9677 31773 9689 31776
rect 9723 31804 9735 31807
rect 10134 31804 10140 31816
rect 9723 31776 10140 31804
rect 9723 31773 9735 31776
rect 9677 31767 9735 31773
rect 10134 31764 10140 31776
rect 10192 31764 10198 31816
rect 11422 31804 11428 31816
rect 11383 31776 11428 31804
rect 11422 31764 11428 31776
rect 11480 31764 11486 31816
rect 11701 31807 11759 31813
rect 11701 31773 11713 31807
rect 11747 31804 11759 31807
rect 12342 31804 12348 31816
rect 11747 31776 12348 31804
rect 11747 31773 11759 31776
rect 11701 31767 11759 31773
rect 12342 31764 12348 31776
rect 12400 31764 12406 31816
rect 13449 31807 13507 31813
rect 13449 31773 13461 31807
rect 13495 31804 13507 31807
rect 13998 31804 14004 31816
rect 13495 31776 14004 31804
rect 13495 31773 13507 31776
rect 13449 31767 13507 31773
rect 13998 31764 14004 31776
rect 14056 31764 14062 31816
rect 14274 31804 14280 31816
rect 14235 31776 14280 31804
rect 14274 31764 14280 31776
rect 14332 31764 14338 31816
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 14642 31804 14648 31816
rect 14507 31776 14648 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 14642 31764 14648 31776
rect 14700 31764 14706 31816
rect 16114 31764 16120 31816
rect 16172 31804 16178 31816
rect 17221 31807 17279 31813
rect 17221 31804 17233 31807
rect 16172 31776 16574 31804
rect 16172 31764 16178 31776
rect 8496 31708 8800 31736
rect 10042 31696 10048 31748
rect 10100 31736 10106 31748
rect 15562 31736 15568 31748
rect 10100 31708 15568 31736
rect 10100 31696 10106 31708
rect 15562 31696 15568 31708
rect 15620 31696 15626 31748
rect 16546 31736 16574 31776
rect 16776 31776 17233 31804
rect 16776 31736 16804 31776
rect 17221 31773 17233 31776
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 17310 31764 17316 31816
rect 17368 31804 17374 31816
rect 17368 31776 17413 31804
rect 17368 31764 17374 31776
rect 16546 31708 16804 31736
rect 16853 31739 16911 31745
rect 16853 31705 16865 31739
rect 16899 31736 16911 31739
rect 17512 31736 17540 31844
rect 17862 31764 17868 31816
rect 17920 31804 17926 31816
rect 18325 31807 18383 31813
rect 18325 31804 18337 31807
rect 17920 31776 18337 31804
rect 17920 31764 17926 31776
rect 18325 31773 18337 31776
rect 18371 31804 18383 31807
rect 18432 31804 18460 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 21082 31872 21088 31884
rect 19429 31835 19487 31841
rect 20272 31844 21088 31872
rect 20272 31813 20300 31844
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 22020 31881 22048 31912
rect 22462 31900 22468 31912
rect 22520 31940 22526 31952
rect 24581 31943 24639 31949
rect 24581 31940 24593 31943
rect 22520 31912 24593 31940
rect 22520 31900 22526 31912
rect 24581 31909 24593 31912
rect 24627 31909 24639 31943
rect 24581 31903 24639 31909
rect 22005 31875 22063 31881
rect 22005 31841 22017 31875
rect 22051 31841 22063 31875
rect 22480 31872 22508 31900
rect 22557 31875 22615 31881
rect 22557 31872 22569 31875
rect 22480 31844 22569 31872
rect 22005 31835 22063 31841
rect 22557 31841 22569 31844
rect 22603 31841 22615 31875
rect 23017 31875 23075 31881
rect 23017 31872 23029 31875
rect 22557 31835 22615 31841
rect 22664 31844 23029 31872
rect 18371 31776 18460 31804
rect 18509 31807 18567 31813
rect 18371 31773 18383 31776
rect 18325 31767 18383 31773
rect 18509 31773 18521 31807
rect 18555 31804 18567 31807
rect 20257 31807 20315 31813
rect 18555 31776 20208 31804
rect 18555 31773 18567 31776
rect 18509 31767 18567 31773
rect 16899 31708 17540 31736
rect 16899 31705 16911 31708
rect 16853 31699 16911 31705
rect 8018 31628 8024 31680
rect 8076 31668 8082 31680
rect 11609 31671 11667 31677
rect 11609 31668 11621 31671
rect 8076 31640 11621 31668
rect 8076 31628 8082 31640
rect 11609 31637 11621 31640
rect 11655 31637 11667 31671
rect 11609 31631 11667 31637
rect 15746 31628 15752 31680
rect 15804 31677 15810 31680
rect 15804 31671 15823 31677
rect 15811 31637 15823 31671
rect 20180 31668 20208 31776
rect 20257 31773 20269 31807
rect 20303 31773 20315 31807
rect 20257 31767 20315 31773
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31804 20499 31807
rect 20806 31804 20812 31816
rect 20487 31776 20812 31804
rect 20487 31773 20499 31776
rect 20441 31767 20499 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 20993 31807 21051 31813
rect 20993 31773 21005 31807
rect 21039 31804 21051 31807
rect 21174 31804 21180 31816
rect 21039 31776 21180 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 21174 31764 21180 31776
rect 21232 31764 21238 31816
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31804 21327 31807
rect 21358 31804 21364 31816
rect 21315 31776 21364 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 21358 31764 21364 31776
rect 21416 31764 21422 31816
rect 22664 31804 22692 31844
rect 23017 31841 23029 31844
rect 23063 31841 23075 31875
rect 25038 31872 25044 31884
rect 24999 31844 25044 31872
rect 23017 31835 23075 31841
rect 25038 31832 25044 31844
rect 25096 31832 25102 31884
rect 25130 31832 25136 31884
rect 25188 31872 25194 31884
rect 25188 31844 25233 31872
rect 25188 31832 25194 31844
rect 22830 31804 22836 31816
rect 21468 31776 22692 31804
rect 22791 31776 22836 31804
rect 21082 31736 21088 31748
rect 21043 31708 21088 31736
rect 21082 31696 21088 31708
rect 21140 31696 21146 31748
rect 21468 31668 21496 31776
rect 20180 31640 21496 31668
rect 22664 31668 22692 31776
rect 22830 31764 22836 31776
rect 22888 31764 22894 31816
rect 23658 31804 23664 31816
rect 23619 31776 23664 31804
rect 23658 31764 23664 31776
rect 23716 31764 23722 31816
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 26421 31807 26479 31813
rect 26421 31773 26433 31807
rect 26467 31773 26479 31807
rect 26602 31804 26608 31816
rect 26563 31776 26608 31804
rect 26421 31767 26479 31773
rect 23382 31696 23388 31748
rect 23440 31736 23446 31748
rect 23860 31736 23888 31767
rect 23440 31708 23888 31736
rect 26436 31736 26464 31767
rect 26602 31764 26608 31776
rect 26660 31764 26666 31816
rect 26694 31736 26700 31748
rect 26436 31708 26700 31736
rect 23440 31696 23446 31708
rect 26694 31696 26700 31708
rect 26752 31696 26758 31748
rect 27706 31736 27712 31748
rect 27554 31708 27712 31736
rect 27706 31696 27712 31708
rect 27764 31696 27770 31748
rect 22738 31668 22744 31680
rect 22664 31640 22744 31668
rect 15804 31631 15823 31637
rect 15804 31628 15810 31631
rect 22738 31628 22744 31640
rect 22796 31628 22802 31680
rect 23474 31668 23480 31680
rect 23435 31640 23480 31668
rect 23474 31628 23480 31640
rect 23532 31628 23538 31680
rect 24762 31628 24768 31680
rect 24820 31668 24826 31680
rect 24949 31671 25007 31677
rect 24949 31668 24961 31671
rect 24820 31640 24961 31668
rect 24820 31628 24826 31640
rect 24949 31637 24961 31640
rect 24995 31637 25007 31671
rect 24949 31631 25007 31637
rect 1104 31578 35027 31600
rect 1104 31526 9390 31578
rect 9442 31526 9454 31578
rect 9506 31526 9518 31578
rect 9570 31526 9582 31578
rect 9634 31526 9646 31578
rect 9698 31526 17831 31578
rect 17883 31526 17895 31578
rect 17947 31526 17959 31578
rect 18011 31526 18023 31578
rect 18075 31526 18087 31578
rect 18139 31526 26272 31578
rect 26324 31526 26336 31578
rect 26388 31526 26400 31578
rect 26452 31526 26464 31578
rect 26516 31526 26528 31578
rect 26580 31526 34713 31578
rect 34765 31526 34777 31578
rect 34829 31526 34841 31578
rect 34893 31526 34905 31578
rect 34957 31526 34969 31578
rect 35021 31526 35027 31578
rect 1104 31504 35027 31526
rect 9493 31467 9551 31473
rect 9493 31433 9505 31467
rect 9539 31464 9551 31467
rect 9858 31464 9864 31476
rect 9539 31436 9864 31464
rect 9539 31433 9551 31436
rect 9493 31427 9551 31433
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 13541 31467 13599 31473
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 14274 31464 14280 31476
rect 13587 31436 14280 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 14274 31424 14280 31436
rect 14332 31424 14338 31476
rect 16114 31464 16120 31476
rect 16075 31436 16120 31464
rect 16114 31424 16120 31436
rect 16172 31464 16178 31476
rect 17037 31467 17095 31473
rect 17037 31464 17049 31467
rect 16172 31436 17049 31464
rect 16172 31424 16178 31436
rect 17037 31433 17049 31436
rect 17083 31433 17095 31467
rect 17037 31427 17095 31433
rect 17310 31424 17316 31476
rect 17368 31464 17374 31476
rect 17589 31467 17647 31473
rect 17589 31464 17601 31467
rect 17368 31436 17601 31464
rect 17368 31424 17374 31436
rect 17589 31433 17601 31436
rect 17635 31433 17647 31467
rect 17589 31427 17647 31433
rect 20806 31424 20812 31476
rect 20864 31473 20870 31476
rect 20864 31467 20892 31473
rect 20880 31433 20892 31467
rect 20864 31427 20892 31433
rect 24765 31467 24823 31473
rect 24765 31433 24777 31467
rect 24811 31464 24823 31467
rect 25130 31464 25136 31476
rect 24811 31436 25136 31464
rect 24811 31433 24823 31436
rect 24765 31427 24823 31433
rect 20864 31424 20870 31427
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 25222 31424 25228 31476
rect 25280 31464 25286 31476
rect 25774 31464 25780 31476
rect 25280 31436 25780 31464
rect 25280 31424 25286 31436
rect 25774 31424 25780 31436
rect 25832 31424 25838 31476
rect 25869 31467 25927 31473
rect 25869 31433 25881 31467
rect 25915 31464 25927 31467
rect 26602 31464 26608 31476
rect 25915 31436 26608 31464
rect 25915 31433 25927 31436
rect 25869 31427 25927 31433
rect 26602 31424 26608 31436
rect 26660 31424 26666 31476
rect 28629 31467 28687 31473
rect 28629 31464 28641 31467
rect 27356 31436 28641 31464
rect 9766 31396 9772 31408
rect 9140 31368 9772 31396
rect 9140 31337 9168 31368
rect 9766 31356 9772 31368
rect 9824 31396 9830 31408
rect 10042 31396 10048 31408
rect 9824 31368 10048 31396
rect 9824 31356 9830 31368
rect 10042 31356 10048 31368
rect 10100 31356 10106 31408
rect 10594 31356 10600 31408
rect 10652 31396 10658 31408
rect 10689 31399 10747 31405
rect 10689 31396 10701 31399
rect 10652 31368 10701 31396
rect 10652 31356 10658 31368
rect 10689 31365 10701 31368
rect 10735 31365 10747 31399
rect 10689 31359 10747 31365
rect 13188 31368 15516 31396
rect 9125 31331 9183 31337
rect 9125 31297 9137 31331
rect 9171 31297 9183 31331
rect 10226 31328 10232 31340
rect 10187 31300 10232 31328
rect 9125 31291 9183 31297
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 10321 31331 10379 31337
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10321 31291 10379 31297
rect 9217 31263 9275 31269
rect 9217 31229 9229 31263
rect 9263 31260 9275 31263
rect 9398 31260 9404 31272
rect 9263 31232 9404 31260
rect 9263 31229 9275 31232
rect 9217 31223 9275 31229
rect 9398 31220 9404 31232
rect 9456 31220 9462 31272
rect 10042 31220 10048 31272
rect 10100 31260 10106 31272
rect 10336 31260 10364 31291
rect 12618 31288 12624 31340
rect 12676 31328 12682 31340
rect 13188 31337 13216 31368
rect 15488 31340 15516 31368
rect 15562 31356 15568 31408
rect 15620 31396 15626 31408
rect 16853 31399 16911 31405
rect 16853 31396 16865 31399
rect 15620 31368 16865 31396
rect 15620 31356 15626 31368
rect 16853 31365 16865 31368
rect 16899 31396 16911 31399
rect 19334 31396 19340 31408
rect 16899 31368 19340 31396
rect 16899 31365 16911 31368
rect 16853 31359 16911 31365
rect 19334 31356 19340 31368
rect 19392 31356 19398 31408
rect 22189 31399 22247 31405
rect 22189 31396 22201 31399
rect 20640 31368 22201 31396
rect 13173 31331 13231 31337
rect 13173 31328 13185 31331
rect 12676 31300 13185 31328
rect 12676 31288 12682 31300
rect 13173 31297 13185 31300
rect 13219 31297 13231 31331
rect 14090 31328 14096 31340
rect 14051 31300 14096 31328
rect 13173 31291 13231 31297
rect 14090 31288 14096 31300
rect 14148 31288 14154 31340
rect 14826 31328 14832 31340
rect 14787 31300 14832 31328
rect 14826 31288 14832 31300
rect 14884 31288 14890 31340
rect 14921 31331 14979 31337
rect 14921 31297 14933 31331
rect 14967 31297 14979 31331
rect 14921 31291 14979 31297
rect 10100 31232 10364 31260
rect 10413 31263 10471 31269
rect 10100 31220 10106 31232
rect 10413 31229 10425 31263
rect 10459 31260 10471 31263
rect 10594 31260 10600 31272
rect 10459 31232 10600 31260
rect 10459 31229 10471 31232
rect 10413 31223 10471 31229
rect 10594 31220 10600 31232
rect 10652 31220 10658 31272
rect 13262 31260 13268 31272
rect 13223 31232 13268 31260
rect 13262 31220 13268 31232
rect 13320 31220 13326 31272
rect 13924 31232 14412 31260
rect 10686 31152 10692 31204
rect 10744 31192 10750 31204
rect 10873 31195 10931 31201
rect 10873 31192 10885 31195
rect 10744 31164 10885 31192
rect 10744 31152 10750 31164
rect 10873 31161 10885 31164
rect 10919 31161 10931 31195
rect 13924 31192 13952 31232
rect 10873 31155 10931 31161
rect 12406 31164 13952 31192
rect 10318 31084 10324 31136
rect 10376 31124 10382 31136
rect 12406 31124 12434 31164
rect 14274 31124 14280 31136
rect 10376 31096 12434 31124
rect 14235 31096 14280 31124
rect 10376 31084 10382 31096
rect 14274 31084 14280 31096
rect 14332 31084 14338 31136
rect 14384 31124 14412 31232
rect 14642 31220 14648 31272
rect 14700 31260 14706 31272
rect 14936 31260 14964 31291
rect 15470 31288 15476 31340
rect 15528 31328 15534 31340
rect 16117 31331 16175 31337
rect 16117 31328 16129 31331
rect 15528 31300 16129 31328
rect 15528 31288 15534 31300
rect 16117 31297 16129 31300
rect 16163 31297 16175 31331
rect 16298 31328 16304 31340
rect 16259 31300 16304 31328
rect 16117 31291 16175 31297
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 17126 31328 17132 31340
rect 17039 31300 17132 31328
rect 17126 31288 17132 31300
rect 17184 31288 17190 31340
rect 17589 31331 17647 31337
rect 17589 31297 17601 31331
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 14700 31232 14964 31260
rect 14700 31220 14706 31232
rect 15746 31220 15752 31272
rect 15804 31260 15810 31272
rect 17144 31260 17172 31288
rect 15804 31232 17172 31260
rect 17604 31260 17632 31291
rect 17678 31288 17684 31340
rect 17736 31328 17742 31340
rect 17773 31331 17831 31337
rect 17773 31328 17785 31331
rect 17736 31300 17785 31328
rect 17736 31288 17742 31300
rect 17773 31297 17785 31300
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 20346 31288 20352 31340
rect 20404 31328 20410 31340
rect 20640 31337 20668 31368
rect 22189 31365 22201 31368
rect 22235 31365 22247 31399
rect 27157 31399 27215 31405
rect 27157 31396 27169 31399
rect 22189 31359 22247 31365
rect 24596 31368 27169 31396
rect 20625 31331 20683 31337
rect 20625 31328 20637 31331
rect 20404 31300 20637 31328
rect 20404 31288 20410 31300
rect 20625 31297 20637 31300
rect 20671 31297 20683 31331
rect 20625 31291 20683 31297
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 21048 31300 21097 31328
rect 21048 31288 21054 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 22646 31328 22652 31340
rect 22607 31300 22652 31328
rect 21085 31291 21143 31297
rect 22646 31288 22652 31300
rect 22704 31288 22710 31340
rect 22738 31288 22744 31340
rect 22796 31328 22802 31340
rect 23014 31328 23020 31340
rect 22796 31300 22841 31328
rect 22975 31300 23020 31328
rect 22796 31288 22802 31300
rect 23014 31288 23020 31300
rect 23072 31288 23078 31340
rect 23293 31331 23351 31337
rect 23293 31297 23305 31331
rect 23339 31297 23351 31331
rect 23474 31328 23480 31340
rect 23435 31300 23480 31328
rect 23293 31291 23351 31297
rect 21364 31272 21416 31278
rect 20530 31260 20536 31272
rect 17604 31232 17724 31260
rect 20491 31232 20536 31260
rect 15804 31220 15810 31232
rect 17696 31192 17724 31232
rect 20530 31220 20536 31232
rect 20588 31220 20594 31272
rect 21450 31220 21456 31272
rect 21508 31260 21514 31272
rect 23308 31260 23336 31291
rect 23474 31288 23480 31300
rect 23532 31288 23538 31340
rect 24213 31331 24271 31337
rect 24213 31297 24225 31331
rect 24259 31328 24271 31331
rect 24486 31328 24492 31340
rect 24259 31300 24492 31328
rect 24259 31297 24271 31300
rect 24213 31291 24271 31297
rect 24486 31288 24492 31300
rect 24544 31288 24550 31340
rect 24596 31337 24624 31368
rect 25608 31340 25636 31368
rect 27157 31365 27169 31368
rect 27203 31365 27215 31399
rect 27157 31359 27215 31365
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 25222 31328 25228 31340
rect 24581 31291 24639 31297
rect 24688 31300 25228 31328
rect 21508 31232 23336 31260
rect 21508 31220 21514 31232
rect 23658 31220 23664 31272
rect 23716 31260 23722 31272
rect 24688 31260 24716 31300
rect 25222 31288 25228 31300
rect 25280 31288 25286 31340
rect 25314 31288 25320 31340
rect 25372 31328 25378 31340
rect 25409 31331 25467 31337
rect 25409 31328 25421 31331
rect 25372 31300 25421 31328
rect 25372 31288 25378 31300
rect 25409 31297 25421 31300
rect 25455 31297 25467 31331
rect 25590 31328 25596 31340
rect 25503 31300 25596 31328
rect 25409 31291 25467 31297
rect 25590 31288 25596 31300
rect 25648 31288 25654 31340
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31297 25743 31331
rect 25685 31291 25743 31297
rect 23716 31232 24716 31260
rect 23716 31220 23722 31232
rect 25038 31220 25044 31272
rect 25096 31260 25102 31272
rect 25700 31260 25728 31291
rect 26694 31288 26700 31340
rect 26752 31328 26758 31340
rect 27356 31337 27384 31436
rect 28629 31433 28641 31436
rect 28675 31433 28687 31467
rect 28629 31427 28687 31433
rect 27341 31331 27399 31337
rect 27341 31328 27353 31331
rect 26752 31300 27353 31328
rect 26752 31288 26758 31300
rect 27341 31297 27353 31300
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 27893 31331 27951 31337
rect 27893 31297 27905 31331
rect 27939 31328 27951 31331
rect 28567 31331 28625 31337
rect 28567 31328 28579 31331
rect 27939 31300 28579 31328
rect 27939 31297 27951 31300
rect 27893 31291 27951 31297
rect 28567 31297 28579 31300
rect 28613 31297 28625 31331
rect 28567 31291 28625 31297
rect 25096 31232 25728 31260
rect 25096 31220 25102 31232
rect 25774 31220 25780 31272
rect 25832 31260 25838 31272
rect 27908 31260 27936 31291
rect 29086 31260 29092 31272
rect 25832 31232 27936 31260
rect 29047 31232 29092 31260
rect 25832 31220 25838 31232
rect 29086 31220 29092 31232
rect 29144 31220 29150 31272
rect 21364 31214 21416 31220
rect 16408 31164 17724 31192
rect 16408 31124 16436 31164
rect 14384 31096 16436 31124
rect 16853 31127 16911 31133
rect 16853 31093 16865 31127
rect 16899 31124 16911 31127
rect 17034 31124 17040 31136
rect 16899 31096 17040 31124
rect 16899 31093 16911 31096
rect 16853 31087 16911 31093
rect 17034 31084 17040 31096
rect 17092 31084 17098 31136
rect 17696 31124 17724 31164
rect 25501 31195 25559 31201
rect 25501 31161 25513 31195
rect 25547 31161 25559 31195
rect 25501 31155 25559 31161
rect 21910 31124 21916 31136
rect 17696 31096 21916 31124
rect 21910 31084 21916 31096
rect 21968 31084 21974 31136
rect 24581 31127 24639 31133
rect 24581 31093 24593 31127
rect 24627 31124 24639 31127
rect 25516 31124 25544 31155
rect 26050 31124 26056 31136
rect 24627 31096 26056 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 26050 31084 26056 31096
rect 26108 31124 26114 31136
rect 28445 31127 28503 31133
rect 28445 31124 28457 31127
rect 26108 31096 28457 31124
rect 26108 31084 26114 31096
rect 28445 31093 28457 31096
rect 28491 31093 28503 31127
rect 28445 31087 28503 31093
rect 28534 31084 28540 31136
rect 28592 31124 28598 31136
rect 28997 31127 29055 31133
rect 28997 31124 29009 31127
rect 28592 31096 29009 31124
rect 28592 31084 28598 31096
rect 28997 31093 29009 31096
rect 29043 31093 29055 31127
rect 28997 31087 29055 31093
rect 1104 31034 34868 31056
rect 1104 30982 5170 31034
rect 5222 30982 5234 31034
rect 5286 30982 5298 31034
rect 5350 30982 5362 31034
rect 5414 30982 5426 31034
rect 5478 30982 13611 31034
rect 13663 30982 13675 31034
rect 13727 30982 13739 31034
rect 13791 30982 13803 31034
rect 13855 30982 13867 31034
rect 13919 30982 22052 31034
rect 22104 30982 22116 31034
rect 22168 30982 22180 31034
rect 22232 30982 22244 31034
rect 22296 30982 22308 31034
rect 22360 30982 30493 31034
rect 30545 30982 30557 31034
rect 30609 30982 30621 31034
rect 30673 30982 30685 31034
rect 30737 30982 30749 31034
rect 30801 30982 34868 31034
rect 1104 30960 34868 30982
rect 9398 30920 9404 30932
rect 9359 30892 9404 30920
rect 9398 30880 9404 30892
rect 9456 30880 9462 30932
rect 10042 30920 10048 30932
rect 10003 30892 10048 30920
rect 10042 30880 10048 30892
rect 10100 30880 10106 30932
rect 10226 30880 10232 30932
rect 10284 30920 10290 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10284 30892 10701 30920
rect 10284 30880 10290 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 13262 30880 13268 30932
rect 13320 30920 13326 30932
rect 13541 30923 13599 30929
rect 13541 30920 13553 30923
rect 13320 30892 13553 30920
rect 13320 30880 13326 30892
rect 13541 30889 13553 30892
rect 13587 30889 13599 30923
rect 13541 30883 13599 30889
rect 17037 30923 17095 30929
rect 17037 30889 17049 30923
rect 17083 30920 17095 30923
rect 17402 30920 17408 30932
rect 17083 30892 17408 30920
rect 17083 30889 17095 30892
rect 17037 30883 17095 30889
rect 17402 30880 17408 30892
rect 17460 30880 17466 30932
rect 20990 30920 20996 30932
rect 20951 30892 20996 30920
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 22741 30923 22799 30929
rect 22741 30889 22753 30923
rect 22787 30920 22799 30923
rect 23014 30920 23020 30932
rect 22787 30892 23020 30920
rect 22787 30889 22799 30892
rect 22741 30883 22799 30889
rect 23014 30880 23020 30892
rect 23072 30880 23078 30932
rect 10060 30784 10088 30880
rect 14826 30812 14832 30864
rect 14884 30852 14890 30864
rect 23109 30855 23167 30861
rect 14884 30824 16160 30852
rect 14884 30812 14890 30824
rect 9324 30756 10088 30784
rect 9324 30725 9352 30756
rect 10502 30744 10508 30796
rect 10560 30784 10566 30796
rect 13449 30787 13507 30793
rect 10560 30756 10824 30784
rect 10560 30744 10566 30756
rect 9309 30719 9367 30725
rect 9309 30685 9321 30719
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 9493 30719 9551 30725
rect 9493 30685 9505 30719
rect 9539 30685 9551 30719
rect 9950 30716 9956 30728
rect 9911 30688 9956 30716
rect 9493 30679 9551 30685
rect 9508 30648 9536 30679
rect 9950 30676 9956 30688
rect 10008 30676 10014 30728
rect 10134 30716 10140 30728
rect 10095 30688 10140 30716
rect 10134 30676 10140 30688
rect 10192 30676 10198 30728
rect 10318 30676 10324 30728
rect 10376 30716 10382 30728
rect 10796 30725 10824 30756
rect 13449 30753 13461 30787
rect 13495 30784 13507 30787
rect 14844 30784 14872 30812
rect 15746 30784 15752 30796
rect 13495 30756 14872 30784
rect 15707 30756 15752 30784
rect 13495 30753 13507 30756
rect 13449 30747 13507 30753
rect 15746 30744 15752 30756
rect 15804 30744 15810 30796
rect 10597 30719 10655 30725
rect 10597 30716 10609 30719
rect 10376 30688 10609 30716
rect 10376 30676 10382 30688
rect 10597 30685 10609 30688
rect 10643 30685 10655 30719
rect 10597 30679 10655 30685
rect 10781 30719 10839 30725
rect 10781 30685 10793 30719
rect 10827 30685 10839 30719
rect 10781 30679 10839 30685
rect 13633 30719 13691 30725
rect 13633 30685 13645 30719
rect 13679 30685 13691 30719
rect 13633 30679 13691 30685
rect 13725 30719 13783 30725
rect 13725 30685 13737 30719
rect 13771 30716 13783 30719
rect 14090 30716 14096 30728
rect 13771 30688 14096 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 13648 30648 13676 30679
rect 14090 30676 14096 30688
rect 14148 30716 14154 30728
rect 14550 30716 14556 30728
rect 14148 30688 14556 30716
rect 14148 30676 14154 30688
rect 14550 30676 14556 30688
rect 14608 30676 14614 30728
rect 14918 30716 14924 30728
rect 14879 30688 14924 30716
rect 14918 30676 14924 30688
rect 14976 30676 14982 30728
rect 15470 30716 15476 30728
rect 15431 30688 15476 30716
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 16132 30725 16160 30824
rect 23109 30821 23121 30855
rect 23155 30852 23167 30855
rect 23382 30852 23388 30864
rect 23155 30824 23388 30852
rect 23155 30821 23167 30824
rect 23109 30815 23167 30821
rect 23382 30812 23388 30824
rect 23440 30852 23446 30864
rect 27525 30855 27583 30861
rect 27525 30852 27537 30855
rect 23440 30824 27537 30852
rect 23440 30812 23446 30824
rect 27525 30821 27537 30824
rect 27571 30821 27583 30855
rect 27525 30815 27583 30821
rect 23658 30784 23664 30796
rect 22940 30756 23664 30784
rect 15933 30719 15991 30725
rect 15933 30685 15945 30719
rect 15979 30685 15991 30719
rect 15933 30679 15991 30685
rect 16117 30719 16175 30725
rect 16117 30685 16129 30719
rect 16163 30685 16175 30719
rect 16850 30716 16856 30728
rect 16811 30688 16856 30716
rect 16117 30679 16175 30685
rect 14936 30648 14964 30676
rect 9508 30620 10640 30648
rect 13648 30620 14964 30648
rect 15948 30648 15976 30679
rect 16850 30676 16856 30688
rect 16908 30676 16914 30728
rect 17034 30716 17040 30728
rect 16995 30688 17040 30716
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 20717 30719 20775 30725
rect 20717 30685 20729 30719
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 20809 30719 20867 30725
rect 20809 30685 20821 30719
rect 20855 30716 20867 30719
rect 21450 30716 21456 30728
rect 20855 30688 21456 30716
rect 20855 30685 20867 30688
rect 20809 30679 20867 30685
rect 16298 30648 16304 30660
rect 15948 30620 16304 30648
rect 10612 30592 10640 30620
rect 10594 30540 10600 30592
rect 10652 30540 10658 30592
rect 13998 30540 14004 30592
rect 14056 30580 14062 30592
rect 15948 30580 15976 30620
rect 16298 30608 16304 30620
rect 16356 30648 16362 30660
rect 18782 30648 18788 30660
rect 16356 30620 18788 30648
rect 16356 30608 16362 30620
rect 18782 30608 18788 30620
rect 18840 30608 18846 30660
rect 20732 30648 20760 30679
rect 21450 30676 21456 30688
rect 21508 30676 21514 30728
rect 22940 30725 22968 30756
rect 23658 30744 23664 30756
rect 23716 30744 23722 30796
rect 25222 30744 25228 30796
rect 25280 30784 25286 30796
rect 29086 30784 29092 30796
rect 25280 30756 26280 30784
rect 25280 30744 25286 30756
rect 22925 30719 22983 30725
rect 22925 30716 22937 30719
rect 22066 30688 22937 30716
rect 22066 30648 22094 30688
rect 22925 30685 22937 30688
rect 22971 30685 22983 30719
rect 23198 30716 23204 30728
rect 23159 30688 23204 30716
rect 22925 30679 22983 30685
rect 23198 30676 23204 30688
rect 23256 30676 23262 30728
rect 25038 30716 25044 30728
rect 24999 30688 25044 30716
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 25590 30716 25596 30728
rect 25551 30688 25596 30716
rect 25590 30676 25596 30688
rect 25648 30676 25654 30728
rect 26050 30716 26056 30728
rect 26011 30688 26056 30716
rect 26050 30676 26056 30688
rect 26108 30676 26114 30728
rect 26252 30725 26280 30756
rect 28460 30756 29092 30784
rect 28460 30725 28488 30756
rect 29086 30744 29092 30756
rect 29144 30744 29150 30796
rect 26237 30719 26295 30725
rect 26237 30685 26249 30719
rect 26283 30685 26295 30719
rect 27709 30719 27767 30725
rect 27709 30716 27721 30719
rect 26237 30679 26295 30685
rect 26988 30688 27721 30716
rect 26988 30660 27016 30688
rect 27709 30685 27721 30688
rect 27755 30685 27767 30719
rect 27709 30679 27767 30685
rect 28077 30719 28135 30725
rect 28077 30685 28089 30719
rect 28123 30685 28135 30719
rect 28077 30679 28135 30685
rect 28445 30719 28503 30725
rect 28445 30685 28457 30719
rect 28491 30685 28503 30719
rect 28902 30716 28908 30728
rect 28863 30688 28908 30716
rect 28445 30679 28503 30685
rect 20732 30620 22094 30648
rect 26145 30651 26203 30657
rect 26145 30617 26157 30651
rect 26191 30648 26203 30651
rect 26970 30648 26976 30660
rect 26191 30620 26976 30648
rect 26191 30617 26203 30620
rect 26145 30611 26203 30617
rect 26970 30608 26976 30620
rect 27028 30608 27034 30660
rect 27614 30608 27620 30660
rect 27672 30648 27678 30660
rect 28092 30648 28120 30679
rect 28902 30676 28908 30688
rect 28960 30676 28966 30728
rect 28718 30648 28724 30660
rect 27672 30620 28724 30648
rect 27672 30608 27678 30620
rect 28718 30608 28724 30620
rect 28776 30608 28782 30660
rect 14056 30552 15976 30580
rect 14056 30540 14062 30552
rect 1104 30490 35027 30512
rect 1104 30438 9390 30490
rect 9442 30438 9454 30490
rect 9506 30438 9518 30490
rect 9570 30438 9582 30490
rect 9634 30438 9646 30490
rect 9698 30438 17831 30490
rect 17883 30438 17895 30490
rect 17947 30438 17959 30490
rect 18011 30438 18023 30490
rect 18075 30438 18087 30490
rect 18139 30438 26272 30490
rect 26324 30438 26336 30490
rect 26388 30438 26400 30490
rect 26452 30438 26464 30490
rect 26516 30438 26528 30490
rect 26580 30438 34713 30490
rect 34765 30438 34777 30490
rect 34829 30438 34841 30490
rect 34893 30438 34905 30490
rect 34957 30438 34969 30490
rect 35021 30438 35027 30490
rect 1104 30416 35027 30438
rect 26050 30376 26056 30388
rect 25608 30348 26056 30376
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 14274 30240 14280 30252
rect 14235 30212 14280 30240
rect 14274 30200 14280 30212
rect 14332 30200 14338 30252
rect 14918 30240 14924 30252
rect 14879 30212 14924 30240
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30240 19763 30243
rect 20162 30240 20168 30252
rect 19751 30212 20168 30240
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20806 30240 20812 30252
rect 20303 30212 20812 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 20898 30200 20904 30252
rect 20956 30240 20962 30252
rect 20993 30243 21051 30249
rect 20993 30240 21005 30243
rect 20956 30212 21005 30240
rect 20956 30200 20962 30212
rect 20993 30209 21005 30212
rect 21039 30209 21051 30243
rect 24670 30240 24676 30252
rect 24631 30212 24676 30240
rect 20993 30203 21051 30209
rect 24670 30200 24676 30212
rect 24728 30200 24734 30252
rect 25130 30240 25136 30252
rect 25091 30212 25136 30240
rect 25130 30200 25136 30212
rect 25188 30200 25194 30252
rect 25222 30200 25228 30252
rect 25280 30240 25286 30252
rect 25608 30249 25636 30348
rect 26050 30336 26056 30348
rect 26108 30336 26114 30388
rect 29086 30376 29092 30388
rect 27632 30348 29092 30376
rect 25317 30243 25375 30249
rect 25317 30240 25329 30243
rect 25280 30212 25329 30240
rect 25280 30200 25286 30212
rect 25317 30209 25329 30212
rect 25363 30209 25375 30243
rect 25317 30203 25375 30209
rect 25593 30243 25651 30249
rect 25593 30209 25605 30243
rect 25639 30209 25651 30243
rect 25593 30203 25651 30209
rect 25682 30200 25688 30252
rect 25740 30240 25746 30252
rect 25869 30243 25927 30249
rect 25869 30240 25881 30243
rect 25740 30212 25881 30240
rect 25740 30200 25746 30212
rect 25869 30209 25881 30212
rect 25915 30209 25927 30243
rect 25869 30203 25927 30209
rect 26053 30243 26111 30249
rect 26053 30209 26065 30243
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 25038 30132 25044 30184
rect 25096 30172 25102 30184
rect 26068 30172 26096 30203
rect 26970 30200 26976 30252
rect 27028 30240 27034 30252
rect 27341 30243 27399 30249
rect 27341 30240 27353 30243
rect 27028 30212 27353 30240
rect 27028 30200 27034 30212
rect 27341 30209 27353 30212
rect 27387 30209 27399 30243
rect 27341 30203 27399 30209
rect 27522 30200 27528 30252
rect 27580 30240 27586 30252
rect 27632 30249 27660 30348
rect 29086 30336 29092 30348
rect 29144 30376 29150 30388
rect 29733 30379 29791 30385
rect 29733 30376 29745 30379
rect 29144 30348 29745 30376
rect 29144 30336 29150 30348
rect 29733 30345 29745 30348
rect 29779 30345 29791 30379
rect 29733 30339 29791 30345
rect 28074 30308 28080 30320
rect 28035 30280 28080 30308
rect 28074 30268 28080 30280
rect 28132 30268 28138 30320
rect 28534 30308 28540 30320
rect 28495 30280 28540 30308
rect 28534 30268 28540 30280
rect 28592 30268 28598 30320
rect 27617 30243 27675 30249
rect 27617 30240 27629 30243
rect 27580 30212 27629 30240
rect 27580 30200 27586 30212
rect 27617 30209 27629 30212
rect 27663 30209 27675 30243
rect 27617 30203 27675 30209
rect 25096 30144 26096 30172
rect 27433 30175 27491 30181
rect 25096 30132 25102 30144
rect 27433 30141 27445 30175
rect 27479 30172 27491 30175
rect 28552 30172 28580 30268
rect 28718 30240 28724 30252
rect 28679 30212 28724 30240
rect 28718 30200 28724 30212
rect 28776 30200 28782 30252
rect 28994 30240 29000 30252
rect 28955 30212 29000 30240
rect 28994 30200 29000 30212
rect 29052 30200 29058 30252
rect 29178 30240 29184 30252
rect 29139 30212 29184 30240
rect 29178 30200 29184 30212
rect 29236 30200 29242 30252
rect 29641 30243 29699 30249
rect 29641 30209 29653 30243
rect 29687 30209 29699 30243
rect 29641 30203 29699 30209
rect 29825 30243 29883 30249
rect 29825 30209 29837 30243
rect 29871 30209 29883 30243
rect 29825 30203 29883 30209
rect 27479 30144 28580 30172
rect 27479 30141 27491 30144
rect 27433 30135 27491 30141
rect 28626 30132 28632 30184
rect 28684 30172 28690 30184
rect 29656 30172 29684 30203
rect 28684 30144 29684 30172
rect 28684 30132 28690 30144
rect 28074 30064 28080 30116
rect 28132 30104 28138 30116
rect 29840 30104 29868 30203
rect 28132 30076 29868 30104
rect 28132 30064 28138 30076
rect 12894 29996 12900 30048
rect 12952 30036 12958 30048
rect 13449 30039 13507 30045
rect 13449 30036 13461 30039
rect 12952 30008 13461 30036
rect 12952 29996 12958 30008
rect 13449 30005 13461 30008
rect 13495 30005 13507 30039
rect 13449 29999 13507 30005
rect 20622 29996 20628 30048
rect 20680 30036 20686 30048
rect 20901 30039 20959 30045
rect 20901 30036 20913 30039
rect 20680 30008 20913 30036
rect 20680 29996 20686 30008
rect 20901 30005 20913 30008
rect 20947 30005 20959 30039
rect 20901 29999 20959 30005
rect 27430 29996 27436 30048
rect 27488 30036 27494 30048
rect 28626 30036 28632 30048
rect 27488 30008 28632 30036
rect 27488 29996 27494 30008
rect 28626 29996 28632 30008
rect 28684 29996 28690 30048
rect 1104 29946 34868 29968
rect 1104 29894 5170 29946
rect 5222 29894 5234 29946
rect 5286 29894 5298 29946
rect 5350 29894 5362 29946
rect 5414 29894 5426 29946
rect 5478 29894 13611 29946
rect 13663 29894 13675 29946
rect 13727 29894 13739 29946
rect 13791 29894 13803 29946
rect 13855 29894 13867 29946
rect 13919 29894 22052 29946
rect 22104 29894 22116 29946
rect 22168 29894 22180 29946
rect 22232 29894 22244 29946
rect 22296 29894 22308 29946
rect 22360 29894 30493 29946
rect 30545 29894 30557 29946
rect 30609 29894 30621 29946
rect 30673 29894 30685 29946
rect 30737 29894 30749 29946
rect 30801 29894 34868 29946
rect 1104 29872 34868 29894
rect 14826 29832 14832 29844
rect 14787 29804 14832 29832
rect 14826 29792 14832 29804
rect 14884 29792 14890 29844
rect 25038 29832 25044 29844
rect 24999 29804 25044 29832
rect 25038 29792 25044 29804
rect 25096 29792 25102 29844
rect 25130 29792 25136 29844
rect 25188 29832 25194 29844
rect 25188 29804 28580 29832
rect 25188 29792 25194 29804
rect 9030 29724 9036 29776
rect 9088 29764 9094 29776
rect 10413 29767 10471 29773
rect 10413 29764 10425 29767
rect 9088 29736 10425 29764
rect 9088 29724 9094 29736
rect 10413 29733 10425 29736
rect 10459 29733 10471 29767
rect 10413 29727 10471 29733
rect 19720 29736 22094 29764
rect 10686 29696 10692 29708
rect 9968 29668 10692 29696
rect 9968 29637 9996 29668
rect 10686 29656 10692 29668
rect 10744 29656 10750 29708
rect 9677 29631 9735 29637
rect 9677 29597 9689 29631
rect 9723 29597 9735 29631
rect 9677 29591 9735 29597
rect 9953 29631 10011 29637
rect 9953 29597 9965 29631
rect 9999 29597 10011 29631
rect 10410 29628 10416 29640
rect 10371 29600 10416 29628
rect 9953 29591 10011 29597
rect 9692 29560 9720 29591
rect 10410 29588 10416 29600
rect 10468 29588 10474 29640
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 12894 29628 12900 29640
rect 10551 29600 12900 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 10134 29560 10140 29572
rect 9692 29532 10140 29560
rect 10134 29520 10140 29532
rect 10192 29560 10198 29572
rect 10520 29560 10548 29591
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 12989 29631 13047 29637
rect 12989 29597 13001 29631
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 13173 29631 13231 29637
rect 13173 29597 13185 29631
rect 13219 29628 13231 29631
rect 14921 29631 14979 29637
rect 14921 29628 14933 29631
rect 13219 29600 14933 29628
rect 13219 29597 13231 29600
rect 13173 29591 13231 29597
rect 14921 29597 14933 29600
rect 14967 29628 14979 29631
rect 15010 29628 15016 29640
rect 14967 29600 15016 29628
rect 14967 29597 14979 29600
rect 14921 29591 14979 29597
rect 10686 29560 10692 29572
rect 10192 29532 10548 29560
rect 10647 29532 10692 29560
rect 10192 29520 10198 29532
rect 10686 29520 10692 29532
rect 10744 29520 10750 29572
rect 13004 29560 13032 29591
rect 15010 29588 15016 29600
rect 15068 29588 15074 29640
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19300 29600 19625 29628
rect 19300 29588 19306 29600
rect 19613 29597 19625 29600
rect 19659 29628 19671 29631
rect 19720 29628 19748 29736
rect 20441 29699 20499 29705
rect 20441 29665 20453 29699
rect 20487 29696 20499 29699
rect 20530 29696 20536 29708
rect 20487 29668 20536 29696
rect 20487 29665 20499 29668
rect 20441 29659 20499 29665
rect 20530 29656 20536 29668
rect 20588 29656 20594 29708
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 21545 29699 21603 29705
rect 21545 29696 21557 29699
rect 20864 29668 21557 29696
rect 20864 29656 20870 29668
rect 21545 29665 21557 29668
rect 21591 29665 21603 29699
rect 22066 29696 22094 29736
rect 23198 29724 23204 29776
rect 23256 29764 23262 29776
rect 27341 29767 27399 29773
rect 27341 29764 27353 29767
rect 23256 29736 27353 29764
rect 23256 29724 23262 29736
rect 27341 29733 27353 29736
rect 27387 29733 27399 29767
rect 27341 29727 27399 29733
rect 27154 29696 27160 29708
rect 22066 29668 27160 29696
rect 21545 29659 21603 29665
rect 27154 29656 27160 29668
rect 27212 29656 27218 29708
rect 27709 29699 27767 29705
rect 27709 29696 27721 29699
rect 27264 29668 27721 29696
rect 19659 29600 19748 29628
rect 20165 29631 20223 29637
rect 19659 29597 19671 29600
rect 19613 29591 19671 29597
rect 20165 29597 20177 29631
rect 20211 29628 20223 29631
rect 20346 29628 20352 29640
rect 20211 29600 20352 29628
rect 20211 29597 20223 29600
rect 20165 29591 20223 29597
rect 20346 29588 20352 29600
rect 20404 29588 20410 29640
rect 20714 29588 20720 29640
rect 20772 29628 20778 29640
rect 20993 29631 21051 29637
rect 20993 29628 21005 29631
rect 20772 29600 21005 29628
rect 20772 29588 20778 29600
rect 20993 29597 21005 29600
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29597 21419 29631
rect 24762 29628 24768 29640
rect 24723 29600 24768 29628
rect 21361 29591 21419 29597
rect 14274 29560 14280 29572
rect 13004 29532 14280 29560
rect 14274 29520 14280 29532
rect 14332 29520 14338 29572
rect 15102 29560 15108 29572
rect 15063 29532 15108 29560
rect 15102 29520 15108 29532
rect 15160 29520 15166 29572
rect 20898 29520 20904 29572
rect 20956 29560 20962 29572
rect 21376 29560 21404 29591
rect 24762 29588 24768 29600
rect 24820 29588 24826 29640
rect 24857 29631 24915 29637
rect 24857 29597 24869 29631
rect 24903 29597 24915 29631
rect 24857 29591 24915 29597
rect 21634 29560 21640 29572
rect 20956 29532 21640 29560
rect 20956 29520 20962 29532
rect 21634 29520 21640 29532
rect 21692 29520 21698 29572
rect 24578 29520 24584 29572
rect 24636 29560 24642 29572
rect 24872 29560 24900 29591
rect 26970 29588 26976 29640
rect 27028 29628 27034 29640
rect 27264 29628 27292 29668
rect 27709 29665 27721 29668
rect 27755 29665 27767 29699
rect 27709 29659 27767 29665
rect 27816 29668 28488 29696
rect 27522 29628 27528 29640
rect 27028 29600 27292 29628
rect 27483 29600 27528 29628
rect 27028 29588 27034 29600
rect 27522 29588 27528 29600
rect 27580 29588 27586 29640
rect 27614 29588 27620 29640
rect 27672 29628 27678 29640
rect 27816 29637 27844 29668
rect 27801 29631 27859 29637
rect 27672 29600 27717 29628
rect 27672 29588 27678 29600
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 28350 29630 28356 29640
rect 28276 29628 28356 29630
rect 28263 29600 28356 29628
rect 27801 29591 27859 29597
rect 24636 29532 24900 29560
rect 24636 29520 24642 29532
rect 27706 29520 27712 29572
rect 27764 29560 27770 29572
rect 28276 29560 28304 29600
rect 28350 29588 28356 29600
rect 28408 29588 28414 29640
rect 27764 29532 28304 29560
rect 28460 29560 28488 29668
rect 28552 29637 28580 29804
rect 28902 29764 28908 29776
rect 28736 29736 28908 29764
rect 28537 29631 28595 29637
rect 28537 29597 28549 29631
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 28736 29560 28764 29736
rect 28902 29724 28908 29736
rect 28960 29764 28966 29776
rect 30009 29767 30067 29773
rect 30009 29764 30021 29767
rect 28960 29736 30021 29764
rect 28960 29724 28966 29736
rect 30009 29733 30021 29736
rect 30055 29733 30067 29767
rect 30009 29727 30067 29733
rect 28813 29699 28871 29705
rect 28813 29665 28825 29699
rect 28859 29696 28871 29699
rect 28994 29696 29000 29708
rect 28859 29668 29000 29696
rect 28859 29665 28871 29668
rect 28813 29659 28871 29665
rect 28994 29656 29000 29668
rect 29052 29696 29058 29708
rect 29052 29668 29960 29696
rect 29052 29656 29058 29668
rect 28902 29628 28908 29640
rect 28863 29600 28908 29628
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 29178 29588 29184 29640
rect 29236 29628 29242 29640
rect 29932 29637 29960 29668
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 29236 29600 29745 29628
rect 29236 29588 29242 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29917 29631 29975 29637
rect 29917 29597 29929 29631
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 28460 29532 28764 29560
rect 27764 29520 27770 29532
rect 9306 29452 9312 29504
rect 9364 29492 9370 29504
rect 9493 29495 9551 29501
rect 9493 29492 9505 29495
rect 9364 29464 9505 29492
rect 9364 29452 9370 29464
rect 9493 29461 9505 29464
rect 9539 29461 9551 29495
rect 9493 29455 9551 29461
rect 9861 29495 9919 29501
rect 9861 29461 9873 29495
rect 9907 29492 9919 29495
rect 9950 29492 9956 29504
rect 9907 29464 9956 29492
rect 9907 29461 9919 29464
rect 9861 29455 9919 29461
rect 9950 29452 9956 29464
rect 10008 29492 10014 29504
rect 10410 29492 10416 29504
rect 10008 29464 10416 29492
rect 10008 29452 10014 29464
rect 10410 29452 10416 29464
rect 10468 29492 10474 29504
rect 12618 29492 12624 29504
rect 10468 29464 12624 29492
rect 10468 29452 10474 29464
rect 12618 29452 12624 29464
rect 12676 29452 12682 29504
rect 12802 29492 12808 29504
rect 12763 29464 12808 29492
rect 12802 29452 12808 29464
rect 12860 29452 12866 29504
rect 19518 29492 19524 29504
rect 19479 29464 19524 29492
rect 19518 29452 19524 29464
rect 19576 29452 19582 29504
rect 21361 29495 21419 29501
rect 21361 29461 21373 29495
rect 21407 29492 21419 29495
rect 21450 29492 21456 29504
rect 21407 29464 21456 29492
rect 21407 29461 21419 29464
rect 21361 29455 21419 29461
rect 21450 29452 21456 29464
rect 21508 29452 21514 29504
rect 1104 29402 35027 29424
rect 1104 29350 9390 29402
rect 9442 29350 9454 29402
rect 9506 29350 9518 29402
rect 9570 29350 9582 29402
rect 9634 29350 9646 29402
rect 9698 29350 17831 29402
rect 17883 29350 17895 29402
rect 17947 29350 17959 29402
rect 18011 29350 18023 29402
rect 18075 29350 18087 29402
rect 18139 29350 26272 29402
rect 26324 29350 26336 29402
rect 26388 29350 26400 29402
rect 26452 29350 26464 29402
rect 26516 29350 26528 29402
rect 26580 29350 34713 29402
rect 34765 29350 34777 29402
rect 34829 29350 34841 29402
rect 34893 29350 34905 29402
rect 34957 29350 34969 29402
rect 35021 29350 35027 29402
rect 1104 29328 35027 29350
rect 12894 29248 12900 29300
rect 12952 29248 12958 29300
rect 14550 29288 14556 29300
rect 14511 29260 14556 29288
rect 14550 29248 14556 29260
rect 14608 29248 14614 29300
rect 14918 29248 14924 29300
rect 14976 29288 14982 29300
rect 20162 29288 20168 29300
rect 14976 29260 17724 29288
rect 20123 29260 20168 29288
rect 14976 29248 14982 29260
rect 12912 29220 12940 29248
rect 12544 29192 12940 29220
rect 9030 29152 9036 29164
rect 8991 29124 9036 29152
rect 9030 29112 9036 29124
rect 9088 29112 9094 29164
rect 9306 29152 9312 29164
rect 9267 29124 9312 29152
rect 9306 29112 9312 29124
rect 9364 29112 9370 29164
rect 9490 29152 9496 29164
rect 9451 29124 9496 29152
rect 9490 29112 9496 29124
rect 9548 29112 9554 29164
rect 11790 29152 11796 29164
rect 11751 29124 11796 29152
rect 11790 29112 11796 29124
rect 11848 29112 11854 29164
rect 12544 29161 12572 29192
rect 15102 29180 15108 29232
rect 15160 29220 15166 29232
rect 17696 29229 17724 29260
rect 20162 29248 20168 29260
rect 20220 29248 20226 29300
rect 21358 29248 21364 29300
rect 21416 29288 21422 29300
rect 22097 29291 22155 29297
rect 22097 29288 22109 29291
rect 21416 29260 22109 29288
rect 21416 29248 21422 29260
rect 22097 29257 22109 29260
rect 22143 29257 22155 29291
rect 22097 29251 22155 29257
rect 27614 29248 27620 29300
rect 27672 29288 27678 29300
rect 27893 29291 27951 29297
rect 27893 29288 27905 29291
rect 27672 29260 27905 29288
rect 27672 29248 27678 29260
rect 27893 29257 27905 29260
rect 27939 29257 27951 29291
rect 27893 29251 27951 29257
rect 28350 29248 28356 29300
rect 28408 29288 28414 29300
rect 28921 29291 28979 29297
rect 28921 29288 28933 29291
rect 28408 29260 28933 29288
rect 28408 29248 28414 29260
rect 28921 29257 28933 29260
rect 28967 29257 28979 29291
rect 28921 29251 28979 29257
rect 29089 29291 29147 29297
rect 29089 29257 29101 29291
rect 29135 29288 29147 29291
rect 29178 29288 29184 29300
rect 29135 29260 29184 29288
rect 29135 29257 29147 29260
rect 29089 29251 29147 29257
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 15381 29223 15439 29229
rect 15381 29220 15393 29223
rect 15160 29192 15393 29220
rect 15160 29180 15166 29192
rect 15381 29189 15393 29192
rect 15427 29189 15439 29223
rect 15381 29183 15439 29189
rect 17681 29223 17739 29229
rect 17681 29189 17693 29223
rect 17727 29189 17739 29223
rect 20530 29220 20536 29232
rect 17681 29183 17739 29189
rect 20364 29192 20536 29220
rect 12529 29155 12587 29161
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 12618 29112 12624 29164
rect 12676 29152 12682 29164
rect 12676 29124 12721 29152
rect 12676 29112 12682 29124
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 12897 29155 12955 29161
rect 12897 29152 12909 29155
rect 12860 29124 12909 29152
rect 12860 29112 12866 29124
rect 12897 29121 12909 29124
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 13173 29155 13231 29161
rect 13173 29121 13185 29155
rect 13219 29152 13231 29155
rect 13446 29152 13452 29164
rect 13219 29124 13452 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 13446 29112 13452 29124
rect 13504 29112 13510 29164
rect 14737 29155 14795 29161
rect 14737 29121 14749 29155
rect 14783 29152 14795 29155
rect 15120 29152 15148 29180
rect 15562 29152 15568 29164
rect 14783 29124 15148 29152
rect 15523 29124 15568 29152
rect 14783 29121 14795 29124
rect 14737 29115 14795 29121
rect 15562 29112 15568 29124
rect 15620 29112 15626 29164
rect 15746 29152 15752 29164
rect 15707 29124 15752 29152
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 19153 29155 19211 29161
rect 19153 29121 19165 29155
rect 19199 29152 19211 29155
rect 19334 29152 19340 29164
rect 19199 29124 19340 29152
rect 19199 29121 19211 29124
rect 19153 29115 19211 29121
rect 19334 29112 19340 29124
rect 19392 29112 19398 29164
rect 19518 29152 19524 29164
rect 19479 29124 19524 29152
rect 19518 29112 19524 29124
rect 19576 29112 19582 29164
rect 20364 29161 20392 29192
rect 20530 29180 20536 29192
rect 20588 29220 20594 29232
rect 20588 29192 21404 29220
rect 20588 29180 20594 29192
rect 20349 29155 20407 29161
rect 20349 29121 20361 29155
rect 20395 29121 20407 29155
rect 20349 29115 20407 29121
rect 20438 29112 20444 29164
rect 20496 29152 20502 29164
rect 20622 29152 20628 29164
rect 20496 29124 20541 29152
rect 20583 29124 20628 29152
rect 20496 29112 20502 29124
rect 20622 29112 20628 29124
rect 20680 29112 20686 29164
rect 20714 29112 20720 29164
rect 20772 29152 20778 29164
rect 21376 29161 21404 29192
rect 21634 29180 21640 29232
rect 21692 29220 21698 29232
rect 25222 29220 25228 29232
rect 21692 29192 22600 29220
rect 25183 29192 25228 29220
rect 21692 29180 21698 29192
rect 21177 29155 21235 29161
rect 21177 29152 21189 29155
rect 20772 29124 20817 29152
rect 20916 29124 21189 29152
rect 20772 29112 20778 29124
rect 14921 29087 14979 29093
rect 14921 29053 14933 29087
rect 14967 29084 14979 29087
rect 15010 29084 15016 29096
rect 14967 29056 15016 29084
rect 14967 29053 14979 29056
rect 14921 29047 14979 29053
rect 15010 29044 15016 29056
rect 15068 29044 15074 29096
rect 20456 29016 20484 29112
rect 20916 29016 20944 29124
rect 21177 29121 21189 29124
rect 21223 29121 21235 29155
rect 21177 29115 21235 29121
rect 21361 29155 21419 29161
rect 21361 29121 21373 29155
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29152 22339 29155
rect 22370 29152 22376 29164
rect 22327 29124 22376 29152
rect 22327 29121 22339 29124
rect 22281 29115 22339 29121
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 22572 29161 22600 29192
rect 25222 29180 25228 29192
rect 25280 29180 25286 29232
rect 27249 29223 27307 29229
rect 27249 29189 27261 29223
rect 27295 29220 27307 29223
rect 28721 29223 28779 29229
rect 27295 29192 28120 29220
rect 27295 29189 27307 29192
rect 27249 29183 27307 29189
rect 28092 29164 28120 29192
rect 28721 29189 28733 29223
rect 28767 29189 28779 29223
rect 28721 29183 28779 29189
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22738 29152 22744 29164
rect 22699 29124 22744 29152
rect 22557 29115 22615 29121
rect 22738 29112 22744 29124
rect 22796 29112 22802 29164
rect 22830 29112 22836 29164
rect 22888 29152 22894 29164
rect 23382 29152 23388 29164
rect 22888 29124 23388 29152
rect 22888 29112 22894 29124
rect 23382 29112 23388 29124
rect 23440 29152 23446 29164
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 23440 29124 25329 29152
rect 23440 29112 23446 29124
rect 25317 29121 25329 29124
rect 25363 29121 25375 29155
rect 25317 29115 25375 29121
rect 25593 29155 25651 29161
rect 25593 29121 25605 29155
rect 25639 29152 25651 29155
rect 25774 29152 25780 29164
rect 25639 29124 25780 29152
rect 25639 29121 25651 29124
rect 25593 29115 25651 29121
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 27154 29152 27160 29164
rect 27115 29124 27160 29152
rect 27154 29112 27160 29124
rect 27212 29112 27218 29164
rect 27338 29152 27344 29164
rect 27299 29124 27344 29152
rect 27338 29112 27344 29124
rect 27396 29112 27402 29164
rect 28074 29152 28080 29164
rect 28035 29124 28080 29152
rect 28074 29112 28080 29124
rect 28132 29112 28138 29164
rect 27172 29084 27200 29112
rect 28166 29084 28172 29096
rect 27172 29056 28172 29084
rect 28166 29044 28172 29056
rect 28224 29044 28230 29096
rect 28261 29087 28319 29093
rect 28261 29053 28273 29087
rect 28307 29084 28319 29087
rect 28626 29084 28632 29096
rect 28307 29056 28632 29084
rect 28307 29053 28319 29056
rect 28261 29047 28319 29053
rect 28626 29044 28632 29056
rect 28684 29044 28690 29096
rect 21266 29016 21272 29028
rect 20456 28988 20944 29016
rect 21227 28988 21272 29016
rect 21266 28976 21272 28988
rect 21324 28976 21330 29028
rect 22373 29019 22431 29025
rect 22373 29016 22385 29019
rect 22066 28988 22385 29016
rect 8938 28908 8944 28960
rect 8996 28948 9002 28960
rect 9401 28951 9459 28957
rect 9401 28948 9413 28951
rect 8996 28920 9413 28948
rect 8996 28908 9002 28920
rect 9401 28917 9413 28920
rect 9447 28917 9459 28951
rect 9401 28911 9459 28917
rect 10594 28908 10600 28960
rect 10652 28948 10658 28960
rect 11793 28951 11851 28957
rect 11793 28948 11805 28951
rect 10652 28920 11805 28948
rect 10652 28908 10658 28920
rect 11793 28917 11805 28920
rect 11839 28917 11851 28951
rect 11793 28911 11851 28917
rect 20714 28908 20720 28960
rect 20772 28948 20778 28960
rect 22066 28948 22094 28988
rect 22373 28985 22385 28988
rect 22419 28985 22431 29019
rect 22373 28979 22431 28985
rect 22462 28976 22468 29028
rect 22520 29016 22526 29028
rect 22520 28988 22565 29016
rect 22520 28976 22526 28988
rect 27522 28976 27528 29028
rect 27580 29016 27586 29028
rect 28736 29016 28764 29183
rect 27580 28988 28764 29016
rect 27580 28976 27586 28988
rect 28902 28948 28908 28960
rect 20772 28920 22094 28948
rect 28863 28920 28908 28948
rect 20772 28908 20778 28920
rect 28902 28908 28908 28920
rect 28960 28908 28966 28960
rect 1104 28858 34868 28880
rect 1104 28806 5170 28858
rect 5222 28806 5234 28858
rect 5286 28806 5298 28858
rect 5350 28806 5362 28858
rect 5414 28806 5426 28858
rect 5478 28806 13611 28858
rect 13663 28806 13675 28858
rect 13727 28806 13739 28858
rect 13791 28806 13803 28858
rect 13855 28806 13867 28858
rect 13919 28806 22052 28858
rect 22104 28806 22116 28858
rect 22168 28806 22180 28858
rect 22232 28806 22244 28858
rect 22296 28806 22308 28858
rect 22360 28806 30493 28858
rect 30545 28806 30557 28858
rect 30609 28806 30621 28858
rect 30673 28806 30685 28858
rect 30737 28806 30749 28858
rect 30801 28806 34868 28858
rect 1104 28784 34868 28806
rect 21174 28744 21180 28756
rect 21135 28716 21180 28744
rect 21174 28704 21180 28716
rect 21232 28704 21238 28756
rect 28813 28747 28871 28753
rect 28813 28713 28825 28747
rect 28859 28744 28871 28747
rect 28902 28744 28908 28756
rect 28859 28716 28908 28744
rect 28859 28713 28871 28716
rect 28813 28707 28871 28713
rect 28902 28704 28908 28716
rect 28960 28704 28966 28756
rect 13446 28636 13452 28688
rect 13504 28676 13510 28688
rect 15197 28679 15255 28685
rect 15197 28676 15209 28679
rect 13504 28648 15209 28676
rect 13504 28636 13510 28648
rect 15197 28645 15209 28648
rect 15243 28645 15255 28679
rect 20714 28676 20720 28688
rect 15197 28639 15255 28645
rect 20180 28648 20720 28676
rect 9490 28608 9496 28620
rect 9324 28580 9496 28608
rect 9324 28549 9352 28580
rect 9490 28568 9496 28580
rect 9548 28608 9554 28620
rect 10965 28611 11023 28617
rect 10965 28608 10977 28611
rect 9548 28580 10977 28608
rect 9548 28568 9554 28580
rect 10965 28577 10977 28580
rect 11011 28577 11023 28611
rect 10965 28571 11023 28577
rect 11609 28611 11667 28617
rect 11609 28577 11621 28611
rect 11655 28608 11667 28611
rect 11790 28608 11796 28620
rect 11655 28580 11796 28608
rect 11655 28577 11667 28580
rect 11609 28571 11667 28577
rect 11790 28568 11796 28580
rect 11848 28608 11854 28620
rect 12526 28608 12532 28620
rect 11848 28580 12532 28608
rect 11848 28568 11854 28580
rect 12526 28568 12532 28580
rect 12584 28608 12590 28620
rect 13173 28611 13231 28617
rect 13173 28608 13185 28611
rect 12584 28580 13185 28608
rect 12584 28568 12590 28580
rect 13173 28577 13185 28580
rect 13219 28577 13231 28611
rect 13173 28571 13231 28577
rect 13358 28611 13416 28617
rect 13358 28577 13370 28611
rect 13404 28608 13416 28611
rect 13464 28608 13492 28636
rect 13404 28580 13492 28608
rect 13404 28577 13416 28580
rect 13358 28571 13416 28577
rect 15010 28568 15016 28620
rect 15068 28608 15074 28620
rect 20180 28617 20208 28648
rect 20714 28636 20720 28648
rect 20772 28636 20778 28688
rect 20165 28611 20223 28617
rect 15068 28580 19840 28608
rect 15068 28568 15074 28580
rect 19812 28552 19840 28580
rect 20165 28577 20177 28611
rect 20211 28577 20223 28611
rect 20165 28571 20223 28577
rect 20806 28568 20812 28620
rect 20864 28608 20870 28620
rect 26237 28611 26295 28617
rect 20864 28580 21036 28608
rect 20864 28568 20870 28580
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28509 9367 28543
rect 9309 28503 9367 28509
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28509 9643 28543
rect 9585 28503 9643 28509
rect 9030 28432 9036 28484
rect 9088 28472 9094 28484
rect 9600 28472 9628 28503
rect 10686 28500 10692 28552
rect 10744 28540 10750 28552
rect 11330 28540 11336 28552
rect 10744 28512 11336 28540
rect 10744 28500 10750 28512
rect 11330 28500 11336 28512
rect 11388 28500 11394 28552
rect 12069 28543 12127 28549
rect 12069 28509 12081 28543
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28540 12403 28543
rect 12802 28540 12808 28552
rect 12391 28512 12808 28540
rect 12391 28509 12403 28512
rect 12345 28503 12403 28509
rect 9088 28444 9628 28472
rect 12084 28472 12112 28503
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 13078 28540 13084 28552
rect 13039 28512 13084 28540
rect 13078 28500 13084 28512
rect 13136 28500 13142 28552
rect 13262 28500 13268 28552
rect 13320 28540 13326 28552
rect 14550 28540 14556 28552
rect 13320 28512 13365 28540
rect 14511 28512 14556 28540
rect 13320 28500 13326 28512
rect 14550 28500 14556 28512
rect 14608 28500 14614 28552
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28540 14979 28543
rect 15102 28540 15108 28552
rect 14967 28512 15108 28540
rect 14967 28509 14979 28512
rect 14921 28503 14979 28509
rect 15102 28500 15108 28512
rect 15160 28500 15166 28552
rect 15378 28540 15384 28552
rect 15339 28512 15384 28540
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 15470 28500 15476 28552
rect 15528 28540 15534 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 15528 28512 16313 28540
rect 15528 28500 15534 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 19794 28540 19800 28552
rect 19755 28512 19800 28540
rect 16301 28503 16359 28509
rect 19794 28500 19800 28512
rect 19852 28500 19858 28552
rect 19978 28540 19984 28552
rect 19939 28512 19984 28540
rect 19978 28500 19984 28512
rect 20036 28500 20042 28552
rect 20714 28549 20720 28552
rect 20615 28543 20673 28549
rect 20615 28540 20627 28543
rect 20548 28512 20627 28540
rect 13446 28472 13452 28484
rect 12084 28444 13452 28472
rect 9088 28432 9094 28444
rect 13446 28432 13452 28444
rect 13504 28432 13510 28484
rect 15746 28432 15752 28484
rect 15804 28472 15810 28484
rect 16669 28475 16727 28481
rect 16669 28472 16681 28475
rect 15804 28444 16681 28472
rect 15804 28432 15810 28444
rect 16669 28441 16681 28444
rect 16715 28472 16727 28475
rect 19242 28472 19248 28484
rect 16715 28444 19248 28472
rect 16715 28441 16727 28444
rect 16669 28435 16727 28441
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 20548 28416 20576 28512
rect 20615 28509 20627 28512
rect 20661 28509 20673 28543
rect 20615 28503 20673 28509
rect 20705 28543 20720 28549
rect 20705 28509 20717 28543
rect 20705 28503 20720 28509
rect 20714 28500 20720 28503
rect 20772 28500 20778 28552
rect 20898 28540 20904 28552
rect 20859 28512 20904 28540
rect 20898 28500 20904 28512
rect 20956 28500 20962 28552
rect 21008 28549 21036 28580
rect 26237 28577 26249 28611
rect 26283 28608 26295 28611
rect 26694 28608 26700 28620
rect 26283 28580 26700 28608
rect 26283 28577 26295 28580
rect 26237 28571 26295 28577
rect 26694 28568 26700 28580
rect 26752 28568 26758 28620
rect 27614 28568 27620 28620
rect 27672 28568 27678 28620
rect 20993 28543 21051 28549
rect 20993 28509 21005 28543
rect 21039 28540 21051 28543
rect 22830 28540 22836 28552
rect 21039 28512 22094 28540
rect 22791 28512 22836 28540
rect 21039 28509 21051 28512
rect 20993 28503 21051 28509
rect 22066 28472 22094 28512
rect 22830 28500 22836 28512
rect 22888 28500 22894 28552
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28540 23443 28543
rect 23566 28540 23572 28552
rect 23431 28512 23572 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 23566 28500 23572 28512
rect 23624 28540 23630 28552
rect 24670 28540 24676 28552
rect 23624 28512 24676 28540
rect 23624 28500 23630 28512
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 27890 28540 27896 28552
rect 27738 28512 27896 28540
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28718 28540 28724 28552
rect 28679 28512 28724 28540
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 22066 28444 22494 28472
rect 9122 28404 9128 28416
rect 9083 28376 9128 28404
rect 9122 28364 9128 28376
rect 9180 28364 9186 28416
rect 9306 28364 9312 28416
rect 9364 28404 9370 28416
rect 9493 28407 9551 28413
rect 9493 28404 9505 28407
rect 9364 28376 9505 28404
rect 9364 28364 9370 28376
rect 9493 28373 9505 28376
rect 9539 28373 9551 28407
rect 12894 28404 12900 28416
rect 12855 28376 12900 28404
rect 9493 28367 9551 28373
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 13078 28364 13084 28416
rect 13136 28404 13142 28416
rect 15930 28404 15936 28416
rect 13136 28376 15936 28404
rect 13136 28364 13142 28376
rect 15930 28364 15936 28376
rect 15988 28364 15994 28416
rect 20530 28404 20536 28416
rect 20443 28376 20536 28404
rect 20530 28364 20536 28376
rect 20588 28404 20594 28416
rect 22738 28404 22744 28416
rect 20588 28376 22744 28404
rect 20588 28364 20594 28376
rect 22738 28364 22744 28376
rect 22796 28364 22802 28416
rect 27246 28404 27252 28416
rect 27207 28376 27252 28404
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 1104 28314 35027 28336
rect 1104 28262 9390 28314
rect 9442 28262 9454 28314
rect 9506 28262 9518 28314
rect 9570 28262 9582 28314
rect 9634 28262 9646 28314
rect 9698 28262 17831 28314
rect 17883 28262 17895 28314
rect 17947 28262 17959 28314
rect 18011 28262 18023 28314
rect 18075 28262 18087 28314
rect 18139 28262 26272 28314
rect 26324 28262 26336 28314
rect 26388 28262 26400 28314
rect 26452 28262 26464 28314
rect 26516 28262 26528 28314
rect 26580 28262 34713 28314
rect 34765 28262 34777 28314
rect 34829 28262 34841 28314
rect 34893 28262 34905 28314
rect 34957 28262 34969 28314
rect 35021 28262 35027 28314
rect 1104 28240 35027 28262
rect 8113 28203 8171 28209
rect 8113 28169 8125 28203
rect 8159 28200 8171 28203
rect 8938 28200 8944 28212
rect 8159 28172 8944 28200
rect 8159 28169 8171 28172
rect 8113 28163 8171 28169
rect 8938 28160 8944 28172
rect 8996 28160 9002 28212
rect 11330 28160 11336 28212
rect 11388 28200 11394 28212
rect 13078 28200 13084 28212
rect 11388 28172 13084 28200
rect 11388 28160 11394 28172
rect 9140 28104 9904 28132
rect 9140 28076 9168 28104
rect 7929 28067 7987 28073
rect 7929 28033 7941 28067
rect 7975 28033 7987 28067
rect 7929 28027 7987 28033
rect 8205 28067 8263 28073
rect 8205 28033 8217 28067
rect 8251 28064 8263 28067
rect 9033 28067 9091 28073
rect 9033 28064 9045 28067
rect 8251 28036 9045 28064
rect 8251 28033 8263 28036
rect 8205 28027 8263 28033
rect 9033 28033 9045 28036
rect 9079 28064 9091 28067
rect 9122 28064 9128 28076
rect 9079 28036 9128 28064
rect 9079 28033 9091 28036
rect 9033 28027 9091 28033
rect 7944 27928 7972 28027
rect 9122 28024 9128 28036
rect 9180 28024 9186 28076
rect 9876 28073 9904 28104
rect 9677 28067 9735 28073
rect 9677 28033 9689 28067
rect 9723 28033 9735 28067
rect 9677 28027 9735 28033
rect 9861 28067 9919 28073
rect 9861 28033 9873 28067
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 12161 28067 12219 28073
rect 12161 28033 12173 28067
rect 12207 28064 12219 28067
rect 12406 28064 12434 28172
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 15378 28200 15384 28212
rect 15339 28172 15384 28200
rect 15378 28160 15384 28172
rect 15436 28160 15442 28212
rect 19794 28160 19800 28212
rect 19852 28200 19858 28212
rect 22281 28203 22339 28209
rect 19852 28172 22094 28200
rect 19852 28160 19858 28172
rect 13446 28132 13452 28144
rect 12912 28104 13452 28132
rect 12526 28064 12532 28076
rect 12207 28036 12434 28064
rect 12487 28036 12532 28064
rect 12207 28033 12219 28036
rect 12161 28027 12219 28033
rect 8754 27996 8760 28008
rect 8715 27968 8760 27996
rect 8754 27956 8760 27968
rect 8812 27956 8818 28008
rect 8849 27999 8907 28005
rect 8849 27965 8861 27999
rect 8895 27965 8907 27999
rect 8849 27959 8907 27965
rect 8864 27928 8892 27959
rect 8938 27956 8944 28008
rect 8996 27996 9002 28008
rect 9692 27996 9720 28027
rect 12526 28024 12532 28036
rect 12584 28024 12590 28076
rect 12912 28073 12940 28104
rect 13446 28092 13452 28104
rect 13504 28092 13510 28144
rect 15010 28132 15016 28144
rect 14016 28104 15016 28132
rect 14016 28076 14044 28104
rect 15010 28092 15016 28104
rect 15068 28092 15074 28144
rect 15562 28092 15568 28144
rect 15620 28132 15626 28144
rect 15933 28135 15991 28141
rect 15933 28132 15945 28135
rect 15620 28104 15945 28132
rect 15620 28092 15626 28104
rect 15933 28101 15945 28104
rect 15979 28132 15991 28135
rect 16022 28132 16028 28144
rect 15979 28104 16028 28132
rect 15979 28101 15991 28104
rect 15933 28095 15991 28101
rect 16022 28092 16028 28104
rect 16080 28092 16086 28144
rect 19334 28092 19340 28144
rect 19392 28132 19398 28144
rect 20625 28135 20683 28141
rect 19392 28104 19472 28132
rect 19392 28092 19398 28104
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 13262 28024 13268 28076
rect 13320 28064 13326 28076
rect 13357 28067 13415 28073
rect 13357 28064 13369 28067
rect 13320 28036 13369 28064
rect 13320 28024 13326 28036
rect 13357 28033 13369 28036
rect 13403 28064 13415 28067
rect 13817 28067 13875 28073
rect 13817 28064 13829 28067
rect 13403 28036 13829 28064
rect 13403 28033 13415 28036
rect 13357 28027 13415 28033
rect 13817 28033 13829 28036
rect 13863 28033 13875 28067
rect 13817 28027 13875 28033
rect 13998 28024 14004 28076
rect 14056 28064 14062 28076
rect 14185 28067 14243 28073
rect 14056 28036 14149 28064
rect 14056 28024 14062 28036
rect 14185 28033 14197 28067
rect 14231 28064 14243 28067
rect 14274 28064 14280 28076
rect 14231 28036 14280 28064
rect 14231 28033 14243 28036
rect 14185 28027 14243 28033
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28064 15439 28067
rect 15470 28064 15476 28076
rect 15427 28036 15476 28064
rect 15427 28033 15439 28036
rect 15381 28027 15439 28033
rect 15470 28024 15476 28036
rect 15528 28024 15534 28076
rect 19242 28064 19248 28076
rect 19203 28036 19248 28064
rect 19242 28024 19248 28036
rect 19300 28024 19306 28076
rect 19444 28073 19472 28104
rect 20625 28101 20637 28135
rect 20671 28132 20683 28135
rect 20898 28132 20904 28144
rect 20671 28104 20904 28132
rect 20671 28101 20683 28104
rect 20625 28095 20683 28101
rect 20898 28092 20904 28104
rect 20956 28092 20962 28144
rect 22066 28132 22094 28172
rect 22281 28169 22293 28203
rect 22327 28200 22339 28203
rect 22370 28200 22376 28212
rect 22327 28172 22376 28200
rect 22327 28169 22339 28172
rect 22281 28163 22339 28169
rect 22370 28160 22376 28172
rect 22428 28160 22434 28212
rect 22462 28160 22468 28212
rect 22520 28200 22526 28212
rect 23201 28203 23259 28209
rect 23201 28200 23213 28203
rect 22520 28172 23213 28200
rect 22520 28160 22526 28172
rect 23201 28169 23213 28172
rect 23247 28169 23259 28203
rect 23201 28163 23259 28169
rect 23566 28132 23572 28144
rect 22066 28104 22416 28132
rect 19429 28067 19487 28073
rect 19429 28033 19441 28067
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 20257 28067 20315 28073
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20257 28027 20315 28033
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28064 20591 28067
rect 22278 28064 22284 28076
rect 20579 28036 22284 28064
rect 20579 28033 20591 28036
rect 20533 28027 20591 28033
rect 8996 27968 9720 27996
rect 8996 27956 9002 27968
rect 9766 27956 9772 28008
rect 9824 27956 9830 28008
rect 12434 27956 12440 28008
rect 12492 27996 12498 28008
rect 12492 27968 12537 27996
rect 12492 27956 12498 27968
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 14608 27968 15301 27996
rect 14608 27956 14614 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15289 27959 15347 27965
rect 19337 27999 19395 28005
rect 19337 27965 19349 27999
rect 19383 27996 19395 27999
rect 19978 27996 19984 28008
rect 19383 27968 19984 27996
rect 19383 27965 19395 27968
rect 19337 27959 19395 27965
rect 19978 27956 19984 27968
rect 20036 27996 20042 28008
rect 20272 27996 20300 28027
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 20036 27968 20300 27996
rect 20036 27956 20042 27968
rect 9784 27928 9812 27956
rect 7944 27900 9812 27928
rect 7745 27863 7803 27869
rect 7745 27829 7757 27863
rect 7791 27860 7803 27863
rect 9122 27860 9128 27872
rect 7791 27832 9128 27860
rect 7791 27829 7803 27832
rect 7745 27823 7803 27829
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9217 27863 9275 27869
rect 9217 27829 9229 27863
rect 9263 27860 9275 27863
rect 9306 27860 9312 27872
rect 9263 27832 9312 27860
rect 9263 27829 9275 27832
rect 9217 27823 9275 27829
rect 9306 27820 9312 27832
rect 9364 27860 9370 27872
rect 9582 27860 9588 27872
rect 9364 27832 9588 27860
rect 9364 27820 9370 27832
rect 9582 27820 9588 27832
rect 9640 27820 9646 27872
rect 9766 27860 9772 27872
rect 9727 27832 9772 27860
rect 9766 27820 9772 27832
rect 9824 27820 9830 27872
rect 22388 27860 22416 28104
rect 22480 28104 23572 28132
rect 22480 27937 22508 28104
rect 23566 28092 23572 28104
rect 23624 28132 23630 28144
rect 23661 28135 23719 28141
rect 23661 28132 23673 28135
rect 23624 28104 23673 28132
rect 23624 28092 23630 28104
rect 23661 28101 23673 28104
rect 23707 28101 23719 28135
rect 27338 28132 27344 28144
rect 23661 28095 23719 28101
rect 24044 28104 27344 28132
rect 22741 27999 22799 28005
rect 22741 27965 22753 27999
rect 22787 27996 22799 27999
rect 22830 27996 22836 28008
rect 22787 27968 22836 27996
rect 22787 27965 22799 27968
rect 22741 27959 22799 27965
rect 22465 27931 22523 27937
rect 22465 27897 22477 27931
rect 22511 27897 22523 27931
rect 22756 27928 22784 27959
rect 22830 27956 22836 27968
rect 22888 27956 22894 28008
rect 23385 27931 23443 27937
rect 23385 27928 23397 27931
rect 22756 27900 23397 27928
rect 22465 27891 22523 27897
rect 23385 27897 23397 27900
rect 23431 27928 23443 27931
rect 24044 27928 24072 28104
rect 27338 28092 27344 28104
rect 27396 28132 27402 28144
rect 30285 28135 30343 28141
rect 30285 28132 30297 28135
rect 27396 28104 30297 28132
rect 27396 28092 27402 28104
rect 30285 28101 30297 28104
rect 30331 28132 30343 28135
rect 31110 28132 31116 28144
rect 30331 28104 31116 28132
rect 30331 28101 30343 28104
rect 30285 28095 30343 28101
rect 31110 28092 31116 28104
rect 31168 28092 31174 28144
rect 24854 28024 24860 28076
rect 24912 28064 24918 28076
rect 25041 28067 25099 28073
rect 25041 28064 25053 28067
rect 24912 28036 25053 28064
rect 24912 28024 24918 28036
rect 25041 28033 25053 28036
rect 25087 28033 25099 28067
rect 25682 28064 25688 28076
rect 25643 28036 25688 28064
rect 25041 28027 25099 28033
rect 25682 28024 25688 28036
rect 25740 28024 25746 28076
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 27249 28067 27307 28073
rect 27249 28064 27261 28067
rect 27120 28036 27261 28064
rect 27120 28024 27126 28036
rect 27249 28033 27261 28036
rect 27295 28033 27307 28067
rect 27249 28027 27307 28033
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28064 27583 28067
rect 27706 28064 27712 28076
rect 27571 28036 27712 28064
rect 27571 28033 27583 28036
rect 27525 28027 27583 28033
rect 27706 28024 27712 28036
rect 27764 28024 27770 28076
rect 28994 28024 29000 28076
rect 29052 28064 29058 28076
rect 30101 28067 30159 28073
rect 30101 28064 30113 28067
rect 29052 28036 30113 28064
rect 29052 28024 29058 28036
rect 30101 28033 30113 28036
rect 30147 28033 30159 28067
rect 30101 28027 30159 28033
rect 30377 28067 30435 28073
rect 30377 28033 30389 28067
rect 30423 28064 30435 28067
rect 32674 28064 32680 28076
rect 30423 28036 32680 28064
rect 30423 28033 30435 28036
rect 30377 28027 30435 28033
rect 32674 28024 32680 28036
rect 32732 28024 32738 28076
rect 25130 27956 25136 28008
rect 25188 27956 25194 28008
rect 25774 27996 25780 28008
rect 25735 27968 25780 27996
rect 25774 27956 25780 27968
rect 25832 27956 25838 28008
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 27157 27999 27215 28005
rect 27157 27996 27169 27999
rect 26292 27968 27169 27996
rect 26292 27956 26298 27968
rect 27157 27965 27169 27968
rect 27203 27965 27215 27999
rect 27157 27959 27215 27965
rect 23431 27900 24072 27928
rect 24857 27931 24915 27937
rect 23431 27897 23443 27900
rect 23385 27891 23443 27897
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25866 27928 25872 27940
rect 24903 27900 25872 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25866 27888 25872 27900
rect 25924 27888 25930 27940
rect 26602 27860 26608 27872
rect 22388 27832 26608 27860
rect 26602 27820 26608 27832
rect 26660 27820 26666 27872
rect 29917 27863 29975 27869
rect 29917 27829 29929 27863
rect 29963 27860 29975 27863
rect 30006 27860 30012 27872
rect 29963 27832 30012 27860
rect 29963 27829 29975 27832
rect 29917 27823 29975 27829
rect 30006 27820 30012 27832
rect 30064 27820 30070 27872
rect 1104 27770 34868 27792
rect 1104 27718 5170 27770
rect 5222 27718 5234 27770
rect 5286 27718 5298 27770
rect 5350 27718 5362 27770
rect 5414 27718 5426 27770
rect 5478 27718 13611 27770
rect 13663 27718 13675 27770
rect 13727 27718 13739 27770
rect 13791 27718 13803 27770
rect 13855 27718 13867 27770
rect 13919 27718 22052 27770
rect 22104 27718 22116 27770
rect 22168 27718 22180 27770
rect 22232 27718 22244 27770
rect 22296 27718 22308 27770
rect 22360 27718 30493 27770
rect 30545 27718 30557 27770
rect 30609 27718 30621 27770
rect 30673 27718 30685 27770
rect 30737 27718 30749 27770
rect 30801 27718 34868 27770
rect 1104 27696 34868 27718
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 24670 27656 24676 27668
rect 22428 27628 24676 27656
rect 22428 27616 22434 27628
rect 24670 27616 24676 27628
rect 24728 27616 24734 27668
rect 16022 27548 16028 27600
rect 16080 27588 16086 27600
rect 16853 27591 16911 27597
rect 16853 27588 16865 27591
rect 16080 27560 16865 27588
rect 16080 27548 16086 27560
rect 16853 27557 16865 27560
rect 16899 27557 16911 27591
rect 16853 27551 16911 27557
rect 24578 27548 24584 27600
rect 24636 27588 24642 27600
rect 25225 27591 25283 27597
rect 25225 27588 25237 27591
rect 24636 27560 25237 27588
rect 24636 27548 24642 27560
rect 25225 27557 25237 27560
rect 25271 27557 25283 27591
rect 27890 27588 27896 27600
rect 27851 27560 27896 27588
rect 25225 27551 25283 27557
rect 27890 27548 27896 27560
rect 27948 27548 27954 27600
rect 9030 27480 9036 27532
rect 9088 27520 9094 27532
rect 9217 27523 9275 27529
rect 9217 27520 9229 27523
rect 9088 27492 9229 27520
rect 9088 27480 9094 27492
rect 9217 27489 9229 27492
rect 9263 27489 9275 27523
rect 9217 27483 9275 27489
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 12805 27523 12863 27529
rect 12805 27520 12817 27523
rect 12584 27492 12817 27520
rect 12584 27480 12590 27492
rect 12805 27489 12817 27492
rect 12851 27489 12863 27523
rect 13998 27520 14004 27532
rect 12805 27483 12863 27489
rect 13188 27492 14004 27520
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9309 27455 9367 27461
rect 9309 27452 9321 27455
rect 9180 27424 9321 27452
rect 9180 27412 9186 27424
rect 9309 27421 9321 27424
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 13188 27461 13216 27492
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 19886 27480 19892 27532
rect 19944 27520 19950 27532
rect 19944 27492 22324 27520
rect 19944 27480 19950 27492
rect 9677 27455 9735 27461
rect 9677 27452 9689 27455
rect 9640 27424 9689 27452
rect 9640 27412 9646 27424
rect 9677 27421 9689 27424
rect 9723 27421 9735 27455
rect 9677 27415 9735 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13814 27452 13820 27464
rect 13403 27424 13820 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27421 14979 27455
rect 14921 27415 14979 27421
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 8202 27344 8208 27396
rect 8260 27384 8266 27396
rect 10137 27387 10195 27393
rect 10137 27384 10149 27387
rect 8260 27356 10149 27384
rect 8260 27344 8266 27356
rect 10137 27353 10149 27356
rect 10183 27384 10195 27387
rect 12342 27384 12348 27396
rect 10183 27356 12348 27384
rect 10183 27353 10195 27356
rect 10137 27347 10195 27353
rect 12342 27344 12348 27356
rect 12400 27344 12406 27396
rect 12618 27344 12624 27396
rect 12676 27384 12682 27396
rect 13722 27384 13728 27396
rect 12676 27356 13728 27384
rect 12676 27344 12682 27356
rect 13722 27344 13728 27356
rect 13780 27384 13786 27396
rect 14369 27387 14427 27393
rect 14369 27384 14381 27387
rect 13780 27356 14381 27384
rect 13780 27344 13786 27356
rect 14369 27353 14381 27356
rect 14415 27353 14427 27387
rect 14369 27347 14427 27353
rect 14936 27316 14964 27415
rect 15948 27384 15976 27415
rect 16022 27412 16028 27464
rect 16080 27452 16086 27464
rect 16209 27455 16267 27461
rect 16080 27424 16125 27452
rect 16080 27412 16086 27424
rect 16209 27421 16221 27455
rect 16255 27452 16267 27455
rect 18230 27452 18236 27464
rect 16255 27424 18092 27452
rect 18191 27424 18236 27452
rect 16255 27421 16267 27424
rect 16209 27415 16267 27421
rect 16298 27384 16304 27396
rect 15948 27356 16304 27384
rect 16298 27344 16304 27356
rect 16356 27344 16362 27396
rect 16393 27387 16451 27393
rect 16393 27353 16405 27387
rect 16439 27384 16451 27387
rect 17966 27387 18024 27393
rect 17966 27384 17978 27387
rect 16439 27356 17978 27384
rect 16439 27353 16451 27356
rect 16393 27347 16451 27353
rect 17966 27353 17978 27356
rect 18012 27353 18024 27387
rect 18064 27384 18092 27424
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 21174 27412 21180 27464
rect 21232 27452 21238 27464
rect 22296 27461 22324 27492
rect 25866 27480 25872 27532
rect 25924 27520 25930 27532
rect 28445 27523 28503 27529
rect 28445 27520 28457 27523
rect 25924 27492 26740 27520
rect 25924 27480 25930 27492
rect 22005 27455 22063 27461
rect 22005 27452 22017 27455
rect 21232 27424 22017 27452
rect 21232 27412 21238 27424
rect 22005 27421 22017 27424
rect 22051 27421 22063 27455
rect 22005 27415 22063 27421
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27452 25467 27455
rect 25682 27452 25688 27464
rect 25455 27424 25544 27452
rect 25643 27424 25688 27452
rect 25455 27421 25467 27424
rect 25409 27415 25467 27421
rect 19518 27384 19524 27396
rect 18064 27356 19524 27384
rect 17966 27347 18024 27353
rect 19518 27344 19524 27356
rect 19576 27384 19582 27396
rect 20990 27384 20996 27396
rect 19576 27356 20996 27384
rect 19576 27344 19582 27356
rect 20990 27344 20996 27356
rect 21048 27344 21054 27396
rect 19794 27316 19800 27328
rect 14936 27288 19800 27316
rect 19794 27276 19800 27288
rect 19852 27276 19858 27328
rect 21910 27276 21916 27328
rect 21968 27316 21974 27328
rect 22097 27319 22155 27325
rect 22097 27316 22109 27319
rect 21968 27288 22109 27316
rect 21968 27276 21974 27288
rect 22097 27285 22109 27288
rect 22143 27285 22155 27319
rect 22097 27279 22155 27285
rect 22370 27276 22376 27328
rect 22428 27316 22434 27328
rect 22465 27319 22523 27325
rect 22465 27316 22477 27319
rect 22428 27288 22477 27316
rect 22428 27276 22434 27288
rect 22465 27285 22477 27288
rect 22511 27285 22523 27319
rect 25516 27316 25544 27424
rect 25682 27412 25688 27424
rect 25740 27412 25746 27464
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 25590 27344 25596 27396
rect 25648 27384 25654 27396
rect 26068 27384 26096 27415
rect 26142 27412 26148 27464
rect 26200 27452 26206 27464
rect 26712 27461 26740 27492
rect 27724 27492 28457 27520
rect 27724 27464 27752 27492
rect 28445 27489 28457 27492
rect 28491 27489 28503 27523
rect 28445 27483 28503 27489
rect 26329 27455 26387 27461
rect 26329 27452 26341 27455
rect 26200 27424 26341 27452
rect 26200 27412 26206 27424
rect 26329 27421 26341 27424
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26697 27455 26755 27461
rect 26697 27421 26709 27455
rect 26743 27421 26755 27455
rect 26697 27415 26755 27421
rect 27433 27455 27491 27461
rect 27433 27421 27445 27455
rect 27479 27421 27491 27455
rect 27706 27452 27712 27464
rect 27667 27424 27712 27452
rect 27433 27415 27491 27421
rect 26234 27384 26240 27396
rect 25648 27356 26240 27384
rect 25648 27344 25654 27356
rect 26234 27344 26240 27356
rect 26292 27344 26298 27396
rect 26344 27384 26372 27415
rect 27448 27384 27476 27415
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 28166 27412 28172 27464
rect 28224 27452 28230 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 28224 27424 28365 27452
rect 28224 27412 28230 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 28353 27415 28411 27421
rect 28537 27455 28595 27461
rect 28537 27421 28549 27455
rect 28583 27421 28595 27455
rect 28537 27415 28595 27421
rect 29825 27455 29883 27461
rect 29825 27421 29837 27455
rect 29871 27452 29883 27455
rect 29914 27452 29920 27464
rect 29871 27424 29920 27452
rect 29871 27421 29883 27424
rect 29825 27415 29883 27421
rect 26344 27356 27476 27384
rect 25774 27316 25780 27328
rect 25516 27288 25780 27316
rect 22465 27279 22523 27285
rect 25774 27276 25780 27288
rect 25832 27316 25838 27328
rect 26694 27316 26700 27328
rect 25832 27288 26700 27316
rect 25832 27276 25838 27288
rect 26694 27276 26700 27288
rect 26752 27276 26758 27328
rect 27062 27276 27068 27328
rect 27120 27316 27126 27328
rect 27525 27319 27583 27325
rect 27525 27316 27537 27319
rect 27120 27288 27537 27316
rect 27120 27276 27126 27288
rect 27525 27285 27537 27288
rect 27571 27285 27583 27319
rect 28552 27316 28580 27415
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 30092 27387 30150 27393
rect 30092 27353 30104 27387
rect 30138 27384 30150 27387
rect 32214 27384 32220 27396
rect 30138 27356 32220 27384
rect 30138 27353 30150 27356
rect 30092 27347 30150 27353
rect 32214 27344 32220 27356
rect 32272 27344 32278 27396
rect 28718 27316 28724 27328
rect 28552 27288 28724 27316
rect 27525 27279 27583 27285
rect 28718 27276 28724 27288
rect 28776 27316 28782 27328
rect 31202 27316 31208 27328
rect 28776 27288 31208 27316
rect 28776 27276 28782 27288
rect 31202 27276 31208 27288
rect 31260 27276 31266 27328
rect 1104 27226 35027 27248
rect 1104 27174 9390 27226
rect 9442 27174 9454 27226
rect 9506 27174 9518 27226
rect 9570 27174 9582 27226
rect 9634 27174 9646 27226
rect 9698 27174 17831 27226
rect 17883 27174 17895 27226
rect 17947 27174 17959 27226
rect 18011 27174 18023 27226
rect 18075 27174 18087 27226
rect 18139 27174 26272 27226
rect 26324 27174 26336 27226
rect 26388 27174 26400 27226
rect 26452 27174 26464 27226
rect 26516 27174 26528 27226
rect 26580 27174 34713 27226
rect 34765 27174 34777 27226
rect 34829 27174 34841 27226
rect 34893 27174 34905 27226
rect 34957 27174 34969 27226
rect 35021 27174 35027 27226
rect 1104 27152 35027 27174
rect 12069 27115 12127 27121
rect 12069 27081 12081 27115
rect 12115 27112 12127 27115
rect 12894 27112 12900 27124
rect 12115 27084 12900 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12894 27072 12900 27084
rect 12952 27072 12958 27124
rect 18230 27072 18236 27124
rect 18288 27112 18294 27124
rect 19521 27115 19579 27121
rect 19521 27112 19533 27115
rect 18288 27084 19533 27112
rect 18288 27072 18294 27084
rect 19521 27081 19533 27084
rect 19567 27081 19579 27115
rect 19521 27075 19579 27081
rect 21177 27115 21235 27121
rect 21177 27081 21189 27115
rect 21223 27112 21235 27115
rect 25222 27112 25228 27124
rect 21223 27084 25228 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 8297 27047 8355 27053
rect 8297 27013 8309 27047
rect 8343 27044 8355 27047
rect 9122 27044 9128 27056
rect 8343 27016 9128 27044
rect 8343 27013 8355 27016
rect 8297 27007 8355 27013
rect 9122 27004 9128 27016
rect 9180 27044 9186 27056
rect 10318 27044 10324 27056
rect 9180 27016 10324 27044
rect 9180 27004 9186 27016
rect 10318 27004 10324 27016
rect 10376 27004 10382 27056
rect 12618 27044 12624 27056
rect 11900 27016 12624 27044
rect 8202 26976 8208 26988
rect 8163 26948 8208 26976
rect 8202 26936 8208 26948
rect 8260 26936 8266 26988
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 9217 26979 9275 26985
rect 9217 26976 9229 26979
rect 8527 26948 9229 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 9217 26945 9229 26948
rect 9263 26976 9275 26979
rect 9766 26976 9772 26988
rect 9263 26948 9772 26976
rect 9263 26945 9275 26948
rect 9217 26939 9275 26945
rect 9766 26936 9772 26948
rect 9824 26936 9830 26988
rect 11900 26985 11928 27016
rect 12618 27004 12624 27016
rect 12676 27004 12682 27056
rect 13814 27004 13820 27056
rect 13872 27044 13878 27056
rect 14274 27044 14280 27056
rect 13872 27016 14280 27044
rect 13872 27004 13878 27016
rect 14274 27004 14280 27016
rect 14332 27044 14338 27056
rect 15473 27047 15531 27053
rect 15473 27044 15485 27047
rect 14332 27016 15485 27044
rect 14332 27004 14338 27016
rect 15473 27013 15485 27016
rect 15519 27013 15531 27047
rect 15473 27007 15531 27013
rect 19794 27004 19800 27056
rect 19852 27044 19858 27056
rect 22664 27053 22692 27084
rect 25222 27072 25228 27084
rect 25280 27112 25286 27124
rect 25498 27112 25504 27124
rect 25280 27084 25504 27112
rect 25280 27072 25286 27084
rect 25498 27072 25504 27084
rect 25556 27072 25562 27124
rect 31110 27112 31116 27124
rect 31071 27084 31116 27112
rect 31110 27072 31116 27084
rect 31168 27072 31174 27124
rect 22649 27047 22707 27053
rect 19852 27016 22140 27044
rect 19852 27004 19858 27016
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 12161 26979 12219 26985
rect 12161 26945 12173 26979
rect 12207 26976 12219 26979
rect 12434 26976 12440 26988
rect 12207 26948 12440 26976
rect 12207 26945 12219 26948
rect 12161 26939 12219 26945
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 13446 26936 13452 26988
rect 13504 26976 13510 26988
rect 13722 26976 13728 26988
rect 13504 26948 13728 26976
rect 13504 26936 13510 26948
rect 13722 26936 13728 26948
rect 13780 26936 13786 26988
rect 15657 26979 15715 26985
rect 15657 26945 15669 26979
rect 15703 26945 15715 26979
rect 15657 26939 15715 26945
rect 9033 26911 9091 26917
rect 9033 26877 9045 26911
rect 9079 26877 9091 26911
rect 9033 26871 9091 26877
rect 8481 26843 8539 26849
rect 8481 26809 8493 26843
rect 8527 26840 8539 26843
rect 9048 26840 9076 26871
rect 9122 26868 9128 26920
rect 9180 26908 9186 26920
rect 9309 26911 9367 26917
rect 9180 26880 9225 26908
rect 9180 26868 9186 26880
rect 9309 26877 9321 26911
rect 9355 26877 9367 26911
rect 15672 26908 15700 26939
rect 15746 26936 15752 26988
rect 15804 26976 15810 26988
rect 16390 26976 16396 26988
rect 15804 26948 16396 26976
rect 15804 26936 15810 26948
rect 16390 26936 16396 26948
rect 16448 26936 16454 26988
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18322 26976 18328 26988
rect 18279 26948 18328 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18322 26936 18328 26948
rect 18380 26936 18386 26988
rect 20990 26976 20996 26988
rect 20951 26948 20996 26976
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 21174 26936 21180 26988
rect 21232 26976 21238 26988
rect 22112 26985 22140 27016
rect 22649 27013 22661 27047
rect 22695 27044 22707 27047
rect 26142 27044 26148 27056
rect 22695 27016 22729 27044
rect 25700 27016 26148 27044
rect 22695 27013 22707 27016
rect 22649 27007 22707 27013
rect 21269 26979 21327 26985
rect 21269 26976 21281 26979
rect 21232 26948 21281 26976
rect 21232 26936 21238 26948
rect 21269 26945 21281 26948
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 22097 26939 22155 26945
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24949 26979 25007 26985
rect 24949 26976 24961 26979
rect 24820 26948 24961 26976
rect 24820 26936 24826 26948
rect 24949 26945 24961 26948
rect 24995 26945 25007 26979
rect 25130 26976 25136 26988
rect 25091 26948 25136 26976
rect 24949 26939 25007 26945
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 25590 26976 25596 26988
rect 25551 26948 25596 26976
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 25700 26985 25728 27016
rect 26142 27004 26148 27016
rect 26200 27044 26206 27056
rect 27525 27047 27583 27053
rect 27525 27044 27537 27047
rect 26200 27016 27537 27044
rect 26200 27004 26206 27016
rect 27525 27013 27537 27016
rect 27571 27013 27583 27047
rect 27525 27007 27583 27013
rect 25685 26979 25743 26985
rect 25685 26945 25697 26979
rect 25731 26945 25743 26979
rect 25866 26976 25872 26988
rect 25827 26948 25872 26976
rect 25685 26939 25743 26945
rect 25866 26936 25872 26948
rect 25924 26936 25930 26988
rect 27246 26976 27252 26988
rect 27207 26948 27252 26976
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27430 26976 27436 26988
rect 27391 26948 27436 26976
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 30006 26976 30012 26988
rect 29967 26948 30012 26976
rect 30006 26936 30012 26948
rect 30064 26936 30070 26988
rect 16666 26908 16672 26920
rect 15672 26880 16672 26908
rect 9309 26871 9367 26877
rect 9324 26840 9352 26871
rect 16666 26868 16672 26880
rect 16724 26868 16730 26920
rect 26142 26868 26148 26920
rect 26200 26908 26206 26920
rect 26421 26911 26479 26917
rect 26421 26908 26433 26911
rect 26200 26880 26433 26908
rect 26200 26868 26206 26880
rect 26421 26877 26433 26880
rect 26467 26908 26479 26911
rect 27614 26908 27620 26920
rect 26467 26880 27620 26908
rect 26467 26877 26479 26880
rect 26421 26871 26479 26877
rect 27614 26868 27620 26880
rect 27672 26868 27678 26920
rect 29733 26911 29791 26917
rect 29733 26877 29745 26911
rect 29779 26908 29791 26911
rect 29914 26908 29920 26920
rect 29779 26880 29920 26908
rect 29779 26877 29791 26880
rect 29733 26871 29791 26877
rect 29914 26868 29920 26880
rect 29972 26868 29978 26920
rect 8527 26812 9076 26840
rect 9140 26812 9352 26840
rect 8527 26809 8539 26812
rect 8481 26803 8539 26809
rect 8754 26732 8760 26784
rect 8812 26772 8818 26784
rect 9140 26772 9168 26812
rect 8812 26744 9168 26772
rect 8812 26732 8818 26744
rect 9214 26732 9220 26784
rect 9272 26772 9278 26784
rect 9493 26775 9551 26781
rect 9493 26772 9505 26775
rect 9272 26744 9505 26772
rect 9272 26732 9278 26744
rect 9493 26741 9505 26744
rect 9539 26741 9551 26775
rect 9493 26735 9551 26741
rect 11146 26732 11152 26784
rect 11204 26772 11210 26784
rect 11701 26775 11759 26781
rect 11701 26772 11713 26775
rect 11204 26744 11713 26772
rect 11204 26732 11210 26744
rect 11701 26741 11713 26744
rect 11747 26741 11759 26775
rect 11701 26735 11759 26741
rect 12618 26732 12624 26784
rect 12676 26772 12682 26784
rect 13633 26775 13691 26781
rect 13633 26772 13645 26775
rect 12676 26744 13645 26772
rect 12676 26732 12682 26744
rect 13633 26741 13645 26744
rect 13679 26772 13691 26775
rect 20530 26772 20536 26784
rect 13679 26744 20536 26772
rect 13679 26741 13691 26744
rect 13633 26735 13691 26741
rect 20530 26732 20536 26744
rect 20588 26732 20594 26784
rect 20809 26775 20867 26781
rect 20809 26741 20821 26775
rect 20855 26772 20867 26775
rect 20898 26772 20904 26784
rect 20855 26744 20904 26772
rect 20855 26741 20867 26744
rect 20809 26735 20867 26741
rect 20898 26732 20904 26744
rect 20956 26732 20962 26784
rect 1104 26682 34868 26704
rect 1104 26630 5170 26682
rect 5222 26630 5234 26682
rect 5286 26630 5298 26682
rect 5350 26630 5362 26682
rect 5414 26630 5426 26682
rect 5478 26630 13611 26682
rect 13663 26630 13675 26682
rect 13727 26630 13739 26682
rect 13791 26630 13803 26682
rect 13855 26630 13867 26682
rect 13919 26630 22052 26682
rect 22104 26630 22116 26682
rect 22168 26630 22180 26682
rect 22232 26630 22244 26682
rect 22296 26630 22308 26682
rect 22360 26630 30493 26682
rect 30545 26630 30557 26682
rect 30609 26630 30621 26682
rect 30673 26630 30685 26682
rect 30737 26630 30749 26682
rect 30801 26630 34868 26682
rect 1104 26608 34868 26630
rect 12345 26571 12403 26577
rect 12345 26537 12357 26571
rect 12391 26568 12403 26571
rect 12434 26568 12440 26580
rect 12391 26540 12440 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 13354 26568 13360 26580
rect 12952 26540 13360 26568
rect 12952 26528 12958 26540
rect 13354 26528 13360 26540
rect 13412 26568 13418 26580
rect 13449 26571 13507 26577
rect 13449 26568 13461 26571
rect 13412 26540 13461 26568
rect 13412 26528 13418 26540
rect 13449 26537 13461 26540
rect 13495 26537 13507 26571
rect 16666 26568 16672 26580
rect 16627 26540 16672 26568
rect 13449 26531 13507 26537
rect 16666 26528 16672 26540
rect 16724 26528 16730 26580
rect 25130 26528 25136 26580
rect 25188 26568 25194 26580
rect 25225 26571 25283 26577
rect 25225 26568 25237 26571
rect 25188 26540 25237 26568
rect 25188 26528 25194 26540
rect 25225 26537 25237 26540
rect 25271 26537 25283 26571
rect 27062 26568 27068 26580
rect 27023 26540 27068 26568
rect 25225 26531 25283 26537
rect 27062 26528 27068 26540
rect 27120 26528 27126 26580
rect 32214 26568 32220 26580
rect 32175 26540 32220 26568
rect 32214 26528 32220 26540
rect 32272 26528 32278 26580
rect 9306 26460 9312 26512
rect 9364 26500 9370 26512
rect 9401 26503 9459 26509
rect 9401 26500 9413 26503
rect 9364 26472 9413 26500
rect 9364 26460 9370 26472
rect 9401 26469 9413 26472
rect 9447 26469 9459 26503
rect 13265 26503 13323 26509
rect 13265 26500 13277 26503
rect 9401 26463 9459 26469
rect 12084 26472 13277 26500
rect 11146 26432 11152 26444
rect 11107 26404 11152 26432
rect 11146 26392 11152 26404
rect 11204 26392 11210 26444
rect 11701 26435 11759 26441
rect 11701 26401 11713 26435
rect 11747 26432 11759 26435
rect 12084 26432 12112 26472
rect 13265 26469 13277 26472
rect 13311 26469 13323 26503
rect 13265 26463 13323 26469
rect 18966 26460 18972 26512
rect 19024 26500 19030 26512
rect 21174 26500 21180 26512
rect 19024 26472 21180 26500
rect 19024 26460 19030 26472
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 11747 26404 12112 26432
rect 12406 26404 12725 26432
rect 11747 26401 11759 26404
rect 11701 26395 11759 26401
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 12406 26364 12434 26404
rect 12713 26401 12725 26404
rect 12759 26432 12771 26435
rect 12802 26432 12808 26444
rect 12759 26404 12808 26432
rect 12759 26401 12771 26404
rect 12713 26395 12771 26401
rect 12802 26392 12808 26404
rect 12860 26392 12866 26444
rect 13446 26392 13452 26444
rect 13504 26432 13510 26444
rect 18049 26435 18107 26441
rect 13504 26404 13676 26432
rect 13504 26392 13510 26404
rect 12618 26364 12624 26376
rect 11379 26336 12434 26364
rect 12579 26336 12624 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 9030 26256 9036 26308
rect 9088 26296 9094 26308
rect 9125 26299 9183 26305
rect 9125 26296 9137 26299
rect 9088 26268 9137 26296
rect 9088 26256 9094 26268
rect 9125 26265 9137 26268
rect 9171 26296 9183 26299
rect 11609 26299 11667 26305
rect 11609 26296 11621 26299
rect 9171 26268 11621 26296
rect 9171 26265 9183 26268
rect 9125 26259 9183 26265
rect 11609 26265 11621 26268
rect 11655 26265 11667 26299
rect 11609 26259 11667 26265
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13446 26305 13452 26308
rect 13417 26299 13452 26305
rect 13417 26296 13429 26299
rect 12584 26268 13429 26296
rect 12584 26256 12590 26268
rect 13417 26265 13429 26268
rect 13504 26296 13510 26308
rect 13648 26305 13676 26404
rect 18049 26401 18061 26435
rect 18095 26432 18107 26435
rect 18230 26432 18236 26444
rect 18095 26404 18236 26432
rect 18095 26401 18107 26404
rect 18049 26395 18107 26401
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19392 26404 19840 26432
rect 19392 26392 19398 26404
rect 19812 26373 19840 26404
rect 19904 26373 19932 26472
rect 21174 26460 21180 26472
rect 21232 26460 21238 26512
rect 22738 26460 22744 26512
rect 22796 26500 22802 26512
rect 22796 26472 25728 26500
rect 22796 26460 22802 26472
rect 25498 26432 25504 26444
rect 25459 26404 25504 26432
rect 25498 26392 25504 26404
rect 25556 26392 25562 26444
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26333 19855 26367
rect 19797 26327 19855 26333
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26333 19947 26367
rect 19889 26327 19947 26333
rect 13633 26299 13691 26305
rect 13504 26268 13565 26296
rect 13417 26259 13452 26265
rect 13446 26256 13452 26259
rect 13504 26256 13510 26268
rect 13633 26265 13645 26299
rect 13679 26265 13691 26299
rect 13633 26259 13691 26265
rect 16850 26256 16856 26308
rect 16908 26296 16914 26308
rect 17782 26299 17840 26305
rect 17782 26296 17794 26299
rect 16908 26268 17794 26296
rect 16908 26256 16914 26268
rect 17782 26265 17794 26268
rect 17828 26265 17840 26299
rect 17782 26259 17840 26265
rect 18230 26256 18236 26308
rect 18288 26296 18294 26308
rect 19429 26299 19487 26305
rect 19429 26296 19441 26299
rect 18288 26268 19441 26296
rect 18288 26256 18294 26268
rect 19429 26265 19441 26268
rect 19475 26265 19487 26299
rect 19628 26296 19656 26327
rect 24854 26324 24860 26376
rect 24912 26364 24918 26376
rect 25314 26364 25320 26376
rect 24912 26336 25320 26364
rect 24912 26324 24918 26336
rect 25314 26324 25320 26336
rect 25372 26364 25378 26376
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 25372 26336 25421 26364
rect 25372 26324 25378 26336
rect 25409 26333 25421 26336
rect 25455 26333 25467 26367
rect 25590 26364 25596 26376
rect 25551 26336 25596 26364
rect 25409 26327 25467 26333
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 25700 26373 25728 26472
rect 26510 26460 26516 26512
rect 26568 26500 26574 26512
rect 26786 26500 26792 26512
rect 26568 26472 26792 26500
rect 26568 26460 26574 26472
rect 26786 26460 26792 26472
rect 26844 26500 26850 26512
rect 26844 26472 27752 26500
rect 26844 26460 26850 26472
rect 27724 26441 27752 26472
rect 28626 26460 28632 26512
rect 28684 26500 28690 26512
rect 31297 26503 31355 26509
rect 31297 26500 31309 26503
rect 28684 26472 31309 26500
rect 28684 26460 28690 26472
rect 31297 26469 31309 26472
rect 31343 26469 31355 26503
rect 31297 26463 31355 26469
rect 27709 26435 27767 26441
rect 25792 26404 27568 26432
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 22554 26296 22560 26308
rect 19628 26268 19932 26296
rect 22515 26268 22560 26296
rect 19429 26259 19487 26265
rect 19904 26240 19932 26268
rect 22554 26256 22560 26268
rect 22612 26256 22618 26308
rect 24578 26256 24584 26308
rect 24636 26296 24642 26308
rect 25792 26296 25820 26404
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26364 25927 26367
rect 26510 26364 26516 26376
rect 25915 26336 26372 26364
rect 26471 26336 26516 26364
rect 25915 26333 25927 26336
rect 25869 26327 25927 26333
rect 24636 26268 25820 26296
rect 24636 26256 24642 26268
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 9585 26231 9643 26237
rect 9585 26228 9597 26231
rect 9364 26200 9597 26228
rect 9364 26188 9370 26200
rect 9585 26197 9597 26200
rect 9631 26197 9643 26231
rect 9585 26191 9643 26197
rect 19886 26188 19892 26240
rect 19944 26188 19950 26240
rect 21085 26231 21143 26237
rect 21085 26197 21097 26231
rect 21131 26228 21143 26231
rect 21174 26228 21180 26240
rect 21131 26200 21180 26228
rect 21131 26197 21143 26200
rect 21085 26191 21143 26197
rect 21174 26188 21180 26200
rect 21232 26188 21238 26240
rect 26344 26228 26372 26336
rect 26510 26324 26516 26336
rect 26568 26324 26574 26376
rect 26602 26324 26608 26376
rect 26660 26364 26666 26376
rect 26896 26373 27016 26374
rect 26789 26367 26847 26373
rect 26660 26336 26705 26364
rect 26660 26324 26666 26336
rect 26789 26333 26801 26367
rect 26835 26333 26847 26367
rect 26789 26327 26847 26333
rect 26881 26367 27016 26373
rect 26881 26333 26893 26367
rect 26927 26364 27016 26367
rect 27154 26364 27160 26376
rect 26927 26346 27160 26364
rect 26927 26333 26939 26346
rect 26988 26336 27160 26346
rect 26881 26327 26939 26333
rect 26804 26296 26832 26327
rect 27154 26324 27160 26336
rect 27212 26324 27218 26376
rect 27540 26373 27568 26404
rect 27709 26401 27721 26435
rect 27755 26401 27767 26435
rect 27709 26395 27767 26401
rect 27525 26367 27583 26373
rect 27525 26333 27537 26367
rect 27571 26333 27583 26367
rect 32398 26364 32404 26376
rect 32359 26336 32404 26364
rect 27525 26327 27583 26333
rect 32398 26324 32404 26336
rect 32456 26324 32462 26376
rect 32674 26364 32680 26376
rect 32635 26336 32680 26364
rect 32674 26324 32680 26336
rect 32732 26324 32738 26376
rect 26804 26268 26921 26296
rect 26602 26228 26608 26240
rect 26344 26200 26608 26228
rect 26602 26188 26608 26200
rect 26660 26188 26666 26240
rect 26893 26228 26921 26268
rect 29086 26256 29092 26308
rect 29144 26296 29150 26308
rect 30009 26299 30067 26305
rect 30009 26296 30021 26299
rect 29144 26268 30021 26296
rect 29144 26256 29150 26268
rect 30009 26265 30021 26268
rect 30055 26265 30067 26299
rect 30009 26259 30067 26265
rect 31202 26256 31208 26308
rect 31260 26296 31266 26308
rect 32585 26299 32643 26305
rect 32585 26296 32597 26299
rect 31260 26268 32597 26296
rect 31260 26256 31266 26268
rect 32585 26265 32597 26268
rect 32631 26265 32643 26299
rect 32585 26259 32643 26265
rect 27522 26228 27528 26240
rect 26893 26200 27528 26228
rect 27522 26188 27528 26200
rect 27580 26188 27586 26240
rect 1104 26138 35027 26160
rect 1104 26086 9390 26138
rect 9442 26086 9454 26138
rect 9506 26086 9518 26138
rect 9570 26086 9582 26138
rect 9634 26086 9646 26138
rect 9698 26086 17831 26138
rect 17883 26086 17895 26138
rect 17947 26086 17959 26138
rect 18011 26086 18023 26138
rect 18075 26086 18087 26138
rect 18139 26086 26272 26138
rect 26324 26086 26336 26138
rect 26388 26086 26400 26138
rect 26452 26086 26464 26138
rect 26516 26086 26528 26138
rect 26580 26086 34713 26138
rect 34765 26086 34777 26138
rect 34829 26086 34841 26138
rect 34893 26086 34905 26138
rect 34957 26086 34969 26138
rect 35021 26086 35027 26138
rect 1104 26064 35027 26086
rect 12253 26027 12311 26033
rect 12253 25993 12265 26027
rect 12299 26024 12311 26027
rect 12526 26024 12532 26036
rect 12299 25996 12532 26024
rect 12299 25993 12311 25996
rect 12253 25987 12311 25993
rect 12526 25984 12532 25996
rect 12584 25984 12590 26036
rect 14734 26024 14740 26036
rect 13188 25996 14740 26024
rect 10505 25959 10563 25965
rect 10505 25956 10517 25959
rect 9508 25928 10517 25956
rect 9306 25848 9312 25900
rect 9364 25888 9370 25900
rect 9508 25897 9536 25928
rect 10505 25925 10517 25928
rect 10551 25925 10563 25959
rect 12342 25956 12348 25968
rect 12303 25928 12348 25956
rect 10505 25919 10563 25925
rect 12342 25916 12348 25928
rect 12400 25916 12406 25968
rect 12434 25916 12440 25968
rect 12492 25956 12498 25968
rect 13081 25959 13139 25965
rect 13081 25956 13093 25959
rect 12492 25928 13093 25956
rect 12492 25916 12498 25928
rect 13081 25925 13093 25928
rect 13127 25925 13139 25959
rect 13081 25919 13139 25925
rect 9493 25891 9551 25897
rect 9493 25888 9505 25891
rect 9364 25860 9505 25888
rect 9364 25848 9370 25860
rect 9493 25857 9505 25860
rect 9539 25857 9551 25891
rect 9493 25851 9551 25857
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25857 9827 25891
rect 10413 25891 10471 25897
rect 10413 25888 10425 25891
rect 9769 25851 9827 25857
rect 9876 25860 10425 25888
rect 9214 25780 9220 25832
rect 9272 25820 9278 25832
rect 9582 25820 9588 25832
rect 9272 25792 9588 25820
rect 9272 25780 9278 25792
rect 9582 25780 9588 25792
rect 9640 25780 9646 25832
rect 9784 25684 9812 25851
rect 9876 25832 9904 25860
rect 10413 25857 10425 25860
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 10689 25891 10747 25897
rect 10689 25857 10701 25891
rect 10735 25888 10747 25891
rect 12250 25888 12256 25900
rect 10735 25860 12256 25888
rect 10735 25857 10747 25860
rect 10689 25851 10747 25857
rect 12250 25848 12256 25860
rect 12308 25848 12314 25900
rect 12360 25888 12388 25916
rect 13188 25888 13216 25996
rect 14734 25984 14740 25996
rect 14792 25984 14798 26036
rect 16850 26024 16856 26036
rect 16811 25996 16856 26024
rect 16850 25984 16856 25996
rect 16908 25984 16914 26036
rect 25038 26024 25044 26036
rect 24504 25996 25044 26024
rect 13354 25956 13360 25968
rect 13315 25928 13360 25956
rect 13354 25916 13360 25928
rect 13412 25916 13418 25968
rect 16666 25916 16672 25968
rect 16724 25956 16730 25968
rect 17221 25959 17279 25965
rect 17221 25956 17233 25959
rect 16724 25928 17233 25956
rect 16724 25916 16730 25928
rect 17221 25925 17233 25928
rect 17267 25925 17279 25959
rect 17221 25919 17279 25925
rect 21361 25959 21419 25965
rect 21361 25925 21373 25959
rect 21407 25956 21419 25959
rect 21910 25956 21916 25968
rect 21407 25928 21916 25956
rect 21407 25925 21419 25928
rect 21361 25919 21419 25925
rect 21910 25916 21916 25928
rect 21968 25916 21974 25968
rect 13265 25891 13323 25897
rect 13265 25888 13277 25891
rect 12360 25860 13277 25888
rect 13265 25857 13277 25860
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 9858 25780 9864 25832
rect 9916 25780 9922 25832
rect 12069 25823 12127 25829
rect 12069 25789 12081 25823
rect 12115 25820 12127 25823
rect 13372 25820 13400 25916
rect 13446 25848 13452 25900
rect 13504 25897 13510 25900
rect 13504 25888 13512 25897
rect 17034 25888 17040 25900
rect 13504 25860 13549 25888
rect 16995 25860 17040 25888
rect 13504 25851 13512 25860
rect 13504 25848 13510 25851
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 17313 25891 17371 25897
rect 17313 25857 17325 25891
rect 17359 25857 17371 25891
rect 19610 25888 19616 25900
rect 19571 25860 19616 25888
rect 17313 25851 17371 25857
rect 12115 25792 13400 25820
rect 12115 25789 12127 25792
rect 12069 25783 12127 25789
rect 16298 25780 16304 25832
rect 16356 25820 16362 25832
rect 16482 25820 16488 25832
rect 16356 25792 16488 25820
rect 16356 25780 16362 25792
rect 16482 25780 16488 25792
rect 16540 25820 16546 25832
rect 17328 25820 17356 25851
rect 19610 25848 19616 25860
rect 19668 25848 19674 25900
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25857 20867 25891
rect 20809 25851 20867 25857
rect 16540 25792 17356 25820
rect 16540 25780 16546 25792
rect 9953 25755 10011 25761
rect 9953 25721 9965 25755
rect 9999 25752 10011 25755
rect 14458 25752 14464 25764
rect 9999 25724 14464 25752
rect 9999 25721 10011 25724
rect 9953 25715 10011 25721
rect 14458 25712 14464 25724
rect 14516 25712 14522 25764
rect 20824 25752 20852 25851
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21232 25860 22017 25888
rect 21232 25848 21238 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25888 22339 25891
rect 22370 25888 22376 25900
rect 22327 25860 22376 25888
rect 22327 25857 22339 25860
rect 22281 25851 22339 25857
rect 22370 25848 22376 25860
rect 22428 25848 22434 25900
rect 24504 25897 24532 25996
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 25593 26027 25651 26033
rect 25593 25993 25605 26027
rect 25639 26024 25651 26027
rect 25682 26024 25688 26036
rect 25639 25996 25688 26024
rect 25639 25993 25651 25996
rect 25593 25987 25651 25993
rect 25682 25984 25688 25996
rect 25740 25984 25746 26036
rect 27157 26027 27215 26033
rect 27157 25993 27169 26027
rect 27203 26024 27215 26027
rect 27246 26024 27252 26036
rect 27203 25996 27252 26024
rect 27203 25993 27215 25996
rect 27157 25987 27215 25993
rect 27246 25984 27252 25996
rect 27304 25984 27310 26036
rect 29914 26024 29920 26036
rect 29875 25996 29920 26024
rect 29914 25984 29920 25996
rect 29972 25984 29978 26036
rect 24581 25959 24639 25965
rect 24581 25925 24593 25959
rect 24627 25956 24639 25959
rect 25133 25959 25191 25965
rect 25133 25956 25145 25959
rect 24627 25928 25145 25956
rect 24627 25925 24639 25928
rect 24581 25919 24639 25925
rect 25133 25925 25145 25928
rect 25179 25956 25191 25959
rect 25498 25956 25504 25968
rect 25179 25928 25504 25956
rect 25179 25925 25191 25928
rect 25133 25919 25191 25925
rect 25498 25916 25504 25928
rect 25556 25916 25562 25968
rect 28626 25956 28632 25968
rect 28587 25928 28632 25956
rect 28626 25916 28632 25928
rect 28684 25916 28690 25968
rect 31478 25916 31484 25968
rect 31536 25956 31542 25968
rect 32677 25959 32735 25965
rect 32677 25956 32689 25959
rect 31536 25928 32689 25956
rect 31536 25916 31542 25928
rect 32677 25925 32689 25928
rect 32723 25925 32735 25959
rect 32677 25919 32735 25925
rect 24489 25891 24547 25897
rect 24489 25857 24501 25891
rect 24535 25857 24547 25891
rect 24670 25888 24676 25900
rect 24631 25860 24676 25888
rect 24489 25851 24547 25857
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 26510 25888 26516 25900
rect 26471 25860 26516 25888
rect 26510 25848 26516 25860
rect 26568 25848 26574 25900
rect 27614 25888 27620 25900
rect 27575 25860 27620 25888
rect 27614 25848 27620 25860
rect 27672 25848 27678 25900
rect 31938 25848 31944 25900
rect 31996 25888 32002 25900
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 31996 25860 32505 25888
rect 31996 25848 32002 25860
rect 32493 25857 32505 25860
rect 32539 25857 32551 25891
rect 32766 25888 32772 25900
rect 32727 25860 32772 25888
rect 32493 25851 32551 25857
rect 32766 25848 32772 25860
rect 32824 25848 32830 25900
rect 23382 25820 23388 25832
rect 21468 25792 23388 25820
rect 21468 25752 21496 25792
rect 23382 25780 23388 25792
rect 23440 25820 23446 25832
rect 23477 25823 23535 25829
rect 23477 25820 23489 25823
rect 23440 25792 23489 25820
rect 23440 25780 23446 25792
rect 23477 25789 23489 25792
rect 23523 25789 23535 25823
rect 23477 25783 23535 25789
rect 26605 25823 26663 25829
rect 26605 25789 26617 25823
rect 26651 25820 26663 25823
rect 26694 25820 26700 25832
rect 26651 25792 26700 25820
rect 26651 25789 26663 25792
rect 26605 25783 26663 25789
rect 26694 25780 26700 25792
rect 26752 25780 26758 25832
rect 27062 25780 27068 25832
rect 27120 25820 27126 25832
rect 27341 25823 27399 25829
rect 27341 25820 27353 25823
rect 27120 25792 27353 25820
rect 27120 25780 27126 25792
rect 27341 25789 27353 25792
rect 27387 25789 27399 25823
rect 27341 25783 27399 25789
rect 27433 25823 27491 25829
rect 27433 25789 27445 25823
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 20824 25724 21496 25752
rect 25038 25712 25044 25764
rect 25096 25752 25102 25764
rect 25409 25755 25467 25761
rect 25409 25752 25421 25755
rect 25096 25724 25421 25752
rect 25096 25712 25102 25724
rect 25409 25721 25421 25724
rect 25455 25752 25467 25755
rect 27154 25752 27160 25764
rect 25455 25724 27160 25752
rect 25455 25721 25467 25724
rect 25409 25715 25467 25721
rect 27154 25712 27160 25724
rect 27212 25752 27218 25764
rect 27448 25752 27476 25783
rect 27522 25780 27528 25832
rect 27580 25820 27586 25832
rect 27580 25792 27625 25820
rect 27580 25780 27586 25792
rect 27212 25724 27476 25752
rect 27212 25712 27218 25724
rect 10689 25687 10747 25693
rect 10689 25684 10701 25687
rect 9784 25656 10701 25684
rect 10689 25653 10701 25656
rect 10735 25653 10747 25687
rect 10689 25647 10747 25653
rect 12621 25687 12679 25693
rect 12621 25653 12633 25687
rect 12667 25684 12679 25687
rect 12710 25684 12716 25696
rect 12667 25656 12716 25684
rect 12667 25653 12679 25656
rect 12621 25647 12679 25653
rect 12710 25644 12716 25656
rect 12768 25644 12774 25696
rect 13078 25684 13084 25696
rect 13039 25656 13084 25684
rect 13078 25644 13084 25656
rect 13136 25644 13142 25696
rect 18322 25684 18328 25696
rect 18283 25656 18328 25684
rect 18322 25644 18328 25656
rect 18380 25644 18386 25696
rect 32306 25684 32312 25696
rect 32267 25656 32312 25684
rect 32306 25644 32312 25656
rect 32364 25644 32370 25696
rect 1104 25594 34868 25616
rect 1104 25542 5170 25594
rect 5222 25542 5234 25594
rect 5286 25542 5298 25594
rect 5350 25542 5362 25594
rect 5414 25542 5426 25594
rect 5478 25542 13611 25594
rect 13663 25542 13675 25594
rect 13727 25542 13739 25594
rect 13791 25542 13803 25594
rect 13855 25542 13867 25594
rect 13919 25542 22052 25594
rect 22104 25542 22116 25594
rect 22168 25542 22180 25594
rect 22232 25542 22244 25594
rect 22296 25542 22308 25594
rect 22360 25542 30493 25594
rect 30545 25542 30557 25594
rect 30609 25542 30621 25594
rect 30673 25542 30685 25594
rect 30737 25542 30749 25594
rect 30801 25542 34868 25594
rect 1104 25520 34868 25542
rect 15381 25483 15439 25489
rect 15381 25449 15393 25483
rect 15427 25480 15439 25483
rect 16666 25480 16672 25492
rect 15427 25452 16672 25480
rect 15427 25449 15439 25452
rect 15381 25443 15439 25449
rect 16298 25412 16304 25424
rect 16259 25384 16304 25412
rect 16298 25372 16304 25384
rect 16356 25372 16362 25424
rect 13078 25344 13084 25356
rect 12544 25316 13084 25344
rect 3326 25236 3332 25288
rect 3384 25276 3390 25288
rect 3421 25279 3479 25285
rect 3421 25276 3433 25279
rect 3384 25248 3433 25276
rect 3384 25236 3390 25248
rect 3421 25245 3433 25248
rect 3467 25245 3479 25279
rect 4062 25276 4068 25288
rect 4023 25248 4068 25276
rect 3421 25239 3479 25245
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 4246 25276 4252 25288
rect 4207 25248 4252 25276
rect 4246 25236 4252 25248
rect 4304 25236 4310 25288
rect 6733 25279 6791 25285
rect 6733 25245 6745 25279
rect 6779 25276 6791 25279
rect 6822 25276 6828 25288
rect 6779 25248 6828 25276
rect 6779 25245 6791 25248
rect 6733 25239 6791 25245
rect 6822 25236 6828 25248
rect 6880 25236 6886 25288
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25276 6975 25279
rect 7834 25276 7840 25288
rect 6963 25248 7840 25276
rect 6963 25245 6975 25248
rect 6917 25239 6975 25245
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 12250 25276 12256 25288
rect 12211 25248 12256 25276
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 12544 25285 12572 25316
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 12710 25276 12716 25288
rect 12671 25248 12716 25276
rect 12529 25239 12587 25245
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 15654 25276 15660 25288
rect 15396 25248 15660 25276
rect 3973 25211 4031 25217
rect 3973 25177 3985 25211
rect 4019 25208 4031 25211
rect 4154 25208 4160 25220
rect 4019 25180 4160 25208
rect 4019 25177 4031 25180
rect 3973 25171 4031 25177
rect 4154 25168 4160 25180
rect 4212 25168 4218 25220
rect 15396 25217 15424 25248
rect 15654 25236 15660 25248
rect 15712 25276 15718 25288
rect 15930 25276 15936 25288
rect 15712 25248 15936 25276
rect 15712 25236 15718 25248
rect 15930 25236 15936 25248
rect 15988 25276 15994 25288
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 15988 25248 16037 25276
rect 15988 25236 15994 25248
rect 16025 25245 16037 25248
rect 16071 25245 16083 25279
rect 16025 25239 16083 25245
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25276 16359 25279
rect 16408 25276 16436 25452
rect 16666 25440 16672 25452
rect 16724 25440 16730 25492
rect 19794 25480 19800 25492
rect 19755 25452 19800 25480
rect 19794 25440 19800 25452
rect 19852 25440 19858 25492
rect 25590 25440 25596 25492
rect 25648 25480 25654 25492
rect 26053 25483 26111 25489
rect 26053 25480 26065 25483
rect 25648 25452 26065 25480
rect 25648 25440 25654 25452
rect 26053 25449 26065 25452
rect 26099 25449 26111 25483
rect 26053 25443 26111 25449
rect 26237 25483 26295 25489
rect 26237 25449 26249 25483
rect 26283 25480 26295 25483
rect 26786 25480 26792 25492
rect 26283 25452 26792 25480
rect 26283 25449 26295 25452
rect 26237 25443 26295 25449
rect 26786 25440 26792 25452
rect 26844 25440 26850 25492
rect 27614 25440 27620 25492
rect 27672 25480 27678 25492
rect 28261 25483 28319 25489
rect 28261 25480 28273 25483
rect 27672 25452 28273 25480
rect 27672 25440 27678 25452
rect 28261 25449 28273 25452
rect 28307 25449 28319 25483
rect 28261 25443 28319 25449
rect 21174 25344 21180 25356
rect 21135 25316 21180 25344
rect 21174 25304 21180 25316
rect 21232 25304 21238 25356
rect 26602 25344 26608 25356
rect 26515 25316 26608 25344
rect 26602 25304 26608 25316
rect 26660 25344 26666 25356
rect 26660 25316 30236 25344
rect 26660 25304 26666 25316
rect 16347 25248 16436 25276
rect 16347 25245 16359 25248
rect 16301 25239 16359 25245
rect 20898 25236 20904 25288
rect 20956 25285 20962 25288
rect 20956 25276 20968 25285
rect 20956 25248 21001 25276
rect 20956 25239 20968 25248
rect 20956 25236 20962 25239
rect 23474 25236 23480 25288
rect 23532 25276 23538 25288
rect 24578 25276 24584 25288
rect 23532 25248 24584 25276
rect 23532 25236 23538 25248
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 24670 25236 24676 25288
rect 24728 25276 24734 25288
rect 24857 25279 24915 25285
rect 24857 25276 24869 25279
rect 24728 25248 24869 25276
rect 24728 25236 24734 25248
rect 24857 25245 24869 25248
rect 24903 25276 24915 25279
rect 27338 25276 27344 25288
rect 24903 25248 27344 25276
rect 24903 25245 24915 25248
rect 24857 25239 24915 25245
rect 27338 25236 27344 25248
rect 27396 25236 27402 25288
rect 28368 25285 28396 25316
rect 27433 25279 27491 25285
rect 27433 25245 27445 25279
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 28353 25279 28411 25285
rect 28353 25245 28365 25279
rect 28399 25245 28411 25279
rect 30098 25276 30104 25288
rect 30059 25248 30104 25276
rect 28353 25239 28411 25245
rect 15365 25211 15424 25217
rect 15365 25177 15377 25211
rect 15411 25180 15424 25211
rect 15411 25177 15423 25180
rect 15365 25171 15423 25177
rect 15470 25168 15476 25220
rect 15528 25208 15534 25220
rect 15565 25211 15623 25217
rect 15565 25208 15577 25211
rect 15528 25180 15577 25208
rect 15528 25168 15534 25180
rect 15565 25177 15577 25180
rect 15611 25177 15623 25211
rect 15565 25171 15623 25177
rect 2866 25100 2872 25152
rect 2924 25140 2930 25152
rect 3329 25143 3387 25149
rect 3329 25140 3341 25143
rect 2924 25112 3341 25140
rect 2924 25100 2930 25112
rect 3329 25109 3341 25112
rect 3375 25109 3387 25143
rect 3329 25103 3387 25109
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 5592 25112 6745 25140
rect 5592 25100 5598 25112
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 6733 25103 6791 25109
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 13446 25140 13452 25152
rect 12115 25112 13452 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 13446 25100 13452 25112
rect 13504 25100 13510 25152
rect 15194 25140 15200 25152
rect 15155 25112 15200 25140
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 15580 25140 15608 25171
rect 21082 25168 21088 25220
rect 21140 25208 21146 25220
rect 21637 25211 21695 25217
rect 21637 25208 21649 25211
rect 21140 25180 21649 25208
rect 21140 25168 21146 25180
rect 21637 25177 21649 25180
rect 21683 25177 21695 25211
rect 21637 25171 21695 25177
rect 25130 25168 25136 25220
rect 25188 25208 25194 25220
rect 26237 25211 26295 25217
rect 26237 25208 26249 25211
rect 25188 25180 26249 25208
rect 25188 25168 25194 25180
rect 26237 25177 26249 25180
rect 26283 25177 26295 25211
rect 26237 25171 26295 25177
rect 26510 25168 26516 25220
rect 26568 25208 26574 25220
rect 27448 25208 27476 25239
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 30208 25276 30236 25316
rect 31478 25276 31484 25288
rect 30208 25248 31484 25276
rect 31478 25236 31484 25248
rect 31536 25236 31542 25288
rect 30374 25217 30380 25220
rect 26568 25180 27476 25208
rect 26568 25168 26574 25180
rect 16114 25140 16120 25152
rect 15580 25112 16120 25140
rect 16114 25100 16120 25112
rect 16172 25100 16178 25152
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 22925 25143 22983 25149
rect 22925 25140 22937 25143
rect 22612 25112 22937 25140
rect 22612 25100 22618 25112
rect 22925 25109 22937 25112
rect 22971 25109 22983 25143
rect 27062 25140 27068 25152
rect 27023 25112 27068 25140
rect 22925 25103 22983 25109
rect 27062 25100 27068 25112
rect 27120 25100 27126 25152
rect 27448 25140 27476 25180
rect 30368 25171 30380 25217
rect 30432 25208 30438 25220
rect 30432 25180 30468 25208
rect 30374 25168 30380 25171
rect 30432 25168 30438 25180
rect 31386 25140 31392 25152
rect 27448 25112 31392 25140
rect 31386 25100 31392 25112
rect 31444 25140 31450 25152
rect 31481 25143 31539 25149
rect 31481 25140 31493 25143
rect 31444 25112 31493 25140
rect 31444 25100 31450 25112
rect 31481 25109 31493 25112
rect 31527 25109 31539 25143
rect 31481 25103 31539 25109
rect 1104 25050 35027 25072
rect 1104 24998 9390 25050
rect 9442 24998 9454 25050
rect 9506 24998 9518 25050
rect 9570 24998 9582 25050
rect 9634 24998 9646 25050
rect 9698 24998 17831 25050
rect 17883 24998 17895 25050
rect 17947 24998 17959 25050
rect 18011 24998 18023 25050
rect 18075 24998 18087 25050
rect 18139 24998 26272 25050
rect 26324 24998 26336 25050
rect 26388 24998 26400 25050
rect 26452 24998 26464 25050
rect 26516 24998 26528 25050
rect 26580 24998 34713 25050
rect 34765 24998 34777 25050
rect 34829 24998 34841 25050
rect 34893 24998 34905 25050
rect 34957 24998 34969 25050
rect 35021 24998 35027 25050
rect 1104 24976 35027 24998
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 15286 24936 15292 24948
rect 12308 24908 15292 24936
rect 12308 24896 12314 24908
rect 15286 24896 15292 24908
rect 15344 24896 15350 24948
rect 17034 24896 17040 24948
rect 17092 24936 17098 24948
rect 23566 24936 23572 24948
rect 17092 24908 23572 24936
rect 17092 24896 17098 24908
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 25130 24936 25136 24948
rect 23676 24908 25136 24936
rect 23676 24880 23704 24908
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 31478 24936 31484 24948
rect 31439 24908 31484 24936
rect 31478 24896 31484 24908
rect 31536 24896 31542 24948
rect 5074 24828 5080 24880
rect 5132 24868 5138 24880
rect 5261 24871 5319 24877
rect 5261 24868 5273 24871
rect 5132 24840 5273 24868
rect 5132 24828 5138 24840
rect 5261 24837 5273 24840
rect 5307 24837 5319 24871
rect 5261 24831 5319 24837
rect 15212 24840 15976 24868
rect 15212 24812 15240 24840
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 3878 24800 3884 24812
rect 2363 24772 3884 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 3878 24760 3884 24772
rect 3936 24760 3942 24812
rect 4154 24760 4160 24812
rect 4212 24800 4218 24812
rect 4212 24772 4646 24800
rect 4212 24760 4218 24772
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 6917 24803 6975 24809
rect 6917 24800 6929 24803
rect 6880 24772 6929 24800
rect 6880 24760 6886 24772
rect 6917 24769 6929 24772
rect 6963 24769 6975 24803
rect 7834 24800 7840 24812
rect 7590 24772 7840 24800
rect 6917 24763 6975 24769
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 14829 24803 14887 24809
rect 14829 24800 14841 24803
rect 12860 24772 14841 24800
rect 12860 24760 12866 24772
rect 14829 24769 14841 24772
rect 14875 24769 14887 24803
rect 14829 24763 14887 24769
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 2593 24735 2651 24741
rect 2593 24701 2605 24735
rect 2639 24732 2651 24735
rect 2774 24732 2780 24744
rect 2639 24704 2780 24732
rect 2639 24701 2651 24704
rect 2593 24695 2651 24701
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 4706 24732 4712 24744
rect 4667 24704 4712 24732
rect 4706 24692 4712 24704
rect 4764 24692 4770 24744
rect 7929 24735 7987 24741
rect 7929 24701 7941 24735
rect 7975 24732 7987 24735
rect 8478 24732 8484 24744
rect 7975 24704 8484 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 8478 24692 8484 24704
rect 8536 24692 8542 24744
rect 3881 24667 3939 24673
rect 3881 24633 3893 24667
rect 3927 24664 3939 24667
rect 4062 24664 4068 24676
rect 3927 24636 4068 24664
rect 3927 24633 3939 24636
rect 3881 24627 3939 24633
rect 4062 24624 4068 24636
rect 4120 24664 4126 24676
rect 4982 24664 4988 24676
rect 4120 24636 4988 24664
rect 4120 24624 4126 24636
rect 4982 24624 4988 24636
rect 5040 24624 5046 24676
rect 15120 24664 15148 24763
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15252 24772 15297 24800
rect 15252 24760 15258 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15948 24809 15976 24840
rect 20622 24828 20628 24880
rect 20680 24868 20686 24880
rect 21085 24871 21143 24877
rect 21085 24868 21097 24871
rect 20680 24840 21097 24868
rect 20680 24828 20686 24840
rect 21085 24837 21097 24840
rect 21131 24837 21143 24871
rect 21085 24831 21143 24837
rect 21453 24871 21511 24877
rect 21453 24837 21465 24871
rect 21499 24868 21511 24871
rect 22094 24868 22100 24880
rect 21499 24840 22100 24868
rect 21499 24837 21511 24840
rect 21453 24831 21511 24837
rect 22094 24828 22100 24840
rect 22152 24828 22158 24880
rect 23658 24868 23664 24880
rect 23571 24840 23664 24868
rect 23658 24828 23664 24840
rect 23716 24828 23722 24880
rect 27062 24868 27068 24880
rect 26160 24840 27068 24868
rect 15933 24803 15991 24809
rect 15436 24772 15481 24800
rect 15436 24760 15442 24772
rect 15933 24769 15945 24803
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 16298 24800 16304 24812
rect 16163 24772 16304 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24732 15347 24735
rect 16132 24732 16160 24763
rect 16298 24760 16304 24772
rect 16356 24760 16362 24812
rect 18141 24803 18199 24809
rect 18141 24769 18153 24803
rect 18187 24800 18199 24803
rect 18230 24800 18236 24812
rect 18187 24772 18236 24800
rect 18187 24769 18199 24772
rect 18141 24763 18199 24769
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 20990 24800 20996 24812
rect 20951 24772 20996 24800
rect 20990 24760 20996 24772
rect 21048 24760 21054 24812
rect 21269 24803 21327 24809
rect 21269 24800 21281 24803
rect 21100 24772 21281 24800
rect 15335 24704 16160 24732
rect 15335 24701 15347 24704
rect 15289 24695 15347 24701
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 17865 24735 17923 24741
rect 17865 24732 17877 24735
rect 17368 24704 17877 24732
rect 17368 24692 17374 24704
rect 17865 24701 17877 24704
rect 17911 24701 17923 24735
rect 19334 24732 19340 24744
rect 19295 24704 19340 24732
rect 17865 24695 17923 24701
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 15470 24664 15476 24676
rect 15120 24636 15476 24664
rect 15470 24624 15476 24636
rect 15528 24624 15534 24676
rect 21100 24664 21128 24772
rect 21269 24769 21281 24772
rect 21315 24800 21327 24803
rect 21542 24800 21548 24812
rect 21315 24772 21548 24800
rect 21315 24769 21327 24772
rect 21269 24763 21327 24769
rect 21542 24760 21548 24772
rect 21600 24800 21606 24812
rect 23750 24800 23756 24812
rect 21600 24772 23756 24800
rect 21600 24760 21606 24772
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 25222 24800 25228 24812
rect 25183 24772 25228 24800
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 25314 24760 25320 24812
rect 25372 24800 25378 24812
rect 26160 24809 26188 24840
rect 27062 24828 27068 24840
rect 27120 24828 27126 24880
rect 27154 24828 27160 24880
rect 27212 24868 27218 24880
rect 28629 24871 28687 24877
rect 28629 24868 28641 24871
rect 27212 24840 28641 24868
rect 27212 24828 27218 24840
rect 28629 24837 28641 24840
rect 28675 24837 28687 24871
rect 28629 24831 28687 24837
rect 28813 24871 28871 24877
rect 28813 24837 28825 24871
rect 28859 24837 28871 24871
rect 28813 24831 28871 24837
rect 26145 24803 26203 24809
rect 25372 24772 25417 24800
rect 25372 24760 25378 24772
rect 26145 24769 26157 24803
rect 26191 24769 26203 24803
rect 26145 24763 26203 24769
rect 28718 24760 28724 24812
rect 28776 24800 28782 24812
rect 28828 24800 28856 24831
rect 29086 24800 29092 24812
rect 28776 24772 28856 24800
rect 29047 24772 29092 24800
rect 28776 24760 28782 24772
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 30368 24803 30426 24809
rect 30368 24769 30380 24803
rect 30414 24800 30426 24803
rect 32306 24800 32312 24812
rect 30414 24772 32312 24800
rect 30414 24769 30426 24772
rect 30368 24763 30426 24769
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 22005 24735 22063 24741
rect 22005 24732 22017 24735
rect 21284 24704 22017 24732
rect 21284 24676 21312 24704
rect 22005 24701 22017 24704
rect 22051 24701 22063 24735
rect 22005 24695 22063 24701
rect 22186 24692 22192 24744
rect 22244 24732 22250 24744
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 22244 24704 22293 24732
rect 22244 24692 22250 24704
rect 22281 24701 22293 24704
rect 22327 24701 22339 24735
rect 22281 24695 22339 24701
rect 26421 24735 26479 24741
rect 26421 24701 26433 24735
rect 26467 24732 26479 24735
rect 28166 24732 28172 24744
rect 26467 24704 28172 24732
rect 26467 24701 26479 24704
rect 26421 24695 26479 24701
rect 28166 24692 28172 24704
rect 28224 24692 28230 24744
rect 30098 24732 30104 24744
rect 30059 24704 30104 24732
rect 30098 24692 30104 24704
rect 30156 24692 30162 24744
rect 18800 24636 21128 24664
rect 15010 24556 15016 24608
rect 15068 24596 15074 24608
rect 16117 24599 16175 24605
rect 16117 24596 16129 24599
rect 15068 24568 16129 24596
rect 15068 24556 15074 24568
rect 16117 24565 16129 24568
rect 16163 24565 16175 24599
rect 16117 24559 16175 24565
rect 18046 24556 18052 24608
rect 18104 24596 18110 24608
rect 18800 24596 18828 24636
rect 21266 24624 21272 24676
rect 21324 24624 21330 24676
rect 23308 24636 23520 24664
rect 18104 24568 18828 24596
rect 18104 24556 18110 24568
rect 20438 24556 20444 24608
rect 20496 24596 20502 24608
rect 23308 24596 23336 24636
rect 20496 24568 23336 24596
rect 23492 24596 23520 24636
rect 25038 24624 25044 24676
rect 25096 24664 25102 24676
rect 25133 24667 25191 24673
rect 25133 24664 25145 24667
rect 25096 24636 25145 24664
rect 25096 24624 25102 24636
rect 25133 24633 25145 24636
rect 25179 24633 25191 24667
rect 25133 24627 25191 24633
rect 25424 24636 28856 24664
rect 25424 24596 25452 24636
rect 25958 24596 25964 24608
rect 23492 24568 25452 24596
rect 25919 24568 25964 24596
rect 20496 24556 20502 24568
rect 25958 24556 25964 24568
rect 26016 24556 26022 24608
rect 26329 24599 26387 24605
rect 26329 24565 26341 24599
rect 26375 24596 26387 24599
rect 26602 24596 26608 24608
rect 26375 24568 26608 24596
rect 26375 24565 26387 24568
rect 26329 24559 26387 24565
rect 26602 24556 26608 24568
rect 26660 24556 26666 24608
rect 28828 24605 28856 24636
rect 28813 24599 28871 24605
rect 28813 24565 28825 24599
rect 28859 24565 28871 24599
rect 28813 24559 28871 24565
rect 1104 24506 34868 24528
rect 1104 24454 5170 24506
rect 5222 24454 5234 24506
rect 5286 24454 5298 24506
rect 5350 24454 5362 24506
rect 5414 24454 5426 24506
rect 5478 24454 13611 24506
rect 13663 24454 13675 24506
rect 13727 24454 13739 24506
rect 13791 24454 13803 24506
rect 13855 24454 13867 24506
rect 13919 24454 22052 24506
rect 22104 24454 22116 24506
rect 22168 24454 22180 24506
rect 22232 24454 22244 24506
rect 22296 24454 22308 24506
rect 22360 24454 30493 24506
rect 30545 24454 30557 24506
rect 30609 24454 30621 24506
rect 30673 24454 30685 24506
rect 30737 24454 30749 24506
rect 30801 24454 34868 24506
rect 1104 24432 34868 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 2832 24364 2877 24392
rect 2832 24352 2838 24364
rect 4338 24352 4344 24404
rect 4396 24392 4402 24404
rect 6822 24392 6828 24404
rect 4396 24364 6684 24392
rect 6783 24364 6828 24392
rect 4396 24352 4402 24364
rect 2317 24327 2375 24333
rect 2317 24293 2329 24327
rect 2363 24324 2375 24327
rect 2682 24324 2688 24336
rect 2363 24296 2688 24324
rect 2363 24293 2375 24296
rect 2317 24287 2375 24293
rect 2682 24284 2688 24296
rect 2740 24284 2746 24336
rect 2958 24284 2964 24336
rect 3016 24324 3022 24336
rect 5261 24327 5319 24333
rect 5261 24324 5273 24327
rect 3016 24296 5273 24324
rect 3016 24284 3022 24296
rect 5261 24293 5273 24296
rect 5307 24293 5319 24327
rect 6656 24324 6684 24364
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 16482 24352 16488 24404
rect 16540 24392 16546 24404
rect 16540 24364 18184 24392
rect 16540 24352 16546 24364
rect 6656 24296 7052 24324
rect 5261 24287 5319 24293
rect 2774 24256 2780 24268
rect 2056 24228 2780 24256
rect 2056 24197 2084 24228
rect 2774 24216 2780 24228
rect 2832 24216 2838 24268
rect 4157 24259 4215 24265
rect 4157 24256 4169 24259
rect 3068 24228 4169 24256
rect 2041 24191 2099 24197
rect 2041 24157 2053 24191
rect 2087 24157 2099 24191
rect 2958 24188 2964 24200
rect 2919 24160 2964 24188
rect 2041 24151 2099 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 3068 24197 3096 24228
rect 4157 24225 4169 24228
rect 4203 24225 4215 24259
rect 4157 24219 4215 24225
rect 4341 24259 4399 24265
rect 4341 24225 4353 24259
rect 4387 24256 4399 24259
rect 5074 24256 5080 24268
rect 4387 24228 5080 24256
rect 4387 24225 4399 24228
rect 4341 24219 4399 24225
rect 5074 24216 5080 24228
rect 5132 24256 5138 24268
rect 5169 24259 5227 24265
rect 5169 24256 5181 24259
rect 5132 24228 5181 24256
rect 5132 24216 5138 24228
rect 5169 24225 5181 24228
rect 5215 24225 5227 24259
rect 6914 24256 6920 24268
rect 5169 24219 5227 24225
rect 5368 24228 6920 24256
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 4433 24191 4491 24197
rect 4433 24157 4445 24191
rect 4479 24157 4491 24191
rect 4433 24151 4491 24157
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24157 4583 24191
rect 4525 24151 4583 24157
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24188 4675 24191
rect 5368 24188 5396 24228
rect 6914 24216 6920 24228
rect 6972 24216 6978 24268
rect 5534 24188 5540 24200
rect 4663 24160 5396 24188
rect 5495 24160 5540 24188
rect 4663 24157 4675 24160
rect 4617 24151 4675 24157
rect 2314 24120 2320 24132
rect 2275 24092 2320 24120
rect 2314 24080 2320 24092
rect 2372 24080 2378 24132
rect 2682 24080 2688 24132
rect 2740 24120 2746 24132
rect 3329 24123 3387 24129
rect 3329 24120 3341 24123
rect 2740 24092 3341 24120
rect 2740 24080 2746 24092
rect 3329 24089 3341 24092
rect 3375 24089 3387 24123
rect 3329 24083 3387 24089
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 3476 24092 3521 24120
rect 3476 24080 3482 24092
rect 2133 24055 2191 24061
rect 2133 24021 2145 24055
rect 2179 24052 2191 24055
rect 4338 24052 4344 24064
rect 2179 24024 4344 24052
rect 2179 24021 2191 24024
rect 2133 24015 2191 24021
rect 4338 24012 4344 24024
rect 4396 24012 4402 24064
rect 4448 24052 4476 24151
rect 4540 24120 4568 24151
rect 5534 24148 5540 24160
rect 5592 24148 5598 24200
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24157 5779 24191
rect 7024 24188 7052 24296
rect 15102 24284 15108 24336
rect 15160 24324 15166 24336
rect 18156 24324 18184 24364
rect 20990 24352 20996 24404
rect 21048 24392 21054 24404
rect 21048 24364 22508 24392
rect 21048 24352 21054 24364
rect 21008 24324 21036 24352
rect 15160 24296 15884 24324
rect 15160 24284 15166 24296
rect 13446 24216 13452 24268
rect 13504 24256 13510 24268
rect 13504 24228 14780 24256
rect 13504 24216 13510 24228
rect 7561 24191 7619 24197
rect 7561 24188 7573 24191
rect 7024 24160 7573 24188
rect 5721 24151 5779 24157
rect 7561 24157 7573 24160
rect 7607 24188 7619 24191
rect 8481 24191 8539 24197
rect 7607 24160 8248 24188
rect 7607 24157 7619 24160
rect 7561 24151 7619 24157
rect 5552 24120 5580 24148
rect 4540 24092 5580 24120
rect 5736 24120 5764 24151
rect 7742 24120 7748 24132
rect 5736 24092 7748 24120
rect 5736 24052 5764 24092
rect 7742 24080 7748 24092
rect 7800 24080 7806 24132
rect 8220 24120 8248 24160
rect 8481 24157 8493 24191
rect 8527 24188 8539 24191
rect 9306 24188 9312 24200
rect 8527 24160 9312 24188
rect 8527 24157 8539 24160
rect 8481 24151 8539 24157
rect 9306 24148 9312 24160
rect 9364 24148 9370 24200
rect 11882 24188 11888 24200
rect 11843 24160 11888 24188
rect 11882 24148 11888 24160
rect 11940 24148 11946 24200
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24188 12127 24191
rect 12434 24188 12440 24200
rect 12115 24160 12440 24188
rect 12115 24157 12127 24160
rect 12069 24151 12127 24157
rect 12434 24148 12440 24160
rect 12492 24188 12498 24200
rect 13262 24188 13268 24200
rect 12492 24160 13268 24188
rect 12492 24148 12498 24160
rect 13262 24148 13268 24160
rect 13320 24148 13326 24200
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 8570 24120 8576 24132
rect 8220 24092 8576 24120
rect 8570 24080 8576 24092
rect 8628 24080 8634 24132
rect 12250 24120 12256 24132
rect 8680 24092 12256 24120
rect 4448 24024 5764 24052
rect 5810 24012 5816 24064
rect 5868 24052 5874 24064
rect 8680 24052 8708 24092
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 14476 24120 14504 24151
rect 14550 24148 14556 24200
rect 14608 24188 14614 24200
rect 14752 24197 14780 24228
rect 15856 24200 15884 24296
rect 18156 24296 21036 24324
rect 14737 24191 14795 24197
rect 14608 24160 14653 24188
rect 14608 24148 14614 24160
rect 14737 24157 14749 24191
rect 14783 24157 14795 24191
rect 14737 24151 14795 24157
rect 14826 24148 14832 24200
rect 14884 24188 14890 24200
rect 15657 24191 15715 24197
rect 14884 24160 14929 24188
rect 14884 24148 14890 24160
rect 15657 24157 15669 24191
rect 15703 24157 15715 24191
rect 15657 24151 15715 24157
rect 15562 24120 15568 24132
rect 14476 24092 15568 24120
rect 15562 24080 15568 24092
rect 15620 24080 15626 24132
rect 15672 24120 15700 24151
rect 15838 24148 15844 24200
rect 15896 24188 15902 24200
rect 15896 24160 15989 24188
rect 15896 24148 15902 24160
rect 16390 24148 16396 24200
rect 16448 24188 16454 24200
rect 17954 24197 17960 24200
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 16448 24160 17049 24188
rect 16448 24148 16454 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24157 17279 24191
rect 17221 24151 17279 24157
rect 17911 24191 17960 24197
rect 17911 24157 17923 24191
rect 17957 24157 17960 24191
rect 17911 24151 17960 24157
rect 17236 24120 17264 24151
rect 17954 24148 17960 24151
rect 18012 24148 18018 24200
rect 18156 24197 18184 24296
rect 20898 24256 20904 24268
rect 20732 24228 20904 24256
rect 20732 24197 20760 24228
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 20993 24259 21051 24265
rect 20993 24225 21005 24259
rect 21039 24256 21051 24259
rect 21082 24256 21088 24268
rect 21039 24228 21088 24256
rect 21039 24225 21051 24228
rect 20993 24219 21051 24225
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 22480 24256 22508 24364
rect 25222 24352 25228 24404
rect 25280 24392 25286 24404
rect 27522 24392 27528 24404
rect 25280 24364 27528 24392
rect 25280 24352 25286 24364
rect 27522 24352 27528 24364
rect 27580 24352 27586 24404
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 30561 24395 30619 24401
rect 30561 24392 30573 24395
rect 30432 24364 30573 24392
rect 30432 24352 30438 24364
rect 30561 24361 30573 24364
rect 30607 24361 30619 24395
rect 30561 24355 30619 24361
rect 22833 24327 22891 24333
rect 22833 24293 22845 24327
rect 22879 24324 22891 24327
rect 23474 24324 23480 24336
rect 22879 24296 23480 24324
rect 22879 24293 22891 24296
rect 22833 24287 22891 24293
rect 23474 24284 23480 24296
rect 23532 24284 23538 24336
rect 23750 24284 23756 24336
rect 23808 24324 23814 24336
rect 28994 24324 29000 24336
rect 23808 24296 29000 24324
rect 23808 24284 23814 24296
rect 28994 24284 29000 24296
rect 29052 24284 29058 24336
rect 32398 24256 32404 24268
rect 22480 24228 23796 24256
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24157 20775 24191
rect 20717 24151 20775 24157
rect 20809 24191 20867 24197
rect 20809 24157 20821 24191
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 18049 24123 18107 24129
rect 18049 24120 18061 24123
rect 15672 24092 17172 24120
rect 17236 24092 18061 24120
rect 17144 24064 17172 24092
rect 18049 24089 18061 24092
rect 18095 24120 18107 24123
rect 18690 24120 18696 24132
rect 18095 24092 18696 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18690 24080 18696 24092
rect 18748 24080 18754 24132
rect 19702 24080 19708 24132
rect 19760 24120 19766 24132
rect 20824 24120 20852 24151
rect 21266 24148 21272 24200
rect 21324 24188 21330 24200
rect 23768 24197 23796 24228
rect 23860 24228 32404 24256
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21324 24160 21465 24188
rect 21324 24148 21330 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24157 23535 24191
rect 23477 24151 23535 24157
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24157 23811 24191
rect 23753 24151 23811 24157
rect 19760 24092 20852 24120
rect 21720 24123 21778 24129
rect 19760 24080 19766 24092
rect 21720 24089 21732 24123
rect 21766 24120 21778 24123
rect 23293 24123 23351 24129
rect 23293 24120 23305 24123
rect 21766 24092 23305 24120
rect 21766 24089 21778 24092
rect 21720 24083 21778 24089
rect 23293 24089 23305 24092
rect 23339 24089 23351 24123
rect 23492 24120 23520 24151
rect 23566 24120 23572 24132
rect 23479 24092 23572 24120
rect 23293 24083 23351 24089
rect 23566 24080 23572 24092
rect 23624 24120 23630 24132
rect 23860 24120 23888 24228
rect 32398 24216 32404 24228
rect 32456 24216 32462 24268
rect 25222 24188 25228 24200
rect 25183 24160 25228 24188
rect 25222 24148 25228 24160
rect 25280 24148 25286 24200
rect 25409 24191 25467 24197
rect 25409 24157 25421 24191
rect 25455 24188 25467 24191
rect 26694 24188 26700 24200
rect 25455 24160 26700 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24188 30803 24191
rect 30926 24188 30932 24200
rect 30791 24160 30932 24188
rect 30791 24157 30803 24160
rect 30745 24151 30803 24157
rect 30926 24148 30932 24160
rect 30984 24148 30990 24200
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24188 31079 24191
rect 32766 24188 32772 24200
rect 31067 24160 32772 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 23624 24092 23888 24120
rect 23624 24080 23630 24092
rect 25130 24080 25136 24132
rect 25188 24120 25194 24132
rect 31036 24120 31064 24151
rect 32766 24148 32772 24160
rect 32824 24148 32830 24200
rect 25188 24092 31064 24120
rect 25188 24080 25194 24092
rect 5868 24024 8708 24052
rect 12069 24055 12127 24061
rect 5868 24012 5874 24024
rect 12069 24021 12081 24055
rect 12115 24052 12127 24055
rect 12618 24052 12624 24064
rect 12115 24024 12624 24052
rect 12115 24021 12127 24024
rect 12069 24015 12127 24021
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 12894 24012 12900 24064
rect 12952 24052 12958 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 12952 24024 14289 24052
rect 12952 24012 12958 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 15470 24052 15476 24064
rect 15431 24024 15476 24052
rect 14277 24015 14335 24021
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 17126 24052 17132 24064
rect 17087 24024 17132 24052
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 17586 24012 17592 24064
rect 17644 24052 17650 24064
rect 17681 24055 17739 24061
rect 17681 24052 17693 24055
rect 17644 24024 17693 24052
rect 17644 24012 17650 24024
rect 17681 24021 17693 24024
rect 17727 24021 17739 24055
rect 17681 24015 17739 24021
rect 23661 24055 23719 24061
rect 23661 24021 23673 24055
rect 23707 24052 23719 24055
rect 24670 24052 24676 24064
rect 23707 24024 24676 24052
rect 23707 24021 23719 24024
rect 23661 24015 23719 24021
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 25314 24052 25320 24064
rect 25275 24024 25320 24052
rect 25314 24012 25320 24024
rect 25372 24012 25378 24064
rect 30929 24055 30987 24061
rect 30929 24021 30941 24055
rect 30975 24052 30987 24055
rect 31386 24052 31392 24064
rect 30975 24024 31392 24052
rect 30975 24021 30987 24024
rect 30929 24015 30987 24021
rect 31386 24012 31392 24024
rect 31444 24012 31450 24064
rect 1104 23962 35027 23984
rect 1104 23910 9390 23962
rect 9442 23910 9454 23962
rect 9506 23910 9518 23962
rect 9570 23910 9582 23962
rect 9634 23910 9646 23962
rect 9698 23910 17831 23962
rect 17883 23910 17895 23962
rect 17947 23910 17959 23962
rect 18011 23910 18023 23962
rect 18075 23910 18087 23962
rect 18139 23910 26272 23962
rect 26324 23910 26336 23962
rect 26388 23910 26400 23962
rect 26452 23910 26464 23962
rect 26516 23910 26528 23962
rect 26580 23910 34713 23962
rect 34765 23910 34777 23962
rect 34829 23910 34841 23962
rect 34893 23910 34905 23962
rect 34957 23910 34969 23962
rect 35021 23910 35027 23962
rect 1104 23888 35027 23910
rect 2314 23808 2320 23860
rect 2372 23848 2378 23860
rect 5077 23851 5135 23857
rect 5077 23848 5089 23851
rect 2372 23820 5089 23848
rect 2372 23808 2378 23820
rect 5077 23817 5089 23820
rect 5123 23817 5135 23851
rect 5077 23811 5135 23817
rect 7742 23808 7748 23860
rect 7800 23848 7806 23860
rect 14921 23851 14979 23857
rect 7800 23820 10272 23848
rect 7800 23808 7806 23820
rect 3326 23780 3332 23792
rect 2976 23752 3332 23780
rect 2976 23721 3004 23752
rect 3326 23740 3332 23752
rect 3384 23780 3390 23792
rect 5810 23780 5816 23792
rect 3384 23752 4660 23780
rect 3384 23740 3390 23752
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23681 3019 23715
rect 3694 23712 3700 23724
rect 3655 23684 3700 23712
rect 2961 23675 3019 23681
rect 3694 23672 3700 23684
rect 3752 23672 3758 23724
rect 4632 23712 4660 23752
rect 5000 23752 5816 23780
rect 5000 23712 5028 23752
rect 5810 23740 5816 23752
rect 5868 23740 5874 23792
rect 8478 23740 8484 23792
rect 8536 23780 8542 23792
rect 10244 23789 10272 23820
rect 14921 23817 14933 23851
rect 14967 23848 14979 23851
rect 15010 23848 15016 23860
rect 14967 23820 15016 23848
rect 14967 23817 14979 23820
rect 14921 23811 14979 23817
rect 15010 23808 15016 23820
rect 15068 23808 15074 23860
rect 15105 23851 15163 23857
rect 15105 23817 15117 23851
rect 15151 23848 15163 23851
rect 15378 23848 15384 23860
rect 15151 23820 15384 23848
rect 15151 23817 15163 23820
rect 15105 23811 15163 23817
rect 15378 23808 15384 23820
rect 15436 23848 15442 23860
rect 15933 23851 15991 23857
rect 15933 23848 15945 23851
rect 15436 23820 15945 23848
rect 15436 23808 15442 23820
rect 15933 23817 15945 23820
rect 15979 23817 15991 23851
rect 15933 23811 15991 23817
rect 16114 23808 16120 23860
rect 16172 23848 16178 23860
rect 19334 23848 19340 23860
rect 16172 23820 19340 23848
rect 16172 23808 16178 23820
rect 19334 23808 19340 23820
rect 19392 23848 19398 23860
rect 20622 23848 20628 23860
rect 19392 23820 20628 23848
rect 19392 23808 19398 23820
rect 20622 23808 20628 23820
rect 20680 23848 20686 23860
rect 30098 23848 30104 23860
rect 20680 23820 22324 23848
rect 30059 23820 30104 23848
rect 20680 23808 20686 23820
rect 10229 23783 10287 23789
rect 8536 23752 9904 23780
rect 8536 23740 8542 23752
rect 4632 23684 5028 23712
rect 4617 23647 4675 23653
rect 4617 23613 4629 23647
rect 4663 23644 4675 23647
rect 4706 23644 4712 23656
rect 4663 23616 4712 23644
rect 4663 23613 4675 23616
rect 4617 23607 4675 23613
rect 4706 23604 4712 23616
rect 4764 23604 4770 23656
rect 5000 23644 5028 23684
rect 5074 23672 5080 23724
rect 5132 23712 5138 23724
rect 5353 23715 5411 23721
rect 5353 23712 5365 23715
rect 5132 23684 5365 23712
rect 5132 23672 5138 23684
rect 5353 23681 5365 23684
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 5537 23715 5595 23721
rect 5537 23681 5549 23715
rect 5583 23712 5595 23715
rect 7190 23712 7196 23724
rect 5583 23684 7196 23712
rect 5583 23681 5595 23684
rect 5537 23675 5595 23681
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 9876 23721 9904 23752
rect 10229 23749 10241 23783
rect 10275 23749 10287 23783
rect 10229 23743 10287 23749
rect 19981 23783 20039 23789
rect 19981 23749 19993 23783
rect 20027 23780 20039 23783
rect 20714 23780 20720 23792
rect 20027 23752 20720 23780
rect 20027 23749 20039 23752
rect 19981 23743 20039 23749
rect 20714 23740 20720 23752
rect 20772 23780 20778 23792
rect 21910 23780 21916 23792
rect 20772 23752 21916 23780
rect 20772 23740 20778 23752
rect 21910 23740 21916 23752
rect 21968 23740 21974 23792
rect 22296 23789 22324 23820
rect 30098 23808 30104 23820
rect 30156 23808 30162 23860
rect 22281 23783 22339 23789
rect 22281 23749 22293 23783
rect 22327 23780 22339 23783
rect 25222 23780 25228 23792
rect 22327 23752 25228 23780
rect 22327 23749 22339 23752
rect 22281 23743 22339 23749
rect 25222 23740 25228 23752
rect 25280 23740 25286 23792
rect 28626 23780 28632 23792
rect 28587 23752 28632 23780
rect 28626 23740 28632 23752
rect 28684 23740 28690 23792
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 7760 23684 9229 23712
rect 5261 23647 5319 23653
rect 5261 23644 5273 23647
rect 5000 23616 5273 23644
rect 5261 23613 5273 23616
rect 5307 23613 5319 23647
rect 5261 23607 5319 23613
rect 5445 23647 5503 23653
rect 5445 23613 5457 23647
rect 5491 23644 5503 23647
rect 6730 23644 6736 23656
rect 5491 23616 6736 23644
rect 5491 23613 5503 23616
rect 5445 23607 5503 23613
rect 6730 23604 6736 23616
rect 6788 23604 6794 23656
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23613 6883 23647
rect 7098 23644 7104 23656
rect 7059 23616 7104 23644
rect 6825 23607 6883 23613
rect 6840 23576 6868 23607
rect 7098 23604 7104 23616
rect 7156 23604 7162 23656
rect 3896 23548 6868 23576
rect 3896 23520 3924 23548
rect 3878 23468 3884 23520
rect 3936 23468 3942 23520
rect 4246 23468 4252 23520
rect 4304 23508 4310 23520
rect 4614 23508 4620 23520
rect 4304 23480 4620 23508
rect 4304 23468 4310 23480
rect 4614 23468 4620 23480
rect 4672 23508 4678 23520
rect 7760 23508 7788 23684
rect 9217 23681 9229 23684
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23681 10103 23715
rect 12894 23712 12900 23724
rect 12855 23684 12900 23712
rect 10045 23675 10103 23681
rect 7926 23604 7932 23656
rect 7984 23644 7990 23656
rect 9033 23647 9091 23653
rect 9033 23644 9045 23647
rect 7984 23616 9045 23644
rect 7984 23604 7990 23616
rect 9033 23613 9045 23616
rect 9079 23613 9091 23647
rect 9033 23607 9091 23613
rect 9401 23647 9459 23653
rect 9401 23613 9413 23647
rect 9447 23644 9459 23647
rect 9490 23644 9496 23656
rect 9447 23616 9496 23644
rect 9447 23613 9459 23616
rect 9401 23607 9459 23613
rect 9490 23604 9496 23616
rect 9548 23604 9554 23656
rect 8294 23536 8300 23588
rect 8352 23576 8358 23588
rect 10060 23576 10088 23675
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 13262 23712 13268 23724
rect 13223 23684 13268 23712
rect 13262 23672 13268 23684
rect 13320 23672 13326 23724
rect 14369 23715 14427 23721
rect 14369 23681 14381 23715
rect 14415 23712 14427 23715
rect 15470 23712 15476 23724
rect 14415 23684 15476 23712
rect 14415 23681 14427 23684
rect 14369 23675 14427 23681
rect 15470 23672 15476 23684
rect 15528 23672 15534 23724
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 16117 23715 16175 23721
rect 16117 23712 16129 23715
rect 15896 23684 16129 23712
rect 15896 23672 15902 23684
rect 16117 23681 16129 23684
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23712 16359 23715
rect 17126 23712 17132 23724
rect 16347 23684 17132 23712
rect 16347 23681 16359 23684
rect 16301 23675 16359 23681
rect 17126 23672 17132 23684
rect 17184 23672 17190 23724
rect 20438 23712 20444 23724
rect 20399 23684 20444 23712
rect 20438 23672 20444 23684
rect 20496 23672 20502 23724
rect 20625 23715 20683 23721
rect 20625 23681 20637 23715
rect 20671 23712 20683 23715
rect 20898 23712 20904 23724
rect 20671 23684 20904 23712
rect 20671 23681 20683 23684
rect 20625 23675 20683 23681
rect 20898 23672 20904 23684
rect 20956 23712 20962 23724
rect 22649 23715 22707 23721
rect 20956 23684 22600 23712
rect 20956 23672 20962 23684
rect 12250 23644 12256 23656
rect 12211 23616 12256 23644
rect 12250 23604 12256 23616
rect 12308 23604 12314 23656
rect 12989 23647 13047 23653
rect 12989 23613 13001 23647
rect 13035 23613 13047 23647
rect 13170 23644 13176 23656
rect 13131 23616 13176 23644
rect 12989 23607 13047 23613
rect 8352 23548 10088 23576
rect 13004 23576 13032 23607
rect 13170 23604 13176 23616
rect 13228 23604 13234 23656
rect 14734 23604 14740 23656
rect 14792 23644 14798 23656
rect 14829 23647 14887 23653
rect 14829 23644 14841 23647
rect 14792 23616 14841 23644
rect 14792 23604 14798 23616
rect 14829 23613 14841 23616
rect 14875 23613 14887 23647
rect 15194 23644 15200 23656
rect 15107 23616 15200 23644
rect 14829 23607 14887 23613
rect 15194 23604 15200 23616
rect 15252 23604 15258 23656
rect 15286 23604 15292 23656
rect 15344 23644 15350 23656
rect 18414 23644 18420 23656
rect 15344 23616 18420 23644
rect 15344 23604 15350 23616
rect 18414 23604 18420 23616
rect 18472 23604 18478 23656
rect 20806 23644 20812 23656
rect 20767 23616 20812 23644
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 22572 23644 22600 23684
rect 22649 23681 22661 23715
rect 22695 23712 22707 23715
rect 23658 23712 23664 23724
rect 22695 23684 23664 23712
rect 22695 23681 22707 23684
rect 22649 23675 22707 23681
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 24670 23672 24676 23724
rect 24728 23712 24734 23724
rect 25501 23715 25559 23721
rect 25501 23712 25513 23715
rect 24728 23684 25513 23712
rect 24728 23672 24734 23684
rect 25501 23681 25513 23684
rect 25547 23681 25559 23715
rect 25501 23675 25559 23681
rect 27154 23644 27160 23656
rect 22572 23616 27160 23644
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 14182 23576 14188 23588
rect 13004 23548 14188 23576
rect 8352 23536 8358 23548
rect 14182 23536 14188 23548
rect 14240 23536 14246 23588
rect 14277 23579 14335 23585
rect 14277 23545 14289 23579
rect 14323 23576 14335 23579
rect 15203 23576 15231 23604
rect 14323 23548 15231 23576
rect 18693 23579 18751 23585
rect 14323 23545 14335 23548
rect 14277 23539 14335 23545
rect 18693 23545 18705 23579
rect 18739 23576 18751 23579
rect 19702 23576 19708 23588
rect 18739 23548 19708 23576
rect 18739 23545 18751 23548
rect 18693 23539 18751 23545
rect 19702 23536 19708 23548
rect 19760 23536 19766 23588
rect 4672 23480 7788 23508
rect 4672 23468 4678 23480
rect 8018 23468 8024 23520
rect 8076 23508 8082 23520
rect 8389 23511 8447 23517
rect 8389 23508 8401 23511
rect 8076 23480 8401 23508
rect 8076 23468 8082 23480
rect 8389 23477 8401 23480
rect 8435 23508 8447 23511
rect 9490 23508 9496 23520
rect 8435 23480 9496 23508
rect 8435 23477 8447 23480
rect 8389 23471 8447 23477
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 15470 23508 15476 23520
rect 15431 23480 15476 23508
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25409 23511 25467 23517
rect 25409 23508 25421 23511
rect 25004 23480 25421 23508
rect 25004 23468 25010 23480
rect 25409 23477 25421 23480
rect 25455 23477 25467 23511
rect 25409 23471 25467 23477
rect 1104 23418 34868 23440
rect 1104 23366 5170 23418
rect 5222 23366 5234 23418
rect 5286 23366 5298 23418
rect 5350 23366 5362 23418
rect 5414 23366 5426 23418
rect 5478 23366 13611 23418
rect 13663 23366 13675 23418
rect 13727 23366 13739 23418
rect 13791 23366 13803 23418
rect 13855 23366 13867 23418
rect 13919 23366 22052 23418
rect 22104 23366 22116 23418
rect 22168 23366 22180 23418
rect 22232 23366 22244 23418
rect 22296 23366 22308 23418
rect 22360 23366 30493 23418
rect 30545 23366 30557 23418
rect 30609 23366 30621 23418
rect 30673 23366 30685 23418
rect 30737 23366 30749 23418
rect 30801 23366 34868 23418
rect 1104 23344 34868 23366
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3237 23307 3295 23313
rect 3237 23304 3249 23307
rect 2924 23276 3249 23304
rect 2924 23264 2930 23276
rect 3237 23273 3249 23276
rect 3283 23273 3295 23307
rect 3237 23267 3295 23273
rect 3329 23307 3387 23313
rect 3329 23273 3341 23307
rect 3375 23304 3387 23307
rect 3418 23304 3424 23316
rect 3375 23276 3424 23304
rect 3375 23273 3387 23276
rect 3329 23267 3387 23273
rect 3418 23264 3424 23276
rect 3476 23264 3482 23316
rect 4157 23307 4215 23313
rect 4157 23273 4169 23307
rect 4203 23304 4215 23307
rect 4246 23304 4252 23316
rect 4203 23276 4252 23304
rect 4203 23273 4215 23276
rect 4157 23267 4215 23273
rect 4246 23264 4252 23276
rect 4304 23264 4310 23316
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7098 23304 7104 23316
rect 6963 23276 7104 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7098 23264 7104 23276
rect 7156 23264 7162 23316
rect 10226 23304 10232 23316
rect 7300 23276 10232 23304
rect 7300 23236 7328 23276
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 18690 23304 18696 23316
rect 10336 23276 12434 23304
rect 18651 23276 18696 23304
rect 3160 23208 7328 23236
rect 3160 23109 3188 23208
rect 7374 23196 7380 23248
rect 7432 23236 7438 23248
rect 9125 23239 9183 23245
rect 9125 23236 9137 23239
rect 7432 23208 9137 23236
rect 7432 23196 7438 23208
rect 9125 23205 9137 23208
rect 9171 23205 9183 23239
rect 9125 23199 9183 23205
rect 9858 23196 9864 23248
rect 9916 23236 9922 23248
rect 10336 23236 10364 23276
rect 9916 23208 10364 23236
rect 9916 23196 9922 23208
rect 3421 23171 3479 23177
rect 3421 23137 3433 23171
rect 3467 23168 3479 23171
rect 4154 23168 4160 23180
rect 3467 23140 4160 23168
rect 3467 23137 3479 23140
rect 3421 23131 3479 23137
rect 4154 23128 4160 23140
rect 4212 23128 4218 23180
rect 7208 23140 7696 23168
rect 3145 23103 3203 23109
rect 3145 23069 3157 23103
rect 3191 23069 3203 23103
rect 7098 23100 7104 23112
rect 7059 23072 7104 23100
rect 3145 23063 3203 23069
rect 7098 23060 7104 23072
rect 7156 23060 7162 23112
rect 7208 23044 7236 23140
rect 7374 23060 7380 23112
rect 7432 23109 7438 23112
rect 7432 23103 7461 23109
rect 7449 23069 7461 23103
rect 7558 23100 7564 23112
rect 7519 23072 7564 23100
rect 7432 23063 7461 23069
rect 7432 23060 7438 23063
rect 7558 23060 7564 23072
rect 7616 23060 7622 23112
rect 7668 23100 7696 23140
rect 8018 23128 8024 23180
rect 8076 23168 8082 23180
rect 8297 23171 8355 23177
rect 8297 23168 8309 23171
rect 8076 23140 8309 23168
rect 8076 23128 8082 23140
rect 8297 23137 8309 23140
rect 8343 23137 8355 23171
rect 8297 23131 8355 23137
rect 8573 23171 8631 23177
rect 8573 23137 8585 23171
rect 8619 23137 8631 23171
rect 8573 23131 8631 23137
rect 8113 23103 8171 23109
rect 8113 23100 8125 23103
rect 7668 23072 8125 23100
rect 8113 23069 8125 23072
rect 8159 23069 8171 23103
rect 8113 23063 8171 23069
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23069 8263 23103
rect 8205 23063 8263 23069
rect 4341 23035 4399 23041
rect 4341 23001 4353 23035
rect 4387 23032 4399 23035
rect 5074 23032 5080 23044
rect 4387 23004 5080 23032
rect 4387 23001 4399 23004
rect 4341 22995 4399 23001
rect 5074 22992 5080 23004
rect 5132 22992 5138 23044
rect 7190 23032 7196 23044
rect 7151 23004 7196 23032
rect 7190 22992 7196 23004
rect 7248 22992 7254 23044
rect 7285 23035 7343 23041
rect 7285 23001 7297 23035
rect 7331 23032 7343 23035
rect 7742 23032 7748 23044
rect 7331 23004 7748 23032
rect 7331 23001 7343 23004
rect 7285 22995 7343 23001
rect 7742 22992 7748 23004
rect 7800 22992 7806 23044
rect 3970 22964 3976 22976
rect 3931 22936 3976 22964
rect 3970 22924 3976 22936
rect 4028 22924 4034 22976
rect 4141 22967 4199 22973
rect 4141 22933 4153 22967
rect 4187 22964 4199 22967
rect 4706 22964 4712 22976
rect 4187 22936 4712 22964
rect 4187 22933 4199 22936
rect 4141 22927 4199 22933
rect 4706 22924 4712 22936
rect 4764 22924 4770 22976
rect 6730 22924 6736 22976
rect 6788 22964 6794 22976
rect 8220 22964 8248 23063
rect 8386 23060 8392 23112
rect 8444 23100 8450 23112
rect 8444 23072 8489 23100
rect 8444 23060 8450 23072
rect 8588 23032 8616 23131
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 10042 23168 10048 23180
rect 9548 23140 10048 23168
rect 9548 23128 9554 23140
rect 10042 23128 10048 23140
rect 10100 23168 10106 23180
rect 10100 23140 12296 23168
rect 10100 23128 10106 23140
rect 8662 23060 8668 23112
rect 8720 23100 8726 23112
rect 9309 23103 9367 23109
rect 8720 23094 9260 23100
rect 9309 23094 9321 23103
rect 8720 23072 9321 23094
rect 8720 23060 8726 23072
rect 9232 23069 9321 23072
rect 9355 23069 9367 23103
rect 9232 23066 9367 23069
rect 9309 23063 9367 23066
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 9456 23072 9501 23100
rect 9456 23060 9462 23072
rect 12066 23060 12072 23112
rect 12124 23100 12130 23112
rect 12124 23072 12169 23100
rect 12124 23060 12130 23072
rect 9125 23035 9183 23041
rect 9125 23032 9137 23035
rect 8588 23004 9137 23032
rect 9125 23001 9137 23004
rect 9171 23001 9183 23035
rect 9125 22995 9183 23001
rect 9766 22992 9772 23044
rect 9824 23032 9830 23044
rect 11793 23035 11851 23041
rect 9824 23004 10626 23032
rect 9824 22992 9830 23004
rect 11793 23001 11805 23035
rect 11839 23032 11851 23035
rect 11882 23032 11888 23044
rect 11839 23004 11888 23032
rect 11839 23001 11851 23004
rect 11793 22995 11851 23001
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 12268 23032 12296 23140
rect 12406 23100 12434 23276
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 21910 23304 21916 23316
rect 21871 23276 21916 23304
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 31846 23264 31852 23316
rect 31904 23304 31910 23316
rect 33134 23304 33140 23316
rect 31904 23276 33140 23304
rect 31904 23264 31910 23276
rect 33134 23264 33140 23276
rect 33192 23264 33198 23316
rect 15378 23236 15384 23248
rect 15304 23208 15384 23236
rect 15194 23168 15200 23180
rect 15155 23140 15200 23168
rect 15194 23128 15200 23140
rect 15252 23128 15258 23180
rect 15304 23177 15332 23208
rect 15378 23196 15384 23208
rect 15436 23196 15442 23248
rect 15565 23239 15623 23245
rect 15565 23205 15577 23239
rect 15611 23236 15623 23239
rect 16117 23239 16175 23245
rect 16117 23236 16129 23239
rect 15611 23208 16129 23236
rect 15611 23205 15623 23208
rect 15565 23199 15623 23205
rect 16117 23205 16129 23208
rect 16163 23205 16175 23239
rect 16117 23199 16175 23205
rect 19610 23196 19616 23248
rect 19668 23236 19674 23248
rect 19705 23239 19763 23245
rect 19705 23236 19717 23239
rect 19668 23208 19717 23236
rect 19668 23196 19674 23208
rect 19705 23205 19717 23208
rect 19751 23205 19763 23239
rect 19705 23199 19763 23205
rect 19978 23196 19984 23248
rect 20036 23236 20042 23248
rect 28718 23236 28724 23248
rect 20036 23208 28724 23236
rect 20036 23196 20042 23208
rect 28718 23196 28724 23208
rect 28776 23196 28782 23248
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 15528 23140 16497 23168
rect 15528 23128 15534 23140
rect 16485 23137 16497 23140
rect 16531 23137 16543 23171
rect 17310 23168 17316 23180
rect 17271 23140 17316 23168
rect 16485 23131 16543 23137
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 24946 23168 24952 23180
rect 24907 23140 24952 23168
rect 24946 23128 24952 23140
rect 25004 23128 25010 23180
rect 25314 23168 25320 23180
rect 25275 23140 25320 23168
rect 25314 23128 25320 23140
rect 25372 23128 25378 23180
rect 31018 23128 31024 23180
rect 31076 23168 31082 23180
rect 32674 23168 32680 23180
rect 31076 23140 32076 23168
rect 32635 23140 32680 23168
rect 31076 23128 31082 23140
rect 32048 23112 32076 23140
rect 32674 23128 32680 23140
rect 32732 23128 32738 23180
rect 33134 23168 33140 23180
rect 33047 23140 33140 23168
rect 33134 23128 33140 23140
rect 33192 23168 33198 23180
rect 33192 23140 33824 23168
rect 33192 23128 33198 23140
rect 12529 23103 12587 23109
rect 12529 23100 12541 23103
rect 12406 23072 12541 23100
rect 12529 23069 12541 23072
rect 12575 23069 12587 23103
rect 13998 23100 14004 23112
rect 12529 23063 12587 23069
rect 13188 23072 14004 23100
rect 13188 23032 13216 23072
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 17586 23109 17592 23112
rect 15105 23103 15163 23109
rect 15105 23100 15117 23103
rect 15068 23072 15117 23100
rect 15068 23060 15074 23072
rect 15105 23069 15117 23072
rect 15151 23069 15163 23103
rect 15105 23063 15163 23069
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23069 15439 23103
rect 17580 23100 17592 23109
rect 17547 23072 17592 23100
rect 15381 23063 15439 23069
rect 17580 23063 17592 23072
rect 12268 23004 13216 23032
rect 13265 23035 13323 23041
rect 13265 23001 13277 23035
rect 13311 23001 13323 23035
rect 13265 22995 13323 23001
rect 10318 22964 10324 22976
rect 6788 22936 10324 22964
rect 6788 22924 6794 22936
rect 10318 22924 10324 22936
rect 10376 22924 10382 22976
rect 10410 22924 10416 22976
rect 10468 22964 10474 22976
rect 13280 22964 13308 22995
rect 14734 22992 14740 23044
rect 14792 23032 14798 23044
rect 15396 23032 15424 23063
rect 17586 23060 17592 23063
rect 17644 23060 17650 23112
rect 19426 23100 19432 23112
rect 19387 23072 19432 23100
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 19702 23100 19708 23112
rect 19663 23072 19708 23100
rect 19702 23060 19708 23072
rect 19760 23060 19766 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 20806 23100 20812 23112
rect 20671 23072 20812 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 22738 23060 22744 23112
rect 22796 23100 22802 23112
rect 24857 23103 24915 23109
rect 24857 23100 24869 23103
rect 22796 23072 24869 23100
rect 22796 23060 22802 23072
rect 24857 23069 24869 23072
rect 24903 23069 24915 23103
rect 27522 23100 27528 23112
rect 27483 23072 27528 23100
rect 24857 23063 24915 23069
rect 27522 23060 27528 23072
rect 27580 23060 27586 23112
rect 27982 23100 27988 23112
rect 27943 23072 27988 23100
rect 27982 23060 27988 23072
rect 28040 23060 28046 23112
rect 28258 23100 28264 23112
rect 28219 23072 28264 23100
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 31754 23100 31760 23112
rect 31715 23072 31760 23100
rect 31754 23060 31760 23072
rect 31812 23060 31818 23112
rect 32030 23100 32036 23112
rect 31991 23072 32036 23100
rect 32030 23060 32036 23072
rect 32088 23060 32094 23112
rect 32398 23060 32404 23112
rect 32456 23100 32462 23112
rect 32769 23103 32827 23109
rect 32769 23100 32781 23103
rect 32456 23072 32781 23100
rect 32456 23060 32462 23072
rect 32769 23069 32781 23072
rect 32815 23069 32827 23103
rect 32769 23063 32827 23069
rect 33318 23060 33324 23112
rect 33376 23100 33382 23112
rect 33796 23109 33824 23140
rect 33597 23103 33655 23109
rect 33597 23100 33609 23103
rect 33376 23072 33609 23100
rect 33376 23060 33382 23072
rect 33597 23069 33609 23072
rect 33643 23069 33655 23103
rect 33597 23063 33655 23069
rect 33781 23103 33839 23109
rect 33781 23069 33793 23103
rect 33827 23069 33839 23103
rect 33781 23063 33839 23069
rect 14792 23004 15424 23032
rect 14792 22992 14798 23004
rect 27614 22992 27620 23044
rect 27672 23032 27678 23044
rect 27801 23035 27859 23041
rect 27801 23032 27813 23035
rect 27672 23004 27813 23032
rect 27672 22992 27678 23004
rect 27801 23001 27813 23004
rect 27847 23032 27859 23035
rect 28534 23032 28540 23044
rect 27847 23004 28540 23032
rect 27847 23001 27859 23004
rect 27801 22995 27859 23001
rect 28534 22992 28540 23004
rect 28592 22992 28598 23044
rect 10468 22936 13308 22964
rect 10468 22924 10474 22936
rect 14642 22924 14648 22976
rect 14700 22964 14706 22976
rect 16025 22967 16083 22973
rect 16025 22964 16037 22967
rect 14700 22936 16037 22964
rect 14700 22924 14706 22936
rect 16025 22933 16037 22936
rect 16071 22933 16083 22967
rect 16025 22927 16083 22933
rect 24673 22967 24731 22973
rect 24673 22933 24685 22967
rect 24719 22964 24731 22967
rect 24854 22964 24860 22976
rect 24719 22936 24860 22964
rect 24719 22933 24731 22936
rect 24673 22927 24731 22933
rect 24854 22924 24860 22936
rect 24912 22924 24918 22976
rect 24946 22924 24952 22976
rect 25004 22964 25010 22976
rect 25041 22967 25099 22973
rect 25041 22964 25053 22967
rect 25004 22936 25053 22964
rect 25004 22924 25010 22936
rect 25041 22933 25053 22936
rect 25087 22933 25099 22967
rect 25222 22964 25228 22976
rect 25183 22936 25228 22964
rect 25041 22927 25099 22933
rect 25222 22924 25228 22936
rect 25280 22924 25286 22976
rect 29730 22924 29736 22976
rect 29788 22964 29794 22976
rect 31021 22967 31079 22973
rect 31021 22964 31033 22967
rect 29788 22936 31033 22964
rect 29788 22924 29794 22936
rect 31021 22933 31033 22936
rect 31067 22933 31079 22967
rect 31021 22927 31079 22933
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 33689 22967 33747 22973
rect 33689 22964 33701 22967
rect 33560 22936 33701 22964
rect 33560 22924 33566 22936
rect 33689 22933 33701 22936
rect 33735 22933 33747 22967
rect 33689 22927 33747 22933
rect 1104 22874 35027 22896
rect 1104 22822 9390 22874
rect 9442 22822 9454 22874
rect 9506 22822 9518 22874
rect 9570 22822 9582 22874
rect 9634 22822 9646 22874
rect 9698 22822 17831 22874
rect 17883 22822 17895 22874
rect 17947 22822 17959 22874
rect 18011 22822 18023 22874
rect 18075 22822 18087 22874
rect 18139 22822 26272 22874
rect 26324 22822 26336 22874
rect 26388 22822 26400 22874
rect 26452 22822 26464 22874
rect 26516 22822 26528 22874
rect 26580 22822 34713 22874
rect 34765 22822 34777 22874
rect 34829 22822 34841 22874
rect 34893 22822 34905 22874
rect 34957 22822 34969 22874
rect 35021 22822 35027 22874
rect 1104 22800 35027 22822
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 7558 22760 7564 22772
rect 7239 22732 7564 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 7558 22720 7564 22732
rect 7616 22720 7622 22772
rect 9306 22720 9312 22772
rect 9364 22760 9370 22772
rect 9364 22732 10272 22760
rect 9364 22720 9370 22732
rect 7098 22652 7104 22704
rect 7156 22692 7162 22704
rect 8113 22695 8171 22701
rect 8113 22692 8125 22695
rect 7156 22664 8125 22692
rect 7156 22652 7162 22664
rect 8113 22661 8125 22664
rect 8159 22661 8171 22695
rect 8294 22692 8300 22704
rect 8255 22664 8300 22692
rect 8113 22655 8171 22661
rect 8294 22652 8300 22664
rect 8352 22652 8358 22704
rect 8478 22692 8484 22704
rect 8439 22664 8484 22692
rect 8478 22652 8484 22664
rect 8536 22652 8542 22704
rect 9677 22695 9735 22701
rect 9677 22661 9689 22695
rect 9723 22692 9735 22695
rect 9766 22692 9772 22704
rect 9723 22664 9772 22692
rect 9723 22661 9735 22664
rect 9677 22655 9735 22661
rect 9766 22652 9772 22664
rect 9824 22652 9830 22704
rect 10244 22692 10272 22732
rect 10318 22720 10324 22772
rect 10376 22760 10382 22772
rect 10778 22760 10784 22772
rect 10376 22732 10784 22760
rect 10376 22720 10382 22732
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 31846 22760 31852 22772
rect 12406 22732 12572 22760
rect 12406 22692 12434 22732
rect 12544 22701 12572 22732
rect 14476 22732 31852 22760
rect 10244 22664 12434 22692
rect 12529 22695 12587 22701
rect 12529 22661 12541 22695
rect 12575 22661 12587 22695
rect 14369 22695 14427 22701
rect 14369 22692 14381 22695
rect 12529 22655 12587 22661
rect 13280 22664 14381 22692
rect 4338 22584 4344 22636
rect 4396 22624 4402 22636
rect 4433 22627 4491 22633
rect 4433 22624 4445 22627
rect 4396 22596 4445 22624
rect 4396 22584 4402 22596
rect 4433 22593 4445 22596
rect 4479 22593 4491 22627
rect 4433 22587 4491 22593
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7466 22624 7472 22636
rect 7423 22596 7472 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 9401 22627 9459 22633
rect 9401 22593 9413 22627
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 9585 22627 9643 22633
rect 9585 22593 9597 22627
rect 9631 22593 9643 22627
rect 9585 22587 9643 22593
rect 10321 22627 10379 22633
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 10410 22624 10416 22636
rect 10367 22596 10416 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 3694 22516 3700 22568
rect 3752 22556 3758 22568
rect 4985 22559 5043 22565
rect 4985 22556 4997 22559
rect 3752 22528 4997 22556
rect 3752 22516 3758 22528
rect 4985 22525 4997 22528
rect 5031 22556 5043 22559
rect 7576 22556 7604 22587
rect 5031 22528 7604 22556
rect 7668 22556 7696 22587
rect 8386 22556 8392 22568
rect 7668 22528 8392 22556
rect 5031 22525 5043 22528
rect 4985 22519 5043 22525
rect 8386 22516 8392 22528
rect 8444 22516 8450 22568
rect 8662 22448 8668 22500
rect 8720 22488 8726 22500
rect 9416 22488 9444 22587
rect 9600 22556 9628 22587
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 11698 22624 11704 22636
rect 11659 22596 11704 22624
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 12434 22624 12440 22636
rect 11931 22596 12440 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12618 22584 12624 22636
rect 12676 22624 12682 22636
rect 13280 22633 13308 22664
rect 14369 22661 14381 22664
rect 14415 22661 14427 22695
rect 14369 22655 14427 22661
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12676 22596 12909 22624
rect 12676 22584 12682 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13265 22627 13323 22633
rect 13265 22593 13277 22627
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 10965 22559 11023 22565
rect 10965 22556 10977 22559
rect 9600 22528 10977 22556
rect 10965 22525 10977 22528
rect 11011 22556 11023 22559
rect 11790 22556 11796 22568
rect 11011 22528 11796 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 11974 22488 11980 22500
rect 8720 22460 9352 22488
rect 9416 22460 11980 22488
rect 8720 22448 8726 22460
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 9214 22420 9220 22432
rect 5132 22392 9220 22420
rect 5132 22380 5138 22392
rect 9214 22380 9220 22392
rect 9272 22380 9278 22432
rect 9324 22420 9352 22460
rect 11974 22448 11980 22460
rect 12032 22448 12038 22500
rect 12894 22448 12900 22500
rect 12952 22488 12958 22500
rect 13372 22488 13400 22587
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 13633 22627 13691 22633
rect 13633 22624 13645 22627
rect 13504 22596 13645 22624
rect 13504 22584 13510 22596
rect 13633 22593 13645 22596
rect 13679 22593 13691 22627
rect 13633 22587 13691 22593
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22624 13967 22627
rect 14476 22624 14504 22732
rect 31846 22720 31852 22732
rect 31904 22720 31910 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32401 22763 32459 22769
rect 32401 22760 32413 22763
rect 32088 22732 32413 22760
rect 32088 22720 32094 22732
rect 32401 22729 32413 22732
rect 32447 22729 32459 22763
rect 32401 22723 32459 22729
rect 14734 22652 14740 22704
rect 14792 22692 14798 22704
rect 23753 22695 23811 22701
rect 14792 22664 17540 22692
rect 14792 22652 14798 22664
rect 14642 22624 14648 22636
rect 13955 22596 14504 22624
rect 14603 22596 14648 22624
rect 13955 22593 13967 22596
rect 13909 22587 13967 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22593 15347 22627
rect 15470 22624 15476 22636
rect 15431 22596 15476 22624
rect 15289 22587 15347 22593
rect 14182 22516 14188 22568
rect 14240 22556 14246 22568
rect 14369 22559 14427 22565
rect 14369 22556 14381 22559
rect 14240 22528 14381 22556
rect 14240 22516 14246 22528
rect 14369 22525 14381 22528
rect 14415 22525 14427 22559
rect 15304 22556 15332 22587
rect 15470 22584 15476 22596
rect 15528 22584 15534 22636
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 16390 22624 16396 22636
rect 15620 22596 16396 22624
rect 15620 22584 15626 22596
rect 16390 22584 16396 22596
rect 16448 22584 16454 22636
rect 17126 22584 17132 22636
rect 17184 22624 17190 22636
rect 17512 22633 17540 22664
rect 18156 22664 20208 22692
rect 18156 22633 18184 22664
rect 17313 22627 17371 22633
rect 17313 22624 17325 22627
rect 17184 22596 17325 22624
rect 17184 22584 17190 22596
rect 17313 22593 17325 22596
rect 17359 22593 17371 22627
rect 17313 22587 17371 22593
rect 17497 22627 17555 22633
rect 17497 22593 17509 22627
rect 17543 22624 17555 22627
rect 18141 22627 18199 22633
rect 18141 22624 18153 22627
rect 17543 22596 18153 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 18141 22593 18153 22596
rect 18187 22593 18199 22627
rect 18141 22587 18199 22593
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22624 18659 22627
rect 18690 22624 18696 22636
rect 18647 22596 18696 22624
rect 18647 22593 18659 22596
rect 18601 22587 18659 22593
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 19978 22584 19984 22636
rect 20036 22624 20042 22636
rect 20180 22633 20208 22664
rect 22020 22664 23704 22692
rect 20146 22627 20208 22633
rect 20036 22596 20081 22624
rect 20036 22584 20042 22596
rect 20146 22593 20158 22627
rect 20192 22596 20208 22627
rect 20257 22627 20315 22633
rect 20192 22593 20204 22596
rect 20146 22587 20204 22593
rect 20257 22593 20269 22627
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22624 20407 22627
rect 20530 22624 20536 22636
rect 20395 22596 20536 22624
rect 20395 22593 20407 22596
rect 20349 22587 20407 22593
rect 18233 22559 18291 22565
rect 15304 22528 18184 22556
rect 14369 22519 14427 22525
rect 12952 22460 13400 22488
rect 17405 22491 17463 22497
rect 12952 22448 12958 22460
rect 17405 22457 17417 22491
rect 17451 22488 17463 22491
rect 18046 22488 18052 22500
rect 17451 22460 18052 22488
rect 17451 22457 17463 22460
rect 17405 22451 17463 22457
rect 18046 22448 18052 22460
rect 18104 22448 18110 22500
rect 18156 22488 18184 22528
rect 18233 22525 18245 22559
rect 18279 22556 18291 22559
rect 19334 22556 19340 22568
rect 18279 22528 19340 22556
rect 18279 22525 18291 22528
rect 18233 22519 18291 22525
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 20272 22488 20300 22587
rect 20530 22584 20536 22596
rect 20588 22584 20594 22636
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 21818 22624 21824 22636
rect 21048 22596 21824 22624
rect 21048 22584 21054 22596
rect 21818 22584 21824 22596
rect 21876 22624 21882 22636
rect 22020 22633 22048 22664
rect 23676 22633 23704 22664
rect 23753 22661 23765 22695
rect 23799 22692 23811 22695
rect 25222 22692 25228 22704
rect 23799 22664 25228 22692
rect 23799 22661 23811 22664
rect 23753 22655 23811 22661
rect 25222 22652 25228 22664
rect 25280 22652 25286 22704
rect 28258 22652 28264 22704
rect 28316 22692 28322 22704
rect 33045 22695 33103 22701
rect 28316 22664 30052 22692
rect 28316 22652 28322 22664
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21876 22596 22017 22624
rect 21876 22584 21882 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22189 22627 22247 22633
rect 22189 22593 22201 22627
rect 22235 22593 22247 22627
rect 22189 22587 22247 22593
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22624 24915 22627
rect 27154 22624 27160 22636
rect 24903 22596 27160 22624
rect 24903 22593 24915 22596
rect 24857 22587 24915 22593
rect 22005 22491 22063 22497
rect 22005 22488 22017 22491
rect 18156 22460 19932 22488
rect 20272 22460 22017 22488
rect 10318 22420 10324 22432
rect 9324 22392 10324 22420
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 11793 22423 11851 22429
rect 11793 22389 11805 22423
rect 11839 22420 11851 22423
rect 12986 22420 12992 22432
rect 11839 22392 12992 22420
rect 11839 22389 11851 22392
rect 11793 22383 11851 22389
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 14553 22423 14611 22429
rect 14553 22389 14565 22423
rect 14599 22420 14611 22423
rect 15105 22423 15163 22429
rect 15105 22420 15117 22423
rect 14599 22392 15117 22420
rect 14599 22389 14611 22392
rect 14553 22383 14611 22389
rect 15105 22389 15117 22392
rect 15151 22389 15163 22423
rect 17954 22420 17960 22432
rect 17915 22392 17960 22420
rect 15105 22383 15163 22389
rect 17954 22380 17960 22392
rect 18012 22380 18018 22432
rect 19794 22420 19800 22432
rect 19755 22392 19800 22420
rect 19794 22380 19800 22392
rect 19852 22380 19858 22432
rect 19904 22420 19932 22460
rect 22005 22457 22017 22460
rect 22051 22457 22063 22491
rect 22204 22488 22232 22587
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 27982 22624 27988 22636
rect 27943 22596 27988 22624
rect 27982 22584 27988 22596
rect 28040 22584 28046 22636
rect 28368 22633 28396 22664
rect 28353 22627 28411 22633
rect 28353 22593 28365 22627
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 28534 22584 28540 22636
rect 28592 22624 28598 22636
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 28592 22596 29929 22624
rect 28592 22584 28598 22596
rect 29917 22593 29929 22596
rect 29963 22593 29975 22627
rect 29917 22587 29975 22593
rect 24762 22556 24768 22568
rect 24723 22528 24768 22556
rect 24762 22516 24768 22528
rect 24820 22516 24826 22568
rect 25133 22559 25191 22565
rect 25133 22525 25145 22559
rect 25179 22556 25191 22559
rect 26142 22556 26148 22568
rect 25179 22528 26148 22556
rect 25179 22525 25191 22528
rect 25133 22519 25191 22525
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 26970 22516 26976 22568
rect 27028 22516 27034 22568
rect 29730 22556 29736 22568
rect 29643 22528 29736 22556
rect 29730 22516 29736 22528
rect 29788 22516 29794 22568
rect 30024 22556 30052 22664
rect 33045 22661 33057 22695
rect 33091 22692 33103 22695
rect 33134 22692 33140 22704
rect 33091 22664 33140 22692
rect 33091 22661 33103 22664
rect 33045 22655 33103 22661
rect 33134 22652 33140 22664
rect 33192 22652 33198 22704
rect 33502 22692 33508 22704
rect 33463 22664 33508 22692
rect 33502 22652 33508 22664
rect 33560 22652 33566 22704
rect 31018 22584 31024 22636
rect 31076 22624 31082 22636
rect 31206 22627 31264 22633
rect 31076 22596 31121 22624
rect 31076 22584 31082 22596
rect 31206 22593 31218 22627
rect 31252 22625 31264 22627
rect 31252 22624 31340 22625
rect 31386 22624 31392 22636
rect 31252 22597 31392 22624
rect 31252 22593 31264 22597
rect 31312 22596 31392 22597
rect 31206 22587 31264 22593
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 32674 22624 32680 22636
rect 32635 22596 32680 22624
rect 32674 22584 32680 22596
rect 32732 22584 32738 22636
rect 33686 22624 33692 22636
rect 33647 22596 33692 22624
rect 33686 22584 33692 22596
rect 33744 22584 33750 22636
rect 31110 22556 31116 22568
rect 30024 22528 30972 22556
rect 31071 22528 31116 22556
rect 26988 22488 27016 22516
rect 22204 22460 27016 22488
rect 22005 22451 22063 22457
rect 27982 22448 27988 22500
rect 28040 22488 28046 22500
rect 29748 22488 29776 22516
rect 30098 22488 30104 22500
rect 28040 22460 29776 22488
rect 30059 22460 30104 22488
rect 28040 22448 28046 22460
rect 30098 22448 30104 22460
rect 30156 22448 30162 22500
rect 23014 22420 23020 22432
rect 19904 22392 23020 22420
rect 23014 22380 23020 22392
rect 23072 22380 23078 22432
rect 24578 22420 24584 22432
rect 24539 22392 24584 22420
rect 24578 22380 24584 22392
rect 24636 22380 24642 22432
rect 26970 22380 26976 22432
rect 27028 22420 27034 22432
rect 27341 22423 27399 22429
rect 27341 22420 27353 22423
rect 27028 22392 27353 22420
rect 27028 22380 27034 22392
rect 27341 22389 27353 22392
rect 27387 22389 27399 22423
rect 27341 22383 27399 22389
rect 30374 22380 30380 22432
rect 30432 22420 30438 22432
rect 30837 22423 30895 22429
rect 30837 22420 30849 22423
rect 30432 22392 30849 22420
rect 30432 22380 30438 22392
rect 30837 22389 30849 22392
rect 30883 22389 30895 22423
rect 30944 22420 30972 22528
rect 31110 22516 31116 22528
rect 31168 22516 31174 22568
rect 31294 22516 31300 22568
rect 31352 22556 31358 22568
rect 31352 22528 31397 22556
rect 31352 22516 31358 22528
rect 32398 22516 32404 22568
rect 32456 22556 32462 22568
rect 32539 22559 32597 22565
rect 32539 22556 32551 22559
rect 32456 22528 32551 22556
rect 32456 22516 32462 22528
rect 32539 22525 32551 22528
rect 32585 22525 32597 22559
rect 32539 22519 32597 22525
rect 32953 22559 33011 22565
rect 32953 22525 32965 22559
rect 32999 22556 33011 22559
rect 33318 22556 33324 22568
rect 32999 22528 33324 22556
rect 32999 22525 33011 22528
rect 32953 22519 33011 22525
rect 33318 22516 33324 22528
rect 33376 22516 33382 22568
rect 33781 22423 33839 22429
rect 33781 22420 33793 22423
rect 30944 22392 33793 22420
rect 30837 22383 30895 22389
rect 33781 22389 33793 22392
rect 33827 22389 33839 22423
rect 33781 22383 33839 22389
rect 1104 22330 34868 22352
rect 1104 22278 5170 22330
rect 5222 22278 5234 22330
rect 5286 22278 5298 22330
rect 5350 22278 5362 22330
rect 5414 22278 5426 22330
rect 5478 22278 13611 22330
rect 13663 22278 13675 22330
rect 13727 22278 13739 22330
rect 13791 22278 13803 22330
rect 13855 22278 13867 22330
rect 13919 22278 22052 22330
rect 22104 22278 22116 22330
rect 22168 22278 22180 22330
rect 22232 22278 22244 22330
rect 22296 22278 22308 22330
rect 22360 22278 30493 22330
rect 30545 22278 30557 22330
rect 30609 22278 30621 22330
rect 30673 22278 30685 22330
rect 30737 22278 30749 22330
rect 30801 22278 34868 22330
rect 1104 22256 34868 22278
rect 4890 22176 4896 22228
rect 4948 22216 4954 22228
rect 9858 22216 9864 22228
rect 4948 22188 9864 22216
rect 4948 22176 4954 22188
rect 9858 22176 9864 22188
rect 9916 22176 9922 22228
rect 10226 22216 10232 22228
rect 10187 22188 10232 22216
rect 10226 22176 10232 22188
rect 10284 22216 10290 22228
rect 10962 22216 10968 22228
rect 10284 22188 10968 22216
rect 10284 22176 10290 22188
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 11698 22176 11704 22228
rect 11756 22225 11762 22228
rect 11756 22219 11771 22225
rect 11759 22185 11771 22219
rect 11756 22179 11771 22185
rect 11756 22176 11762 22179
rect 16390 22176 16396 22228
rect 16448 22216 16454 22228
rect 19978 22216 19984 22228
rect 16448 22188 19984 22216
rect 16448 22176 16454 22188
rect 19978 22176 19984 22188
rect 20036 22176 20042 22228
rect 23014 22216 23020 22228
rect 22975 22188 23020 22216
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 23201 22219 23259 22225
rect 23201 22185 23213 22219
rect 23247 22185 23259 22219
rect 23201 22179 23259 22185
rect 12809 22151 12867 22157
rect 12809 22117 12821 22151
rect 12855 22148 12867 22151
rect 13354 22148 13360 22160
rect 12855 22120 13360 22148
rect 12855 22117 12867 22120
rect 12809 22111 12867 22117
rect 13354 22108 13360 22120
rect 13412 22108 13418 22160
rect 17954 22108 17960 22160
rect 18012 22108 18018 22160
rect 22646 22108 22652 22160
rect 22704 22148 22710 22160
rect 23216 22148 23244 22179
rect 23842 22176 23848 22228
rect 23900 22216 23906 22228
rect 24762 22216 24768 22228
rect 23900 22188 24768 22216
rect 23900 22176 23906 22188
rect 24762 22176 24768 22188
rect 24820 22216 24826 22228
rect 28442 22216 28448 22228
rect 24820 22188 28448 22216
rect 24820 22176 24826 22188
rect 28442 22176 28448 22188
rect 28500 22176 28506 22228
rect 33505 22219 33563 22225
rect 33505 22185 33517 22219
rect 33551 22216 33563 22219
rect 33686 22216 33692 22228
rect 33551 22188 33692 22216
rect 33551 22185 33563 22188
rect 33505 22179 33563 22185
rect 33686 22176 33692 22188
rect 33744 22176 33750 22228
rect 24946 22148 24952 22160
rect 22704 22120 23244 22148
rect 24872 22120 24952 22148
rect 22704 22108 22710 22120
rect 11606 22040 11612 22092
rect 11664 22080 11670 22092
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11664 22052 11989 22080
rect 11664 22040 11670 22052
rect 11977 22049 11989 22052
rect 12023 22080 12035 22083
rect 12066 22080 12072 22092
rect 12023 22052 12072 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 17773 22083 17831 22089
rect 17773 22049 17785 22083
rect 17819 22080 17831 22083
rect 17972 22080 18000 22108
rect 17819 22052 18000 22080
rect 17819 22049 17831 22052
rect 17773 22043 17831 22049
rect 20070 22040 20076 22092
rect 20128 22080 20134 22092
rect 24872 22089 24900 22120
rect 24946 22108 24952 22120
rect 25004 22108 25010 22160
rect 30374 22148 30380 22160
rect 30024 22120 30380 22148
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 20128 22052 24777 22080
rect 20128 22040 20134 22052
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 24857 22083 24915 22089
rect 24857 22049 24869 22083
rect 24903 22049 24915 22083
rect 24857 22043 24915 22049
rect 25041 22083 25099 22089
rect 25041 22049 25053 22083
rect 25087 22080 25099 22083
rect 25222 22080 25228 22092
rect 25087 22052 25228 22080
rect 25087 22049 25099 22052
rect 25041 22043 25099 22049
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 26142 22040 26148 22092
rect 26200 22040 26206 22092
rect 26970 22080 26976 22092
rect 26252 22052 26976 22080
rect 7190 22012 7196 22024
rect 7103 21984 7196 22012
rect 7190 21972 7196 21984
rect 7248 22012 7254 22024
rect 7466 22012 7472 22024
rect 7248 21984 7472 22012
rect 7248 21972 7254 21984
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 9306 22012 9312 22024
rect 8619 21984 9312 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 12710 22012 12716 22024
rect 12671 21984 12716 22012
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 12894 22012 12900 22024
rect 12855 21984 12900 22012
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 12986 21972 12992 22024
rect 13044 22012 13050 22024
rect 17957 22015 18015 22021
rect 13044 21984 13089 22012
rect 13044 21972 13050 21984
rect 17957 21981 17969 22015
rect 18003 22012 18015 22015
rect 18046 22012 18052 22024
rect 18003 21984 18052 22012
rect 18003 21981 18015 21984
rect 17957 21975 18015 21981
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 22012 18383 22015
rect 18414 22012 18420 22024
rect 18371 21984 18420 22012
rect 18371 21981 18383 21984
rect 18325 21975 18383 21981
rect 18414 21972 18420 21984
rect 18472 22012 18478 22024
rect 19426 22012 19432 22024
rect 18472 21984 19432 22012
rect 18472 21972 18478 21984
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 19518 21972 19524 22024
rect 19576 22012 19582 22024
rect 19797 22015 19855 22021
rect 19797 22012 19809 22015
rect 19576 21984 19809 22012
rect 19576 21972 19582 21984
rect 19797 21981 19809 21984
rect 19843 21981 19855 22015
rect 19797 21975 19855 21981
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 20809 22015 20867 22021
rect 20809 22012 20821 22015
rect 20772 21984 20821 22012
rect 20772 21972 20778 21984
rect 20809 21981 20821 21984
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23201 22015 23259 22021
rect 23201 22012 23213 22015
rect 22980 21984 23213 22012
rect 22980 21972 22986 21984
rect 23201 21981 23213 21984
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 23385 22015 23443 22021
rect 23385 21981 23397 22015
rect 23431 22012 23443 22015
rect 24578 22012 24584 22024
rect 23431 21984 24584 22012
rect 23431 21981 23443 21984
rect 23385 21975 23443 21981
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 22012 25007 22015
rect 25958 22012 25964 22024
rect 24995 21984 25964 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 25958 21972 25964 21984
rect 26016 21972 26022 22024
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 22012 26111 22015
rect 26160 22012 26188 22040
rect 26252 22021 26280 22052
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 30024 22080 30052 22120
rect 30374 22108 30380 22120
rect 30432 22108 30438 22160
rect 30193 22083 30251 22089
rect 30193 22080 30205 22083
rect 30024 22052 30205 22080
rect 30193 22049 30205 22052
rect 30239 22049 30251 22083
rect 33134 22080 33140 22092
rect 33095 22052 33140 22080
rect 30193 22043 30251 22049
rect 33134 22040 33140 22052
rect 33192 22040 33198 22092
rect 26099 21984 26188 22012
rect 26237 22015 26295 22021
rect 26099 21981 26111 21984
rect 26053 21975 26111 21981
rect 26237 21981 26249 22015
rect 26283 21981 26295 22015
rect 26237 21975 26295 21981
rect 26326 21972 26332 22024
rect 26384 22012 26390 22024
rect 27062 22012 27068 22024
rect 26384 21984 27068 22012
rect 26384 21972 26390 21984
rect 27062 21972 27068 21984
rect 27120 21972 27126 22024
rect 27801 22015 27859 22021
rect 27801 21981 27813 22015
rect 27847 22012 27859 22015
rect 28629 22015 28687 22021
rect 28629 22012 28641 22015
rect 27847 21984 28641 22012
rect 27847 21981 27859 21984
rect 27801 21975 27859 21981
rect 28629 21981 28641 21984
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 21981 30159 22015
rect 31018 22012 31024 22024
rect 30979 21984 31024 22012
rect 30101 21975 30159 21981
rect 11698 21944 11704 21956
rect 11270 21916 11704 21944
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 19334 21904 19340 21956
rect 19392 21944 19398 21956
rect 19886 21944 19892 21956
rect 19392 21916 19892 21944
rect 19392 21904 19398 21916
rect 19886 21904 19892 21916
rect 19944 21944 19950 21956
rect 20165 21947 20223 21953
rect 20165 21944 20177 21947
rect 19944 21916 20177 21944
rect 19944 21904 19950 21916
rect 20165 21913 20177 21916
rect 20211 21944 20223 21947
rect 20211 21916 22508 21944
rect 20211 21913 20223 21916
rect 20165 21907 20223 21913
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7190 21876 7196 21888
rect 6972 21848 7196 21876
rect 6972 21836 6978 21848
rect 7190 21836 7196 21848
rect 7248 21836 7254 21888
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 8481 21879 8539 21885
rect 8481 21876 8493 21879
rect 8444 21848 8493 21876
rect 8444 21836 8450 21848
rect 8481 21845 8493 21848
rect 8527 21876 8539 21879
rect 9030 21876 9036 21888
rect 8527 21848 9036 21876
rect 8527 21845 8539 21848
rect 8481 21839 8539 21845
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 10686 21836 10692 21888
rect 10744 21876 10750 21888
rect 12529 21879 12587 21885
rect 12529 21876 12541 21879
rect 10744 21848 12541 21876
rect 10744 21836 10750 21848
rect 12529 21845 12541 21848
rect 12575 21845 12587 21879
rect 12529 21839 12587 21845
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 19610 21876 19616 21888
rect 18279 21848 19616 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 19610 21836 19616 21848
rect 19668 21836 19674 21888
rect 22278 21876 22284 21888
rect 22239 21848 22284 21876
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 22480 21876 22508 21916
rect 23106 21904 23112 21956
rect 23164 21944 23170 21956
rect 26145 21947 26203 21953
rect 23164 21916 25360 21944
rect 23164 21904 23170 21916
rect 24946 21876 24952 21888
rect 22480 21848 24952 21876
rect 24946 21836 24952 21848
rect 25004 21836 25010 21888
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 25096 21848 25237 21876
rect 25096 21836 25102 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25332 21876 25360 21916
rect 26145 21913 26157 21947
rect 26191 21944 26203 21947
rect 27522 21944 27528 21956
rect 26191 21916 27528 21944
rect 26191 21913 26203 21916
rect 26145 21907 26203 21913
rect 27522 21904 27528 21916
rect 27580 21944 27586 21956
rect 28261 21947 28319 21953
rect 28261 21944 28273 21947
rect 27580 21916 28273 21944
rect 27580 21904 27586 21916
rect 28261 21913 28273 21916
rect 28307 21913 28319 21947
rect 28442 21944 28448 21956
rect 28403 21916 28448 21944
rect 28261 21907 28319 21913
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 30116 21944 30144 21975
rect 31018 21972 31024 21984
rect 31076 22012 31082 22024
rect 31386 22012 31392 22024
rect 31076 21984 31248 22012
rect 31347 21984 31392 22012
rect 31076 21972 31082 21984
rect 30282 21944 30288 21956
rect 30116 21916 30288 21944
rect 30282 21904 30288 21916
rect 30340 21944 30346 21956
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 30340 21916 31125 21944
rect 30340 21904 30346 21916
rect 31113 21913 31125 21916
rect 31159 21913 31171 21947
rect 31220 21944 31248 21984
rect 31386 21972 31392 21984
rect 31444 21972 31450 22024
rect 31570 22012 31576 22024
rect 31531 21984 31576 22012
rect 31570 21972 31576 21984
rect 31628 22012 31634 22024
rect 32033 22015 32091 22021
rect 32033 22012 32045 22015
rect 31628 21984 32045 22012
rect 31628 21972 31634 21984
rect 32033 21981 32045 21984
rect 32079 21981 32091 22015
rect 32398 22012 32404 22024
rect 32359 21984 32404 22012
rect 32033 21975 32091 21981
rect 32398 21972 32404 21984
rect 32456 21972 32462 22024
rect 32582 22012 32588 22024
rect 32543 21984 32588 22012
rect 32582 21972 32588 21984
rect 32640 21972 32646 22024
rect 33318 22012 33324 22024
rect 33279 21984 33324 22012
rect 33318 21972 33324 21984
rect 33376 21972 33382 22024
rect 32125 21947 32183 21953
rect 32125 21944 32137 21947
rect 31220 21916 32137 21944
rect 31113 21907 31171 21913
rect 32125 21913 32137 21916
rect 32171 21913 32183 21947
rect 32125 21907 32183 21913
rect 27709 21879 27767 21885
rect 27709 21876 27721 21879
rect 25332 21848 27721 21876
rect 25225 21839 25283 21845
rect 27709 21845 27721 21848
rect 27755 21845 27767 21879
rect 29730 21876 29736 21888
rect 29691 21848 29736 21876
rect 27709 21839 27767 21845
rect 29730 21836 29736 21848
rect 29788 21836 29794 21888
rect 1104 21786 35027 21808
rect 1104 21734 9390 21786
rect 9442 21734 9454 21786
rect 9506 21734 9518 21786
rect 9570 21734 9582 21786
rect 9634 21734 9646 21786
rect 9698 21734 17831 21786
rect 17883 21734 17895 21786
rect 17947 21734 17959 21786
rect 18011 21734 18023 21786
rect 18075 21734 18087 21786
rect 18139 21734 26272 21786
rect 26324 21734 26336 21786
rect 26388 21734 26400 21786
rect 26452 21734 26464 21786
rect 26516 21734 26528 21786
rect 26580 21734 34713 21786
rect 34765 21734 34777 21786
rect 34829 21734 34841 21786
rect 34893 21734 34905 21786
rect 34957 21734 34969 21786
rect 35021 21734 35027 21786
rect 1104 21712 35027 21734
rect 12710 21632 12716 21684
rect 12768 21672 12774 21684
rect 27154 21672 27160 21684
rect 12768 21644 23244 21672
rect 27115 21644 27160 21672
rect 12768 21632 12774 21644
rect 11698 21604 11704 21616
rect 11659 21576 11704 21604
rect 11698 21564 11704 21576
rect 11756 21564 11762 21616
rect 20438 21604 20444 21616
rect 19444 21576 20444 21604
rect 19444 21548 19472 21576
rect 20438 21564 20444 21576
rect 20496 21564 20502 21616
rect 23106 21604 23112 21616
rect 20548 21576 23112 21604
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 2915 21508 3801 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 3789 21505 3801 21508
rect 3835 21536 3847 21539
rect 3970 21536 3976 21548
rect 3835 21508 3976 21536
rect 3835 21505 3847 21508
rect 3789 21499 3847 21505
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21536 4123 21539
rect 4154 21536 4160 21548
rect 4111 21508 4160 21536
rect 4111 21505 4123 21508
rect 4065 21499 4123 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 11790 21536 11796 21548
rect 11751 21508 11796 21536
rect 11790 21496 11796 21508
rect 11848 21496 11854 21548
rect 11974 21496 11980 21548
rect 12032 21536 12038 21548
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 12032 21508 12081 21536
rect 12032 21496 12038 21508
rect 12069 21505 12081 21508
rect 12115 21536 12127 21539
rect 12342 21536 12348 21548
rect 12115 21508 12348 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 14056 21508 14473 21536
rect 14056 21496 14062 21508
rect 14461 21505 14473 21508
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21536 14611 21539
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 14599 21508 15301 21536
rect 14599 21505 14611 21508
rect 14553 21499 14611 21505
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21536 15531 21539
rect 16022 21536 16028 21548
rect 15519 21508 16028 21536
rect 15519 21505 15531 21508
rect 15473 21499 15531 21505
rect 16022 21496 16028 21508
rect 16080 21536 16086 21548
rect 16482 21536 16488 21548
rect 16080 21508 16488 21536
rect 16080 21496 16086 21508
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 19426 21536 19432 21548
rect 19339 21508 19432 21536
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 19794 21536 19800 21548
rect 19755 21508 19800 21536
rect 19794 21496 19800 21508
rect 19852 21496 19858 21548
rect 20548 21545 20576 21576
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20625 21539 20683 21545
rect 20625 21505 20637 21539
rect 20671 21505 20683 21539
rect 20625 21499 20683 21505
rect 22005 21539 22063 21545
rect 22005 21505 22017 21539
rect 22051 21505 22063 21539
rect 22278 21536 22284 21548
rect 22239 21508 22284 21536
rect 22005 21499 22063 21505
rect 2958 21468 2964 21480
rect 2919 21440 2964 21468
rect 2958 21428 2964 21440
rect 3016 21428 3022 21480
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21468 3203 21471
rect 3191 21440 4016 21468
rect 3191 21437 3203 21440
rect 3145 21431 3203 21437
rect 2976 21400 3004 21428
rect 3988 21409 4016 21440
rect 10962 21428 10968 21480
rect 11020 21468 11026 21480
rect 19521 21471 19579 21477
rect 19521 21468 19533 21471
rect 11020 21440 19533 21468
rect 11020 21428 11026 21440
rect 19521 21437 19533 21440
rect 19567 21437 19579 21471
rect 19521 21431 19579 21437
rect 19610 21428 19616 21480
rect 19668 21468 19674 21480
rect 20640 21468 20668 21499
rect 19668 21440 20668 21468
rect 19668 21428 19674 21440
rect 3881 21403 3939 21409
rect 3881 21400 3893 21403
rect 2976 21372 3893 21400
rect 3881 21369 3893 21372
rect 3927 21369 3939 21403
rect 3881 21363 3939 21369
rect 3973 21403 4031 21409
rect 3973 21369 3985 21403
rect 4019 21400 4031 21403
rect 4062 21400 4068 21412
rect 4019 21372 4068 21400
rect 4019 21369 4031 21372
rect 3973 21363 4031 21369
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 3050 21332 3056 21344
rect 3011 21304 3056 21332
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 3602 21332 3608 21344
rect 3563 21304 3608 21332
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21332 15531 21335
rect 16850 21332 16856 21344
rect 15519 21304 16856 21332
rect 15519 21301 15531 21304
rect 15473 21295 15531 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 19886 21292 19892 21344
rect 19944 21332 19950 21344
rect 22020 21332 22048 21499
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 23216 21536 23244 21644
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 30098 21672 30104 21684
rect 27264 21644 30104 21672
rect 27264 21536 27292 21644
rect 30098 21632 30104 21644
rect 30156 21632 30162 21684
rect 30282 21672 30288 21684
rect 30243 21644 30288 21672
rect 30282 21632 30288 21644
rect 30340 21632 30346 21684
rect 31665 21675 31723 21681
rect 31665 21641 31677 21675
rect 31711 21672 31723 21675
rect 31754 21672 31760 21684
rect 31711 21644 31760 21672
rect 31711 21641 31723 21644
rect 31665 21635 31723 21641
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 28442 21604 28448 21616
rect 28184 21576 28448 21604
rect 23216 21508 27292 21536
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 27982 21536 27988 21548
rect 27571 21508 27988 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 28184 21545 28212 21576
rect 28442 21564 28448 21576
rect 28500 21564 28506 21616
rect 30469 21607 30527 21613
rect 30469 21573 30481 21607
rect 30515 21604 30527 21607
rect 31018 21604 31024 21616
rect 30515 21576 31024 21604
rect 30515 21573 30527 21576
rect 30469 21567 30527 21573
rect 31018 21564 31024 21576
rect 31076 21564 31082 21616
rect 31386 21564 31392 21616
rect 31444 21604 31450 21616
rect 31444 21576 31708 21604
rect 31444 21564 31450 21576
rect 28169 21539 28227 21545
rect 28169 21505 28181 21539
rect 28215 21505 28227 21539
rect 28169 21499 28227 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21536 28411 21539
rect 29730 21536 29736 21548
rect 28399 21508 29736 21536
rect 28399 21505 28411 21508
rect 28353 21499 28411 21505
rect 29730 21496 29736 21508
rect 29788 21496 29794 21548
rect 30193 21539 30251 21545
rect 30193 21505 30205 21539
rect 30239 21536 30251 21539
rect 30374 21536 30380 21548
rect 30239 21508 30380 21536
rect 30239 21505 30251 21508
rect 30193 21499 30251 21505
rect 30374 21496 30380 21508
rect 30432 21496 30438 21548
rect 31110 21496 31116 21548
rect 31168 21536 31174 21548
rect 31680 21545 31708 21576
rect 31481 21539 31539 21545
rect 31481 21536 31493 21539
rect 31168 21508 31493 21536
rect 31168 21496 31174 21508
rect 31481 21505 31493 21508
rect 31527 21505 31539 21539
rect 31481 21499 31539 21505
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21536 31723 21539
rect 32582 21536 32588 21548
rect 31711 21508 32588 21536
rect 31711 21505 31723 21508
rect 31665 21499 31723 21505
rect 32582 21496 32588 21508
rect 32640 21496 32646 21548
rect 22370 21468 22376 21480
rect 22331 21440 22376 21468
rect 22370 21428 22376 21440
rect 22428 21428 22434 21480
rect 23198 21468 23204 21480
rect 23159 21440 23204 21468
rect 23198 21428 23204 21440
rect 23256 21428 23262 21480
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 23566 21468 23572 21480
rect 23523 21440 23572 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 27614 21468 27620 21480
rect 27575 21440 27620 21468
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 24765 21403 24823 21409
rect 24765 21369 24777 21403
rect 24811 21400 24823 21403
rect 30098 21400 30104 21412
rect 24811 21372 30104 21400
rect 24811 21369 24823 21372
rect 24765 21363 24823 21369
rect 23842 21332 23848 21344
rect 19944 21304 23848 21332
rect 19944 21292 19950 21304
rect 23842 21292 23848 21304
rect 23900 21292 23906 21344
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 24780 21332 24808 21363
rect 30098 21360 30104 21372
rect 30156 21400 30162 21412
rect 32214 21400 32220 21412
rect 30156 21372 32220 21400
rect 30156 21360 30162 21372
rect 32214 21360 32220 21372
rect 32272 21360 32278 21412
rect 23992 21304 24808 21332
rect 23992 21292 23998 21304
rect 27890 21292 27896 21344
rect 27948 21332 27954 21344
rect 28353 21335 28411 21341
rect 28353 21332 28365 21335
rect 27948 21304 28365 21332
rect 27948 21292 27954 21304
rect 28353 21301 28365 21304
rect 28399 21301 28411 21335
rect 28353 21295 28411 21301
rect 28442 21292 28448 21344
rect 28500 21332 28506 21344
rect 30469 21335 30527 21341
rect 30469 21332 30481 21335
rect 28500 21304 30481 21332
rect 28500 21292 28506 21304
rect 30469 21301 30481 21304
rect 30515 21301 30527 21335
rect 30469 21295 30527 21301
rect 1104 21242 34868 21264
rect 1104 21190 5170 21242
rect 5222 21190 5234 21242
rect 5286 21190 5298 21242
rect 5350 21190 5362 21242
rect 5414 21190 5426 21242
rect 5478 21190 13611 21242
rect 13663 21190 13675 21242
rect 13727 21190 13739 21242
rect 13791 21190 13803 21242
rect 13855 21190 13867 21242
rect 13919 21190 22052 21242
rect 22104 21190 22116 21242
rect 22168 21190 22180 21242
rect 22232 21190 22244 21242
rect 22296 21190 22308 21242
rect 22360 21190 30493 21242
rect 30545 21190 30557 21242
rect 30609 21190 30621 21242
rect 30673 21190 30685 21242
rect 30737 21190 30749 21242
rect 30801 21190 34868 21242
rect 1104 21168 34868 21190
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 13449 21131 13507 21137
rect 13449 21128 13461 21131
rect 12952 21100 13461 21128
rect 12952 21088 12958 21100
rect 13449 21097 13461 21100
rect 13495 21097 13507 21131
rect 13449 21091 13507 21097
rect 14645 21131 14703 21137
rect 14645 21097 14657 21131
rect 14691 21097 14703 21131
rect 14645 21091 14703 21097
rect 16117 21131 16175 21137
rect 16117 21097 16129 21131
rect 16163 21128 16175 21131
rect 17310 21128 17316 21140
rect 16163 21100 17316 21128
rect 16163 21097 16175 21100
rect 16117 21091 16175 21097
rect 7377 20995 7435 21001
rect 7377 20961 7389 20995
rect 7423 20992 7435 20995
rect 7466 20992 7472 21004
rect 7423 20964 7472 20992
rect 7423 20961 7435 20964
rect 7377 20955 7435 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 3234 20924 3240 20936
rect 3195 20896 3240 20924
rect 3234 20884 3240 20896
rect 3292 20884 3298 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 3694 20924 3700 20936
rect 3467 20896 3700 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 3694 20884 3700 20896
rect 3752 20884 3758 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7340 20896 7573 20924
rect 7340 20884 7346 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 7708 20896 7753 20924
rect 7708 20884 7714 20896
rect 10318 20884 10324 20936
rect 10376 20924 10382 20936
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 10376 20896 10425 20924
rect 10376 20884 10382 20896
rect 10413 20893 10425 20896
rect 10459 20893 10471 20927
rect 10686 20924 10692 20936
rect 10647 20896 10692 20924
rect 10413 20887 10471 20893
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 13446 20884 13452 20936
rect 13504 20924 13510 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13504 20896 13553 20924
rect 13504 20884 13510 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 14553 20927 14611 20933
rect 14553 20924 14565 20927
rect 14516 20896 14565 20924
rect 14516 20884 14522 20896
rect 14553 20893 14565 20896
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 14660 20856 14688 21091
rect 17310 21088 17316 21100
rect 17368 21088 17374 21140
rect 21266 21128 21272 21140
rect 21227 21100 21272 21128
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 23566 21128 23572 21140
rect 23527 21100 23572 21128
rect 23566 21088 23572 21100
rect 23624 21088 23630 21140
rect 24946 21088 24952 21140
rect 25004 21128 25010 21140
rect 30926 21128 30932 21140
rect 25004 21100 30932 21128
rect 25004 21088 25010 21100
rect 30926 21088 30932 21100
rect 30984 21088 30990 21140
rect 31938 21128 31944 21140
rect 31588 21100 31944 21128
rect 19521 21063 19579 21069
rect 19521 21029 19533 21063
rect 19567 21029 19579 21063
rect 31588 21060 31616 21100
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 32398 21128 32404 21140
rect 32359 21100 32404 21128
rect 32398 21088 32404 21100
rect 32456 21088 32462 21140
rect 33137 21063 33195 21069
rect 33137 21060 33149 21063
rect 19521 21023 19579 21029
rect 23768 21032 31616 21060
rect 31680 21032 33149 21060
rect 19536 20992 19564 21023
rect 14752 20964 19564 20992
rect 19705 20995 19763 21001
rect 14752 20933 14780 20964
rect 19705 20961 19717 20995
rect 19751 20992 19763 20995
rect 19886 20992 19892 21004
rect 19751 20964 19892 20992
rect 19751 20961 19763 20964
rect 19705 20955 19763 20961
rect 19886 20952 19892 20964
rect 19944 20952 19950 21004
rect 19978 20952 19984 21004
rect 20036 20992 20042 21004
rect 20073 20995 20131 21001
rect 20073 20992 20085 20995
rect 20036 20964 20085 20992
rect 20036 20952 20042 20964
rect 20073 20961 20085 20964
rect 20119 20961 20131 20995
rect 20073 20955 20131 20961
rect 20165 20995 20223 21001
rect 20165 20961 20177 20995
rect 20211 20992 20223 20995
rect 21174 20992 21180 21004
rect 20211 20964 21180 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 21174 20952 21180 20964
rect 21232 20952 21238 21004
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20924 17463 20927
rect 18322 20924 18328 20936
rect 17451 20896 18328 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 19794 20924 19800 20936
rect 19755 20896 19800 20924
rect 19794 20884 19800 20896
rect 19852 20884 19858 20936
rect 22554 20924 22560 20936
rect 22515 20896 22560 20924
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 23768 20933 23796 21032
rect 24946 20992 24952 21004
rect 24799 20964 24952 20992
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 22664 20896 23765 20924
rect 14660 20828 14872 20856
rect 3142 20748 3148 20800
rect 3200 20788 3206 20800
rect 3329 20791 3387 20797
rect 3329 20788 3341 20791
rect 3200 20760 3341 20788
rect 3200 20748 3206 20760
rect 3329 20757 3341 20760
rect 3375 20757 3387 20791
rect 7374 20788 7380 20800
rect 7335 20760 7380 20788
rect 3329 20751 3387 20757
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 10226 20788 10232 20800
rect 10187 20760 10232 20788
rect 10226 20748 10232 20760
rect 10284 20748 10290 20800
rect 10597 20791 10655 20797
rect 10597 20757 10609 20791
rect 10643 20788 10655 20791
rect 10962 20788 10968 20800
rect 10643 20760 10968 20788
rect 10643 20757 10655 20760
rect 10597 20751 10655 20757
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 14366 20788 14372 20800
rect 14327 20760 14372 20788
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 14844 20788 14872 20828
rect 19702 20816 19708 20868
rect 19760 20856 19766 20868
rect 22664 20856 22692 20896
rect 23753 20893 23765 20896
rect 23799 20893 23811 20927
rect 23934 20924 23940 20936
rect 23895 20896 23940 20924
rect 23753 20887 23811 20893
rect 23934 20884 23940 20896
rect 23992 20884 23998 20936
rect 24799 20933 24827 20964
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 31110 20952 31116 21004
rect 31168 20992 31174 21004
rect 31297 20995 31355 21001
rect 31297 20992 31309 20995
rect 31168 20964 31309 20992
rect 31168 20952 31174 20964
rect 31297 20961 31309 20964
rect 31343 20961 31355 20995
rect 31297 20955 31355 20961
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20924 24087 20927
rect 24784 20927 24842 20933
rect 24075 20896 24716 20924
rect 24075 20893 24087 20896
rect 24029 20887 24087 20893
rect 19760 20828 22692 20856
rect 19760 20816 19766 20828
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 23440 20828 24593 20856
rect 23440 20816 23446 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24688 20856 24716 20896
rect 24784 20893 24796 20927
rect 24830 20893 24842 20927
rect 24784 20887 24842 20893
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20924 25099 20927
rect 25130 20924 25136 20936
rect 25087 20896 25136 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 25056 20856 25084 20887
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 31680 20933 31708 21032
rect 33137 21029 33149 21032
rect 33183 21029 33195 21063
rect 33137 21023 33195 21029
rect 31572 20927 31630 20933
rect 31572 20893 31584 20927
rect 31618 20893 31630 20927
rect 31572 20887 31630 20893
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20893 31723 20927
rect 32214 20924 32220 20936
rect 32175 20896 32220 20924
rect 31665 20887 31723 20893
rect 24688 20828 25084 20856
rect 31588 20856 31616 20887
rect 32214 20884 32220 20896
rect 32272 20884 32278 20936
rect 32490 20924 32496 20936
rect 32451 20896 32496 20924
rect 32490 20884 32496 20896
rect 32548 20884 32554 20936
rect 32950 20924 32956 20936
rect 32911 20896 32956 20924
rect 32950 20884 32956 20896
rect 33008 20884 33014 20936
rect 33042 20884 33048 20936
rect 33100 20924 33106 20936
rect 33137 20927 33195 20933
rect 33137 20924 33149 20927
rect 33100 20896 33149 20924
rect 33100 20884 33106 20896
rect 33137 20893 33149 20896
rect 33183 20893 33195 20927
rect 33137 20887 33195 20893
rect 32766 20856 32772 20868
rect 31588 20828 32772 20856
rect 24581 20819 24639 20825
rect 32766 20816 32772 20828
rect 32824 20816 32830 20868
rect 22554 20788 22560 20800
rect 14844 20760 22560 20788
rect 22554 20748 22560 20760
rect 22612 20748 22618 20800
rect 24949 20791 25007 20797
rect 24949 20757 24961 20791
rect 24995 20788 25007 20791
rect 25222 20788 25228 20800
rect 24995 20760 25228 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 1104 20698 35027 20720
rect 1104 20646 9390 20698
rect 9442 20646 9454 20698
rect 9506 20646 9518 20698
rect 9570 20646 9582 20698
rect 9634 20646 9646 20698
rect 9698 20646 17831 20698
rect 17883 20646 17895 20698
rect 17947 20646 17959 20698
rect 18011 20646 18023 20698
rect 18075 20646 18087 20698
rect 18139 20646 26272 20698
rect 26324 20646 26336 20698
rect 26388 20646 26400 20698
rect 26452 20646 26464 20698
rect 26516 20646 26528 20698
rect 26580 20646 34713 20698
rect 34765 20646 34777 20698
rect 34829 20646 34841 20698
rect 34893 20646 34905 20698
rect 34957 20646 34969 20698
rect 35021 20646 35027 20698
rect 1104 20624 35027 20646
rect 7837 20587 7895 20593
rect 7837 20553 7849 20587
rect 7883 20584 7895 20587
rect 8294 20584 8300 20596
rect 7883 20556 8300 20584
rect 7883 20553 7895 20556
rect 7837 20547 7895 20553
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 8389 20587 8447 20593
rect 8389 20553 8401 20587
rect 8435 20553 8447 20587
rect 14182 20584 14188 20596
rect 8389 20547 8447 20553
rect 13280 20556 14188 20584
rect 3602 20516 3608 20528
rect 3563 20488 3608 20516
rect 3602 20476 3608 20488
rect 3660 20476 3666 20528
rect 7469 20519 7527 20525
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 7742 20516 7748 20528
rect 7515 20488 7748 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 7742 20476 7748 20488
rect 7800 20516 7806 20528
rect 8404 20516 8432 20547
rect 7800 20488 8432 20516
rect 7800 20476 7806 20488
rect 3142 20448 3148 20460
rect 3103 20420 3148 20448
rect 3142 20408 3148 20420
rect 3200 20408 3206 20460
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3970 20448 3976 20460
rect 3283 20420 3976 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4522 20448 4528 20460
rect 4479 20420 4528 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 7340 20420 7389 20448
rect 7340 20408 7346 20420
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20448 7711 20451
rect 8018 20448 8024 20460
rect 7699 20420 8024 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8478 20448 8484 20460
rect 8439 20420 8484 20448
rect 8297 20411 8355 20417
rect 3050 20340 3056 20392
rect 3108 20380 3114 20392
rect 3418 20380 3424 20392
rect 3108 20352 3424 20380
rect 3108 20340 3114 20352
rect 3418 20340 3424 20352
rect 3476 20380 3482 20392
rect 3513 20383 3571 20389
rect 3513 20380 3525 20383
rect 3476 20352 3525 20380
rect 3476 20340 3482 20352
rect 3513 20349 3525 20352
rect 3559 20349 3571 20383
rect 4062 20380 4068 20392
rect 4023 20352 4068 20380
rect 3513 20343 3571 20349
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20349 4399 20383
rect 8312 20380 8340 20411
rect 8478 20408 8484 20420
rect 8536 20408 8542 20460
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 10226 20448 10232 20460
rect 8619 20420 10232 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 11054 20448 11060 20460
rect 11015 20420 11060 20448
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 13280 20457 13308 20556
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 19058 20584 19064 20596
rect 18340 20556 19064 20584
rect 14366 20516 14372 20528
rect 13464 20488 14372 20516
rect 13464 20457 13492 20488
rect 14366 20476 14372 20488
rect 14424 20476 14430 20528
rect 16206 20516 16212 20528
rect 14476 20488 16212 20516
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13449 20411 13507 20417
rect 13556 20420 13829 20448
rect 8938 20380 8944 20392
rect 8312 20352 8944 20380
rect 4341 20343 4399 20349
rect 2406 20272 2412 20324
rect 2464 20312 2470 20324
rect 4356 20312 4384 20343
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 10318 20380 10324 20392
rect 10279 20352 10324 20380
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 12406 20352 12817 20380
rect 2464 20284 4384 20312
rect 2464 20272 2470 20284
rect 7834 20272 7840 20324
rect 7892 20312 7898 20324
rect 12406 20312 12434 20352
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 13556 20380 13584 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 13817 20411 13875 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20448 14059 20451
rect 14476 20448 14504 20488
rect 16206 20476 16212 20488
rect 16264 20476 16270 20528
rect 14047 20420 14504 20448
rect 15105 20451 15163 20457
rect 14047 20417 14059 20420
rect 14001 20411 14059 20417
rect 15105 20417 15117 20451
rect 15151 20417 15163 20451
rect 15654 20448 15660 20460
rect 15615 20420 15660 20448
rect 15105 20411 15163 20417
rect 13412 20352 13584 20380
rect 13412 20340 13418 20352
rect 7892 20284 12434 20312
rect 7892 20272 7898 20284
rect 12894 20272 12900 20324
rect 12952 20312 12958 20324
rect 14016 20312 14044 20411
rect 14182 20340 14188 20392
rect 14240 20380 14246 20392
rect 14642 20380 14648 20392
rect 14240 20352 14648 20380
rect 14240 20340 14246 20352
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15120 20380 15148 20411
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16022 20448 16028 20460
rect 15887 20420 16028 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 18340 20457 18368 20556
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19153 20587 19211 20593
rect 19153 20553 19165 20587
rect 19199 20584 19211 20587
rect 19610 20584 19616 20596
rect 19199 20556 19616 20584
rect 19199 20553 19211 20556
rect 19153 20547 19211 20553
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 19794 20544 19800 20596
rect 19852 20584 19858 20596
rect 21085 20587 21143 20593
rect 19852 20556 20852 20584
rect 19852 20544 19858 20556
rect 18782 20516 18788 20528
rect 18432 20488 18788 20516
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18432 20380 18460 20488
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 20824 20525 20852 20556
rect 21085 20553 21097 20587
rect 21131 20584 21143 20587
rect 22738 20584 22744 20596
rect 21131 20556 22744 20584
rect 21131 20553 21143 20556
rect 21085 20547 21143 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 31570 20584 31576 20596
rect 31531 20556 31576 20584
rect 31570 20544 31576 20556
rect 31628 20544 31634 20596
rect 32582 20584 32588 20596
rect 32543 20556 32588 20584
rect 32582 20544 32588 20556
rect 32640 20544 32646 20596
rect 20809 20519 20867 20525
rect 20809 20485 20821 20519
rect 20855 20485 20867 20519
rect 20809 20479 20867 20485
rect 22370 20476 22376 20528
rect 22428 20516 22434 20528
rect 23201 20519 23259 20525
rect 23201 20516 23213 20519
rect 22428 20488 23213 20516
rect 22428 20476 22434 20488
rect 23201 20485 23213 20488
rect 23247 20485 23259 20519
rect 23201 20479 23259 20485
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20448 18659 20451
rect 18966 20448 18972 20460
rect 18647 20420 18972 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 14792 20352 18460 20380
rect 18524 20380 18552 20411
rect 18966 20408 18972 20420
rect 19024 20448 19030 20460
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 19024 20420 19073 20448
rect 19024 20408 19030 20420
rect 19061 20417 19073 20420
rect 19107 20448 19119 20451
rect 19150 20448 19156 20460
rect 19107 20420 19156 20448
rect 19107 20417 19119 20420
rect 19061 20411 19119 20417
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19702 20448 19708 20460
rect 19392 20420 19708 20448
rect 19392 20408 19398 20420
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 20438 20408 20444 20460
rect 20496 20448 20502 20460
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 20496 20420 20545 20448
rect 20496 20408 20502 20420
rect 20533 20417 20545 20420
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 20717 20451 20775 20457
rect 20717 20448 20729 20451
rect 20680 20420 20729 20448
rect 20680 20408 20686 20420
rect 20717 20417 20729 20420
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 20947 20451 21005 20457
rect 20947 20417 20959 20451
rect 20993 20448 21005 20451
rect 21082 20448 21088 20460
rect 20993 20420 21088 20448
rect 20993 20417 21005 20420
rect 20947 20411 21005 20417
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 27982 20448 27988 20460
rect 27943 20420 27988 20448
rect 27982 20408 27988 20420
rect 28040 20408 28046 20460
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20448 31815 20451
rect 32398 20448 32404 20460
rect 31803 20420 32404 20448
rect 31803 20417 31815 20420
rect 31757 20411 31815 20417
rect 19794 20380 19800 20392
rect 18524 20352 19800 20380
rect 14792 20340 14798 20352
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 25866 20380 25872 20392
rect 22612 20352 25872 20380
rect 22612 20340 22618 20352
rect 25866 20340 25872 20352
rect 25924 20340 25930 20392
rect 27890 20380 27896 20392
rect 27851 20352 27896 20380
rect 27890 20340 27896 20352
rect 27948 20340 27954 20392
rect 31588 20380 31616 20411
rect 32398 20408 32404 20420
rect 32456 20408 32462 20460
rect 32766 20448 32772 20460
rect 32727 20420 32772 20448
rect 32766 20408 32772 20420
rect 32824 20408 32830 20460
rect 33042 20448 33048 20460
rect 33003 20420 33048 20448
rect 33042 20408 33048 20420
rect 33100 20408 33106 20460
rect 31938 20380 31944 20392
rect 31588 20352 31944 20380
rect 31938 20340 31944 20352
rect 31996 20340 32002 20392
rect 12952 20284 14044 20312
rect 12952 20272 12958 20284
rect 16666 20272 16672 20324
rect 16724 20312 16730 20324
rect 20254 20312 20260 20324
rect 16724 20284 20260 20312
rect 16724 20272 16730 20284
rect 20254 20272 20260 20284
rect 20312 20272 20318 20324
rect 21358 20272 21364 20324
rect 21416 20312 21422 20324
rect 27617 20315 27675 20321
rect 27617 20312 27629 20315
rect 21416 20284 27629 20312
rect 21416 20272 21422 20284
rect 27617 20281 27629 20284
rect 27663 20281 27675 20315
rect 27617 20275 27675 20281
rect 32306 20272 32312 20324
rect 32364 20312 32370 20324
rect 32950 20312 32956 20324
rect 32364 20284 32956 20312
rect 32364 20272 32370 20284
rect 32950 20272 32956 20284
rect 33008 20272 33014 20324
rect 2958 20244 2964 20256
rect 2919 20216 2964 20244
rect 2958 20204 2964 20216
rect 3016 20204 3022 20256
rect 15838 20244 15844 20256
rect 15799 20216 15844 20244
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 18141 20247 18199 20253
rect 18141 20213 18153 20247
rect 18187 20244 18199 20247
rect 19058 20244 19064 20256
rect 18187 20216 19064 20244
rect 18187 20213 18199 20216
rect 18141 20207 18199 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19521 20247 19579 20253
rect 19521 20213 19533 20247
rect 19567 20244 19579 20247
rect 19702 20244 19708 20256
rect 19567 20216 19708 20244
rect 19567 20213 19579 20216
rect 19521 20207 19579 20213
rect 19702 20204 19708 20216
rect 19760 20204 19766 20256
rect 21726 20204 21732 20256
rect 21784 20244 21790 20256
rect 24489 20247 24547 20253
rect 24489 20244 24501 20247
rect 21784 20216 24501 20244
rect 21784 20204 21790 20216
rect 24489 20213 24501 20216
rect 24535 20213 24547 20247
rect 24489 20207 24547 20213
rect 27985 20247 28043 20253
rect 27985 20213 27997 20247
rect 28031 20244 28043 20247
rect 28074 20244 28080 20256
rect 28031 20216 28080 20244
rect 28031 20213 28043 20216
rect 27985 20207 28043 20213
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 1104 20154 34868 20176
rect 1104 20102 5170 20154
rect 5222 20102 5234 20154
rect 5286 20102 5298 20154
rect 5350 20102 5362 20154
rect 5414 20102 5426 20154
rect 5478 20102 13611 20154
rect 13663 20102 13675 20154
rect 13727 20102 13739 20154
rect 13791 20102 13803 20154
rect 13855 20102 13867 20154
rect 13919 20102 22052 20154
rect 22104 20102 22116 20154
rect 22168 20102 22180 20154
rect 22232 20102 22244 20154
rect 22296 20102 22308 20154
rect 22360 20102 30493 20154
rect 30545 20102 30557 20154
rect 30609 20102 30621 20154
rect 30673 20102 30685 20154
rect 30737 20102 30749 20154
rect 30801 20102 34868 20154
rect 1104 20080 34868 20102
rect 3970 20040 3976 20052
rect 3931 20012 3976 20040
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 7466 20040 7472 20052
rect 4212 20012 7472 20040
rect 4212 20000 4218 20012
rect 2406 19904 2412 19916
rect 1688 19876 2412 19904
rect 1688 19845 1716 19876
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 3234 19904 3240 19916
rect 3147 19876 3240 19904
rect 3234 19864 3240 19876
rect 3292 19904 3298 19916
rect 4632 19904 4660 20012
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 7650 20040 7656 20052
rect 7607 20012 7656 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 7098 19972 7104 19984
rect 7059 19944 7104 19972
rect 7098 19932 7104 19944
rect 7156 19932 7162 19984
rect 5149 19907 5207 19913
rect 5149 19904 5161 19907
rect 3292 19876 4200 19904
rect 3292 19864 3298 19876
rect 4172 19848 4200 19876
rect 4540 19876 4660 19904
rect 4816 19876 5161 19904
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1673 19799 1731 19805
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3694 19836 3700 19848
rect 3191 19808 3700 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 4154 19836 4160 19848
rect 4115 19808 4160 19836
rect 4154 19796 4160 19808
rect 4212 19796 4218 19848
rect 4540 19845 4568 19876
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19805 4583 19839
rect 4525 19799 4583 19805
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 4816 19836 4844 19876
rect 5149 19873 5161 19876
rect 5195 19873 5207 19907
rect 7576 19904 7604 20003
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 14461 20043 14519 20049
rect 14461 20009 14473 20043
rect 14507 20040 14519 20043
rect 15654 20040 15660 20052
rect 14507 20012 15660 20040
rect 14507 20009 14519 20012
rect 14461 20003 14519 20009
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 18785 20043 18843 20049
rect 18785 20009 18797 20043
rect 18831 20040 18843 20043
rect 19242 20040 19248 20052
rect 18831 20012 19248 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 19242 20000 19248 20012
rect 19300 20000 19306 20052
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19518 20040 19524 20052
rect 19392 20012 19524 20040
rect 19392 20000 19398 20012
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 20070 20040 20076 20052
rect 20031 20012 20076 20040
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 7742 19972 7748 19984
rect 7703 19944 7748 19972
rect 7742 19932 7748 19944
rect 7800 19932 7806 19984
rect 9125 19975 9183 19981
rect 9125 19941 9137 19975
rect 9171 19941 9183 19975
rect 9125 19935 9183 19941
rect 13633 19975 13691 19981
rect 13633 19941 13645 19975
rect 13679 19972 13691 19975
rect 14734 19972 14740 19984
rect 13679 19944 14740 19972
rect 13679 19941 13691 19944
rect 13633 19935 13691 19941
rect 9140 19904 9168 19935
rect 14734 19932 14740 19944
rect 14792 19932 14798 19984
rect 14826 19932 14832 19984
rect 14884 19972 14890 19984
rect 21358 19972 21364 19984
rect 14884 19944 21364 19972
rect 14884 19932 14890 19944
rect 21358 19932 21364 19944
rect 21416 19932 21422 19984
rect 32306 19972 32312 19984
rect 32267 19944 32312 19972
rect 32306 19932 32312 19944
rect 32364 19932 32370 19984
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 5149 19867 5207 19873
rect 6932 19876 7604 19904
rect 8312 19876 9168 19904
rect 9416 19876 10517 19904
rect 4663 19808 4844 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 5350 19796 5356 19848
rect 5408 19836 5414 19848
rect 6932 19845 6960 19876
rect 6825 19839 6883 19845
rect 5408 19808 6684 19836
rect 5408 19796 5414 19808
rect 1765 19771 1823 19777
rect 1765 19737 1777 19771
rect 1811 19768 1823 19771
rect 3326 19768 3332 19780
rect 1811 19740 3332 19768
rect 1811 19737 1823 19740
rect 1765 19731 1823 19737
rect 3326 19728 3332 19740
rect 3384 19728 3390 19780
rect 4246 19768 4252 19780
rect 4207 19740 4252 19768
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19737 4399 19771
rect 5074 19768 5080 19780
rect 5035 19740 5080 19768
rect 4341 19731 4399 19737
rect 4356 19700 4384 19731
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 5258 19768 5264 19780
rect 5219 19740 5264 19768
rect 5258 19728 5264 19740
rect 5316 19728 5322 19780
rect 6546 19700 6552 19712
rect 4356 19672 6552 19700
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 6656 19700 6684 19808
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7374 19836 7380 19848
rect 7147 19808 7380 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 6840 19768 6868 19799
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 8018 19836 8024 19848
rect 7931 19808 8024 19836
rect 8018 19796 8024 19808
rect 8076 19836 8082 19848
rect 8312 19836 8340 19876
rect 8076 19808 8340 19836
rect 8076 19796 8082 19808
rect 8478 19796 8484 19848
rect 8536 19836 8542 19848
rect 9416 19845 9444 19876
rect 10505 19873 10517 19876
rect 10551 19873 10563 19907
rect 10962 19904 10968 19916
rect 10505 19867 10563 19873
rect 10796 19876 10968 19904
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8536 19808 9413 19836
rect 8536 19796 8542 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9950 19796 9956 19848
rect 10008 19836 10014 19848
rect 10318 19836 10324 19848
rect 10008 19808 10324 19836
rect 10008 19796 10014 19808
rect 10318 19796 10324 19808
rect 10376 19836 10382 19848
rect 10796 19845 10824 19876
rect 10962 19864 10968 19876
rect 11020 19904 11026 19916
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 11020 19876 11897 19904
rect 11020 19864 11026 19876
rect 11885 19873 11897 19876
rect 11931 19873 11943 19907
rect 19334 19904 19340 19916
rect 11885 19867 11943 19873
rect 15120 19876 19340 19904
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 10376 19808 10425 19836
rect 10376 19796 10382 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11103 19808 11713 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 7282 19768 7288 19780
rect 6840 19740 7288 19768
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 9125 19771 9183 19777
rect 9125 19768 9137 19771
rect 8996 19740 9137 19768
rect 8996 19728 9002 19740
rect 9125 19737 9137 19740
rect 9171 19737 9183 19771
rect 9125 19731 9183 19737
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 9766 19768 9772 19780
rect 9355 19740 9772 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 9766 19728 9772 19740
rect 9824 19768 9830 19780
rect 10226 19768 10232 19780
rect 9824 19740 10232 19768
rect 9824 19728 9830 19740
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 10686 19728 10692 19780
rect 10744 19768 10750 19780
rect 11072 19768 11100 19799
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 13354 19836 13360 19848
rect 12768 19808 13360 19836
rect 12768 19796 12774 19808
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13504 19808 13553 19836
rect 13504 19796 13510 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 14366 19836 14372 19848
rect 14327 19808 14372 19836
rect 13541 19799 13599 19805
rect 14366 19796 14372 19808
rect 14424 19796 14430 19848
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 15120 19845 15148 19876
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 20622 19904 20628 19916
rect 19720 19876 20628 19904
rect 15105 19839 15163 19845
rect 15105 19836 15117 19839
rect 14608 19808 15117 19836
rect 14608 19796 14614 19808
rect 15105 19805 15117 19808
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 16301 19839 16359 19845
rect 16301 19836 16313 19839
rect 15896 19808 16313 19836
rect 15896 19796 15902 19808
rect 16301 19805 16313 19808
rect 16347 19836 16359 19839
rect 18509 19839 18567 19845
rect 18509 19836 18521 19839
rect 16347 19808 18521 19836
rect 16347 19805 16359 19808
rect 16301 19799 16359 19805
rect 18509 19805 18521 19808
rect 18555 19805 18567 19839
rect 18509 19799 18567 19805
rect 19429 19839 19487 19845
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 15654 19768 15660 19780
rect 10744 19740 11100 19768
rect 15615 19740 15660 19768
rect 10744 19728 10750 19740
rect 15654 19728 15660 19740
rect 15712 19728 15718 19780
rect 16853 19771 16911 19777
rect 16853 19737 16865 19771
rect 16899 19768 16911 19771
rect 17126 19768 17132 19780
rect 16899 19740 17132 19768
rect 16899 19737 16911 19740
rect 16853 19731 16911 19737
rect 17126 19728 17132 19740
rect 17184 19728 17190 19780
rect 7834 19700 7840 19712
rect 6656 19672 7840 19700
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 11514 19700 11520 19712
rect 11475 19672 11520 19700
rect 11514 19660 11520 19672
rect 11572 19660 11578 19712
rect 19444 19700 19472 19799
rect 19518 19796 19524 19848
rect 19576 19836 19582 19848
rect 19720 19845 19748 19876
rect 20180 19848 20208 19876
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 22557 19907 22615 19913
rect 22557 19873 22569 19907
rect 22603 19904 22615 19907
rect 23198 19904 23204 19916
rect 22603 19876 23204 19904
rect 22603 19873 22615 19876
rect 22557 19867 22615 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 32490 19904 32496 19916
rect 32140 19876 32496 19904
rect 19705 19839 19763 19845
rect 19576 19808 19621 19836
rect 19576 19796 19582 19808
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19894 19839 19952 19845
rect 19894 19805 19906 19839
rect 19940 19836 19952 19839
rect 19940 19805 19978 19836
rect 19894 19799 19978 19805
rect 19610 19728 19616 19780
rect 19668 19768 19674 19780
rect 19797 19771 19855 19777
rect 19797 19768 19809 19771
rect 19668 19740 19809 19768
rect 19668 19728 19674 19740
rect 19797 19737 19809 19740
rect 19843 19737 19855 19771
rect 19950 19768 19978 19799
rect 20162 19796 20168 19848
rect 20220 19796 20226 19848
rect 21082 19836 21088 19848
rect 20272 19808 21088 19836
rect 20070 19768 20076 19780
rect 19950 19740 20076 19768
rect 19797 19731 19855 19737
rect 20070 19728 20076 19740
rect 20128 19768 20134 19780
rect 20272 19768 20300 19808
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 31938 19836 31944 19848
rect 31899 19808 31944 19836
rect 31938 19796 31944 19808
rect 31996 19796 32002 19848
rect 32140 19845 32168 19876
rect 32490 19864 32496 19876
rect 32548 19864 32554 19916
rect 32125 19839 32183 19845
rect 32125 19805 32137 19839
rect 32171 19805 32183 19839
rect 32125 19799 32183 19805
rect 32214 19796 32220 19848
rect 32272 19836 32278 19848
rect 32401 19839 32459 19845
rect 32401 19836 32413 19839
rect 32272 19808 32413 19836
rect 32272 19796 32278 19808
rect 32401 19805 32413 19808
rect 32447 19805 32459 19839
rect 32401 19799 32459 19805
rect 32585 19839 32643 19845
rect 32585 19805 32597 19839
rect 32631 19805 32643 19839
rect 32585 19799 32643 19805
rect 20806 19768 20812 19780
rect 20128 19740 20300 19768
rect 20767 19740 20812 19768
rect 20128 19728 20134 19740
rect 20806 19728 20812 19740
rect 20864 19768 20870 19780
rect 21726 19768 21732 19780
rect 20864 19740 21732 19768
rect 20864 19728 20870 19740
rect 21726 19728 21732 19740
rect 21784 19728 21790 19780
rect 32600 19768 32628 19799
rect 32416 19740 32628 19768
rect 32416 19712 32444 19740
rect 19886 19700 19892 19712
rect 19444 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 32398 19660 32404 19712
rect 32456 19660 32462 19712
rect 1104 19610 35027 19632
rect 1104 19558 9390 19610
rect 9442 19558 9454 19610
rect 9506 19558 9518 19610
rect 9570 19558 9582 19610
rect 9634 19558 9646 19610
rect 9698 19558 17831 19610
rect 17883 19558 17895 19610
rect 17947 19558 17959 19610
rect 18011 19558 18023 19610
rect 18075 19558 18087 19610
rect 18139 19558 26272 19610
rect 26324 19558 26336 19610
rect 26388 19558 26400 19610
rect 26452 19558 26464 19610
rect 26516 19558 26528 19610
rect 26580 19558 34713 19610
rect 34765 19558 34777 19610
rect 34829 19558 34841 19610
rect 34893 19558 34905 19610
rect 34957 19558 34969 19610
rect 35021 19558 35027 19610
rect 1104 19536 35027 19558
rect 1854 19456 1860 19508
rect 1912 19496 1918 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 1912 19468 4445 19496
rect 1912 19456 1918 19468
rect 4433 19465 4445 19468
rect 4479 19496 4491 19499
rect 4522 19496 4528 19508
rect 4479 19468 4528 19496
rect 4479 19465 4491 19468
rect 4433 19459 4491 19465
rect 4522 19456 4528 19468
rect 4580 19496 4586 19508
rect 5074 19496 5080 19508
rect 4580 19468 5080 19496
rect 4580 19456 4586 19468
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 17221 19499 17279 19505
rect 17221 19496 17233 19499
rect 16347 19468 17233 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 17221 19465 17233 19468
rect 17267 19496 17279 19499
rect 19518 19496 19524 19508
rect 17267 19468 19524 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 19794 19456 19800 19508
rect 19852 19496 19858 19508
rect 20349 19499 20407 19505
rect 20349 19496 20361 19499
rect 19852 19468 20361 19496
rect 19852 19456 19858 19468
rect 20349 19465 20361 19468
rect 20395 19465 20407 19499
rect 29178 19496 29184 19508
rect 20349 19459 20407 19465
rect 25240 19468 29184 19496
rect 25240 19440 25268 19468
rect 29178 19456 29184 19468
rect 29236 19456 29242 19508
rect 32214 19456 32220 19508
rect 32272 19496 32278 19508
rect 32493 19499 32551 19505
rect 32493 19496 32505 19499
rect 32272 19468 32505 19496
rect 32272 19456 32278 19468
rect 32493 19465 32505 19468
rect 32539 19465 32551 19499
rect 32493 19459 32551 19465
rect 32582 19456 32588 19508
rect 32640 19496 32646 19508
rect 32677 19499 32735 19505
rect 32677 19496 32689 19499
rect 32640 19468 32689 19496
rect 32640 19456 32646 19468
rect 32677 19465 32689 19468
rect 32723 19465 32735 19499
rect 32677 19459 32735 19465
rect 32861 19499 32919 19505
rect 32861 19465 32873 19499
rect 32907 19496 32919 19499
rect 33042 19496 33048 19508
rect 32907 19468 33048 19496
rect 32907 19465 32919 19468
rect 32861 19459 32919 19465
rect 33042 19456 33048 19468
rect 33100 19456 33106 19508
rect 2768 19431 2826 19437
rect 2768 19397 2780 19431
rect 2814 19428 2826 19431
rect 2958 19428 2964 19440
rect 2814 19400 2964 19428
rect 2814 19397 2826 19400
rect 2768 19391 2826 19397
rect 2958 19388 2964 19400
rect 3016 19388 3022 19440
rect 4264 19400 7144 19428
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 3510 19360 3516 19372
rect 2547 19332 3516 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 3510 19320 3516 19332
rect 3568 19360 3574 19372
rect 3878 19360 3884 19372
rect 3568 19332 3884 19360
rect 3568 19320 3574 19332
rect 3878 19320 3884 19332
rect 3936 19360 3942 19372
rect 4264 19360 4292 19400
rect 4614 19360 4620 19372
rect 3936 19332 4292 19360
rect 4575 19332 4620 19360
rect 3936 19320 3942 19332
rect 4614 19320 4620 19332
rect 4672 19360 4678 19372
rect 6638 19360 6644 19372
rect 4672 19332 6644 19360
rect 4672 19320 4678 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 7116 19369 7144 19400
rect 16022 19388 16028 19440
rect 16080 19428 16086 19440
rect 19426 19428 19432 19440
rect 16080 19400 17356 19428
rect 16080 19388 16086 19400
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 7368 19363 7426 19369
rect 7368 19329 7380 19363
rect 7414 19360 7426 19363
rect 7650 19360 7656 19372
rect 7414 19332 7656 19360
rect 7414 19329 7426 19332
rect 7368 19323 7426 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8996 19332 9045 19360
rect 8996 19320 9002 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 9766 19360 9772 19372
rect 9263 19332 9772 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 10778 19360 10784 19372
rect 10739 19332 10784 19360
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12713 19363 12771 19369
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13354 19360 13360 19372
rect 12759 19332 13360 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 15188 19363 15246 19369
rect 15188 19329 15200 19363
rect 15234 19360 15246 19363
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 15234 19332 16865 19360
rect 15234 19329 15246 19332
rect 15188 19323 15246 19329
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19360 17095 19363
rect 17126 19360 17132 19372
rect 17083 19332 17132 19360
rect 17083 19329 17095 19332
rect 17037 19323 17095 19329
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 17328 19369 17356 19400
rect 18984 19400 19432 19428
rect 18984 19369 19012 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 24765 19431 24823 19437
rect 24765 19397 24777 19431
rect 24811 19428 24823 19431
rect 25222 19428 25228 19440
rect 24811 19400 25228 19428
rect 24811 19397 24823 19400
rect 24765 19391 24823 19397
rect 25222 19388 25228 19400
rect 25280 19388 25286 19440
rect 28166 19388 28172 19440
rect 28224 19428 28230 19440
rect 28353 19431 28411 19437
rect 28353 19428 28365 19431
rect 28224 19400 28365 19428
rect 28224 19388 28230 19400
rect 28353 19397 28365 19400
rect 28399 19397 28411 19431
rect 29196 19428 29224 19456
rect 31938 19428 31944 19440
rect 29196 19400 31944 19428
rect 28353 19391 28411 19397
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19225 19363 19283 19369
rect 19225 19360 19237 19363
rect 19116 19332 19237 19360
rect 19116 19320 19122 19332
rect 19225 19329 19237 19332
rect 19271 19329 19283 19363
rect 19225 19323 19283 19329
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 23198 19360 23204 19372
rect 23155 19332 23204 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 23198 19320 23204 19332
rect 23256 19320 23262 19372
rect 27246 19360 27252 19372
rect 27207 19332 27252 19360
rect 27246 19320 27252 19332
rect 27304 19320 27310 19372
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19360 27491 19363
rect 27890 19360 27896 19372
rect 27479 19332 27896 19360
rect 27479 19329 27491 19332
rect 27433 19323 27491 19329
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 28994 19360 29000 19372
rect 28955 19332 29000 19360
rect 28994 19320 29000 19332
rect 29052 19320 29058 19372
rect 29362 19360 29368 19372
rect 29323 19332 29368 19360
rect 29362 19320 29368 19332
rect 29420 19320 29426 19372
rect 31220 19369 31248 19400
rect 31938 19388 31944 19400
rect 31996 19428 32002 19440
rect 32309 19431 32367 19437
rect 32309 19428 32321 19431
rect 31996 19400 32321 19428
rect 31996 19388 32002 19400
rect 32309 19397 32321 19400
rect 32355 19397 32367 19431
rect 32309 19391 32367 19397
rect 31205 19363 31263 19369
rect 31205 19329 31217 19363
rect 31251 19329 31263 19363
rect 31386 19360 31392 19372
rect 31347 19332 31392 19360
rect 31205 19323 31263 19329
rect 31386 19320 31392 19332
rect 31444 19320 31450 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 32585 19363 32643 19369
rect 32585 19360 32597 19363
rect 32456 19332 32597 19360
rect 32456 19320 32462 19332
rect 32585 19329 32597 19332
rect 32631 19329 32643 19363
rect 32585 19323 32643 19329
rect 4801 19295 4859 19301
rect 4801 19261 4813 19295
rect 4847 19261 4859 19295
rect 4801 19255 4859 19261
rect 10505 19295 10563 19301
rect 10505 19261 10517 19295
rect 10551 19292 10563 19295
rect 11054 19292 11060 19304
rect 10551 19264 11060 19292
rect 10551 19261 10563 19264
rect 10505 19255 10563 19261
rect 3881 19159 3939 19165
rect 3881 19125 3893 19159
rect 3927 19156 3939 19159
rect 4246 19156 4252 19168
rect 3927 19128 4252 19156
rect 3927 19125 3939 19128
rect 3881 19119 3939 19125
rect 4246 19116 4252 19128
rect 4304 19156 4310 19168
rect 4816 19156 4844 19255
rect 11054 19252 11060 19264
rect 11112 19292 11118 19304
rect 11514 19292 11520 19304
rect 11112 19264 11520 19292
rect 11112 19252 11118 19264
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14792 19264 14933 19292
rect 14792 19252 14798 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 23382 19292 23388 19304
rect 23343 19264 23388 19292
rect 14921 19255 14979 19261
rect 23382 19252 23388 19264
rect 23440 19252 23446 19304
rect 28534 19252 28540 19304
rect 28592 19292 28598 19304
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28592 19264 28825 19292
rect 28592 19252 28598 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 29270 19292 29276 19304
rect 29231 19264 29276 19292
rect 28813 19255 28871 19261
rect 29270 19252 29276 19264
rect 29328 19292 29334 19304
rect 31113 19295 31171 19301
rect 31113 19292 31125 19295
rect 29328 19264 31125 19292
rect 29328 19252 29334 19264
rect 31113 19261 31125 19264
rect 31159 19261 31171 19295
rect 31113 19255 31171 19261
rect 10134 19224 10140 19236
rect 8036 19196 10140 19224
rect 8036 19156 8064 19196
rect 10134 19184 10140 19196
rect 10192 19184 10198 19236
rect 31128 19224 31156 19255
rect 32674 19224 32680 19236
rect 31128 19196 32680 19224
rect 32674 19184 32680 19196
rect 32732 19184 32738 19236
rect 4304 19128 8064 19156
rect 4304 19116 4310 19128
rect 8110 19116 8116 19168
rect 8168 19156 8174 19168
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 8168 19128 8493 19156
rect 8168 19116 8174 19128
rect 8481 19125 8493 19128
rect 8527 19125 8539 19159
rect 9122 19156 9128 19168
rect 9083 19128 9128 19156
rect 8481 19119 8539 19125
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 10226 19156 10232 19168
rect 10187 19128 10232 19156
rect 10226 19116 10232 19128
rect 10284 19116 10290 19168
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 20990 19156 20996 19168
rect 19208 19128 20996 19156
rect 19208 19116 19214 19128
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 27338 19156 27344 19168
rect 27299 19128 27344 19156
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 1104 19066 34868 19088
rect 1104 19014 5170 19066
rect 5222 19014 5234 19066
rect 5286 19014 5298 19066
rect 5350 19014 5362 19066
rect 5414 19014 5426 19066
rect 5478 19014 13611 19066
rect 13663 19014 13675 19066
rect 13727 19014 13739 19066
rect 13791 19014 13803 19066
rect 13855 19014 13867 19066
rect 13919 19014 22052 19066
rect 22104 19014 22116 19066
rect 22168 19014 22180 19066
rect 22232 19014 22244 19066
rect 22296 19014 22308 19066
rect 22360 19014 30493 19066
rect 30545 19014 30557 19066
rect 30609 19014 30621 19066
rect 30673 19014 30685 19066
rect 30737 19014 30749 19066
rect 30801 19014 34868 19066
rect 1104 18992 34868 19014
rect 7650 18952 7656 18964
rect 7611 18924 7656 18952
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 14553 18955 14611 18961
rect 14553 18921 14565 18955
rect 14599 18952 14611 18955
rect 14642 18952 14648 18964
rect 14599 18924 14648 18952
rect 14599 18921 14611 18924
rect 14553 18915 14611 18921
rect 14642 18912 14648 18924
rect 14700 18952 14706 18964
rect 16666 18952 16672 18964
rect 14700 18924 16252 18952
rect 16627 18924 16672 18952
rect 14700 18912 14706 18924
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3145 18887 3203 18893
rect 3145 18884 3157 18887
rect 3016 18856 3157 18884
rect 3016 18844 3022 18856
rect 3145 18853 3157 18856
rect 3191 18853 3203 18887
rect 8478 18884 8484 18896
rect 3145 18847 3203 18853
rect 7944 18856 8484 18884
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7944 18825 7972 18856
rect 8478 18844 8484 18856
rect 8536 18844 8542 18896
rect 16224 18884 16252 18924
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 18693 18955 18751 18961
rect 18693 18921 18705 18955
rect 18739 18952 18751 18955
rect 19334 18952 19340 18964
rect 18739 18924 19340 18952
rect 18739 18921 18751 18924
rect 18693 18915 18751 18921
rect 18708 18884 18736 18915
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 19610 18912 19616 18964
rect 19668 18952 19674 18964
rect 20809 18955 20867 18961
rect 20809 18952 20821 18955
rect 19668 18924 20821 18952
rect 19668 18912 19674 18924
rect 20809 18921 20821 18924
rect 20855 18921 20867 18955
rect 25866 18952 25872 18964
rect 25827 18924 25872 18952
rect 20809 18915 20867 18921
rect 25866 18912 25872 18924
rect 25924 18912 25930 18964
rect 33137 18955 33195 18961
rect 33137 18921 33149 18955
rect 33183 18952 33195 18955
rect 33318 18952 33324 18964
rect 33183 18924 33324 18952
rect 33183 18921 33195 18924
rect 33137 18915 33195 18921
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 27706 18884 27712 18896
rect 16224 18856 18736 18884
rect 26068 18856 27712 18884
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 7156 18788 7849 18816
rect 7156 18776 7162 18788
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 7929 18819 7987 18825
rect 7929 18785 7941 18819
rect 7975 18785 7987 18819
rect 7929 18779 7987 18785
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 9122 18816 9128 18828
rect 8251 18788 9128 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 9122 18776 9128 18788
rect 9180 18776 9186 18828
rect 26068 18825 26096 18856
rect 27706 18844 27712 18856
rect 27764 18844 27770 18896
rect 32766 18844 32772 18896
rect 32824 18844 32830 18896
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18816 12403 18819
rect 26053 18819 26111 18825
rect 12391 18788 15424 18816
rect 12391 18785 12403 18788
rect 12345 18779 12403 18785
rect 15396 18760 15424 18788
rect 26053 18785 26065 18819
rect 26099 18785 26111 18819
rect 26053 18779 26111 18785
rect 26145 18819 26203 18825
rect 26145 18785 26157 18819
rect 26191 18816 26203 18819
rect 27338 18816 27344 18828
rect 26191 18788 27344 18816
rect 26191 18785 26203 18788
rect 26145 18779 26203 18785
rect 27338 18776 27344 18788
rect 27396 18776 27402 18828
rect 31849 18819 31907 18825
rect 31849 18785 31861 18819
rect 31895 18816 31907 18819
rect 32398 18816 32404 18828
rect 31895 18788 32404 18816
rect 31895 18785 31907 18788
rect 31849 18779 31907 18785
rect 32398 18776 32404 18788
rect 32456 18776 32462 18828
rect 32784 18816 32812 18844
rect 32784 18788 32996 18816
rect 3326 18748 3332 18760
rect 3287 18720 3332 18748
rect 3326 18708 3332 18720
rect 3384 18708 3390 18760
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 8297 18751 8355 18757
rect 3476 18720 3521 18748
rect 3476 18708 3482 18720
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 10226 18748 10232 18760
rect 8343 18720 10232 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18717 10471 18751
rect 10413 18711 10471 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10686 18748 10692 18760
rect 10551 18720 10692 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 3234 18680 3240 18692
rect 3191 18652 3240 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3234 18640 3240 18652
rect 3292 18680 3298 18692
rect 7190 18680 7196 18692
rect 3292 18652 7196 18680
rect 3292 18640 3298 18652
rect 7190 18640 7196 18652
rect 7248 18680 7254 18692
rect 7248 18652 8064 18680
rect 7248 18640 7254 18652
rect 8036 18621 8064 18652
rect 8110 18640 8116 18692
rect 8168 18680 8174 18692
rect 10428 18680 10456 18711
rect 10686 18708 10692 18720
rect 10744 18748 10750 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 10744 18720 11989 18748
rect 10744 18708 10750 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12434 18748 12440 18760
rect 12299 18720 12440 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14792 18720 15301 18748
rect 14792 18708 14798 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15378 18708 15384 18760
rect 15436 18708 15442 18760
rect 19426 18748 19432 18760
rect 19387 18720 19432 18748
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 20898 18748 20904 18760
rect 19628 18720 20904 18748
rect 8168 18652 10456 18680
rect 8168 18640 8174 18652
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 12400 18652 14381 18680
rect 12400 18640 12406 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14553 18683 14611 18689
rect 14553 18649 14565 18683
rect 14599 18680 14611 18683
rect 15556 18683 15614 18689
rect 14599 18652 15516 18680
rect 14599 18649 14611 18652
rect 14553 18643 14611 18649
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 14737 18615 14795 18621
rect 14737 18581 14749 18615
rect 14783 18612 14795 18615
rect 15194 18612 15200 18624
rect 14783 18584 15200 18612
rect 14783 18581 14795 18584
rect 14737 18575 14795 18581
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 15488 18612 15516 18652
rect 15556 18649 15568 18683
rect 15602 18680 15614 18683
rect 15746 18680 15752 18692
rect 15602 18652 15752 18680
rect 15602 18649 15614 18652
rect 15556 18643 15614 18649
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 18877 18683 18935 18689
rect 18877 18649 18889 18683
rect 18923 18680 18935 18683
rect 19334 18680 19340 18692
rect 18923 18652 19340 18680
rect 18923 18649 18935 18652
rect 18877 18643 18935 18649
rect 19334 18640 19340 18652
rect 19392 18680 19398 18692
rect 19628 18680 19656 18720
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23532 18720 23765 18748
rect 23532 18708 23538 18720
rect 23753 18717 23765 18720
rect 23799 18748 23811 18751
rect 23842 18748 23848 18760
rect 23799 18720 23848 18748
rect 23799 18717 23811 18720
rect 23753 18711 23811 18717
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18717 24087 18751
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24029 18711 24087 18717
rect 19702 18689 19708 18692
rect 19392 18652 19656 18680
rect 19392 18640 19398 18652
rect 19696 18643 19708 18689
rect 19760 18680 19766 18692
rect 24044 18680 24072 18711
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25041 18751 25099 18757
rect 25041 18717 25053 18751
rect 25087 18748 25099 18751
rect 25130 18748 25136 18760
rect 25087 18720 25136 18748
rect 25087 18717 25099 18720
rect 25041 18711 25099 18717
rect 25056 18680 25084 18711
rect 25130 18708 25136 18720
rect 25188 18748 25194 18760
rect 25958 18748 25964 18760
rect 25188 18720 25964 18748
rect 25188 18708 25194 18720
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 26234 18748 26240 18760
rect 26195 18720 26240 18748
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26329 18751 26387 18757
rect 26329 18717 26341 18751
rect 26375 18717 26387 18751
rect 26329 18711 26387 18717
rect 19760 18652 19796 18680
rect 24044 18652 25084 18680
rect 19702 18640 19708 18643
rect 19760 18640 19766 18652
rect 25682 18640 25688 18692
rect 25740 18680 25746 18692
rect 26344 18680 26372 18711
rect 27246 18708 27252 18760
rect 27304 18748 27310 18760
rect 27709 18751 27767 18757
rect 27709 18748 27721 18751
rect 27304 18720 27721 18748
rect 27304 18708 27310 18720
rect 27709 18717 27721 18720
rect 27755 18717 27767 18751
rect 27890 18748 27896 18760
rect 27851 18720 27896 18748
rect 27709 18711 27767 18717
rect 27890 18708 27896 18720
rect 27948 18708 27954 18760
rect 28534 18748 28540 18760
rect 28495 18720 28540 18748
rect 28534 18708 28540 18720
rect 28592 18708 28598 18760
rect 28626 18708 28632 18760
rect 28684 18748 28690 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28684 18720 28825 18748
rect 28684 18708 28690 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29270 18748 29276 18760
rect 29043 18720 29276 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 25740 18652 26372 18680
rect 27341 18683 27399 18689
rect 25740 18640 25746 18652
rect 27341 18649 27353 18683
rect 27387 18649 27399 18683
rect 28828 18680 28856 18711
rect 29270 18708 29276 18720
rect 29328 18708 29334 18760
rect 29822 18748 29828 18760
rect 29783 18720 29828 18748
rect 29822 18708 29828 18720
rect 29880 18708 29886 18760
rect 30098 18748 30104 18760
rect 30059 18720 30104 18748
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 32030 18748 32036 18760
rect 31991 18720 32036 18748
rect 32030 18708 32036 18720
rect 32088 18708 32094 18760
rect 32217 18751 32275 18757
rect 32217 18717 32229 18751
rect 32263 18748 32275 18751
rect 32677 18751 32735 18757
rect 32677 18748 32689 18751
rect 32263 18720 32689 18748
rect 32263 18717 32275 18720
rect 32217 18711 32275 18717
rect 32677 18717 32689 18720
rect 32723 18717 32735 18751
rect 32677 18711 32735 18717
rect 32766 18708 32772 18760
rect 32824 18748 32830 18760
rect 32968 18757 32996 18788
rect 32953 18751 33011 18757
rect 32824 18720 32869 18748
rect 32824 18708 32830 18720
rect 32953 18717 32965 18751
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 29362 18680 29368 18692
rect 28828 18652 29368 18680
rect 27341 18643 27399 18649
rect 16942 18612 16948 18624
rect 15488 18584 16948 18612
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 18506 18612 18512 18624
rect 18467 18584 18512 18612
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 18693 18615 18751 18621
rect 18693 18581 18705 18615
rect 18739 18612 18751 18615
rect 19610 18612 19616 18624
rect 18739 18584 19616 18612
rect 18739 18581 18751 18584
rect 18693 18575 18751 18581
rect 19610 18572 19616 18584
rect 19668 18612 19674 18624
rect 20070 18612 20076 18624
rect 19668 18584 20076 18612
rect 19668 18572 19674 18584
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 23566 18612 23572 18624
rect 23527 18584 23572 18612
rect 23566 18572 23572 18584
rect 23624 18572 23630 18624
rect 23937 18615 23995 18621
rect 23937 18581 23949 18615
rect 23983 18612 23995 18615
rect 24394 18612 24400 18624
rect 23983 18584 24400 18612
rect 23983 18581 23995 18584
rect 23937 18575 23995 18581
rect 24394 18572 24400 18584
rect 24452 18572 24458 18624
rect 24578 18612 24584 18624
rect 24539 18584 24584 18612
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 24946 18612 24952 18624
rect 24907 18584 24952 18612
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 27062 18612 27068 18624
rect 26292 18584 27068 18612
rect 26292 18572 26298 18584
rect 27062 18572 27068 18584
rect 27120 18612 27126 18624
rect 27356 18612 27384 18643
rect 29362 18640 29368 18652
rect 29420 18680 29426 18692
rect 29733 18683 29791 18689
rect 29733 18680 29745 18683
rect 29420 18652 29745 18680
rect 29420 18640 29426 18652
rect 29733 18649 29745 18652
rect 29779 18649 29791 18683
rect 29733 18643 29791 18649
rect 28350 18612 28356 18624
rect 27120 18584 27384 18612
rect 28311 18584 28356 18612
rect 27120 18572 27126 18584
rect 28350 18572 28356 18584
rect 28408 18572 28414 18624
rect 1104 18522 35027 18544
rect 1104 18470 9390 18522
rect 9442 18470 9454 18522
rect 9506 18470 9518 18522
rect 9570 18470 9582 18522
rect 9634 18470 9646 18522
rect 9698 18470 17831 18522
rect 17883 18470 17895 18522
rect 17947 18470 17959 18522
rect 18011 18470 18023 18522
rect 18075 18470 18087 18522
rect 18139 18470 26272 18522
rect 26324 18470 26336 18522
rect 26388 18470 26400 18522
rect 26452 18470 26464 18522
rect 26516 18470 26528 18522
rect 26580 18470 34713 18522
rect 34765 18470 34777 18522
rect 34829 18470 34841 18522
rect 34893 18470 34905 18522
rect 34957 18470 34969 18522
rect 35021 18470 35027 18522
rect 1104 18448 35027 18470
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8938 18408 8944 18420
rect 8251 18380 8944 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 15746 18408 15752 18420
rect 12492 18380 15608 18408
rect 15707 18380 15752 18408
rect 12492 18368 12498 18380
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 7098 18340 7104 18352
rect 6871 18312 7104 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 12066 18300 12072 18352
rect 12124 18340 12130 18352
rect 12342 18340 12348 18352
rect 12124 18312 12348 18340
rect 12124 18300 12130 18312
rect 12342 18300 12348 18312
rect 12400 18340 12406 18352
rect 14734 18340 14740 18352
rect 12400 18312 12480 18340
rect 14695 18312 14740 18340
rect 12400 18300 12406 18312
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 6696 18244 8033 18272
rect 6696 18232 6702 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8021 18235 8079 18241
rect 8110 18232 8116 18284
rect 8168 18272 8174 18284
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 8168 18244 8217 18272
rect 8168 18232 8174 18244
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8205 18235 8263 18241
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 11054 18272 11060 18284
rect 10367 18244 11060 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12452 18281 12480 18312
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 15580 18340 15608 18380
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 16117 18411 16175 18417
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 16666 18408 16672 18420
rect 16163 18380 16672 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 24765 18411 24823 18417
rect 24765 18377 24777 18411
rect 24811 18408 24823 18411
rect 24946 18408 24952 18420
rect 24811 18380 24952 18408
rect 24811 18377 24823 18380
rect 24765 18371 24823 18377
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 25682 18408 25688 18420
rect 25643 18380 25688 18408
rect 25682 18368 25688 18380
rect 25740 18368 25746 18420
rect 29086 18408 29092 18420
rect 28736 18380 29092 18408
rect 16022 18340 16028 18352
rect 15580 18312 16028 18340
rect 16022 18300 16028 18312
rect 16080 18340 16086 18352
rect 16080 18312 16252 18340
rect 16080 18300 16086 18312
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 11848 18244 12265 18272
rect 11848 18232 11854 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12437 18235 12495 18241
rect 6730 18204 6736 18216
rect 6691 18176 6736 18204
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 6914 18204 6920 18216
rect 6875 18176 6920 18204
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 12158 18204 12164 18216
rect 12119 18176 12164 18204
rect 12158 18164 12164 18176
rect 12216 18164 12222 18216
rect 7282 18136 7288 18148
rect 7243 18108 7288 18136
rect 7282 18096 7288 18108
rect 7340 18096 7346 18148
rect 12268 18136 12296 18235
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 16224 18281 16252 18312
rect 18506 18300 18512 18352
rect 18564 18340 18570 18352
rect 19245 18343 19303 18349
rect 19245 18340 19257 18343
rect 18564 18312 19257 18340
rect 18564 18300 18570 18312
rect 19245 18309 19257 18312
rect 19291 18309 19303 18343
rect 24964 18340 24992 18368
rect 28736 18340 28764 18380
rect 29086 18368 29092 18380
rect 29144 18368 29150 18420
rect 32490 18408 32496 18420
rect 31726 18380 32496 18408
rect 31386 18340 31392 18352
rect 24964 18312 28764 18340
rect 28828 18312 31392 18340
rect 19245 18303 19303 18309
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15712 18244 15945 18272
rect 15712 18232 15718 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 16209 18275 16267 18281
rect 16209 18241 16221 18275
rect 16255 18241 16267 18275
rect 16209 18235 16267 18241
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18272 23535 18275
rect 24578 18272 24584 18284
rect 23523 18244 24584 18272
rect 23523 18241 23535 18244
rect 23477 18235 23535 18241
rect 15948 18204 15976 18235
rect 24578 18232 24584 18244
rect 24636 18232 24642 18284
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 25317 18275 25375 18281
rect 25317 18272 25329 18275
rect 24912 18244 25329 18272
rect 24912 18232 24918 18244
rect 25317 18241 25329 18244
rect 25363 18241 25375 18275
rect 25498 18272 25504 18284
rect 25459 18244 25504 18272
rect 25317 18235 25375 18241
rect 25498 18232 25504 18244
rect 25556 18232 25562 18284
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18272 27951 18275
rect 28350 18272 28356 18284
rect 27939 18244 28356 18272
rect 27939 18241 27951 18244
rect 27893 18235 27951 18241
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 28828 18281 28856 18312
rect 31386 18300 31392 18312
rect 31444 18300 31450 18352
rect 28813 18275 28871 18281
rect 28813 18241 28825 18275
rect 28859 18241 28871 18275
rect 28813 18235 28871 18241
rect 29089 18275 29147 18281
rect 29089 18241 29101 18275
rect 29135 18241 29147 18275
rect 29089 18235 29147 18241
rect 20346 18204 20352 18216
rect 15948 18176 20352 18204
rect 20346 18164 20352 18176
rect 20404 18164 20410 18216
rect 23106 18164 23112 18216
rect 23164 18204 23170 18216
rect 23201 18207 23259 18213
rect 23201 18204 23213 18207
rect 23164 18176 23213 18204
rect 23164 18164 23170 18176
rect 23201 18173 23213 18176
rect 23247 18173 23259 18207
rect 23201 18167 23259 18173
rect 23842 18164 23848 18216
rect 23900 18204 23906 18216
rect 23900 18176 25452 18204
rect 23900 18164 23906 18176
rect 12434 18136 12440 18148
rect 12268 18108 12440 18136
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 10226 18068 10232 18080
rect 10187 18040 10232 18068
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 18230 18028 18236 18080
rect 18288 18068 18294 18080
rect 20533 18071 20591 18077
rect 20533 18068 20545 18071
rect 18288 18040 20545 18068
rect 18288 18028 18294 18040
rect 20533 18037 20545 18040
rect 20579 18037 20591 18071
rect 25314 18068 25320 18080
rect 25275 18040 25320 18068
rect 20533 18031 20591 18037
rect 25314 18028 25320 18040
rect 25372 18028 25378 18080
rect 25424 18068 25452 18176
rect 27246 18164 27252 18216
rect 27304 18204 27310 18216
rect 27525 18207 27583 18213
rect 27525 18204 27537 18207
rect 27304 18176 27537 18204
rect 27304 18164 27310 18176
rect 27525 18173 27537 18176
rect 27571 18173 27583 18207
rect 27525 18167 27583 18173
rect 27985 18207 28043 18213
rect 27985 18173 27997 18207
rect 28031 18204 28043 18207
rect 28994 18204 29000 18216
rect 28031 18176 29000 18204
rect 28031 18173 28043 18176
rect 27985 18167 28043 18173
rect 28994 18164 29000 18176
rect 29052 18164 29058 18216
rect 29104 18204 29132 18235
rect 29178 18232 29184 18284
rect 29236 18272 29242 18284
rect 29365 18275 29423 18281
rect 29365 18272 29377 18275
rect 29236 18244 29377 18272
rect 29236 18232 29242 18244
rect 29365 18241 29377 18244
rect 29411 18241 29423 18275
rect 29730 18272 29736 18284
rect 29691 18244 29736 18272
rect 29365 18235 29423 18241
rect 29730 18232 29736 18244
rect 29788 18232 29794 18284
rect 30098 18204 30104 18216
rect 29104 18176 30104 18204
rect 30098 18164 30104 18176
rect 30156 18164 30162 18216
rect 28534 18096 28540 18148
rect 28592 18136 28598 18148
rect 28629 18139 28687 18145
rect 28629 18136 28641 18139
rect 28592 18108 28641 18136
rect 28592 18096 28598 18108
rect 28629 18105 28641 18108
rect 28675 18105 28687 18139
rect 28629 18099 28687 18105
rect 31726 18068 31754 18380
rect 32490 18368 32496 18380
rect 32548 18368 32554 18420
rect 32674 18368 32680 18420
rect 32732 18408 32738 18420
rect 32769 18411 32827 18417
rect 32769 18408 32781 18411
rect 32732 18380 32781 18408
rect 32732 18368 32738 18380
rect 32769 18377 32781 18380
rect 32815 18377 32827 18411
rect 32769 18371 32827 18377
rect 32398 18232 32404 18284
rect 32456 18272 32462 18284
rect 32493 18275 32551 18281
rect 32493 18272 32505 18275
rect 32456 18244 32505 18272
rect 32456 18232 32462 18244
rect 32493 18241 32505 18244
rect 32539 18241 32551 18275
rect 32493 18235 32551 18241
rect 32306 18204 32312 18216
rect 32267 18176 32312 18204
rect 32306 18164 32312 18176
rect 32364 18164 32370 18216
rect 32858 18204 32864 18216
rect 32819 18176 32864 18204
rect 32858 18164 32864 18176
rect 32916 18164 32922 18216
rect 34330 18204 34336 18216
rect 34291 18176 34336 18204
rect 34330 18164 34336 18176
rect 34388 18164 34394 18216
rect 25424 18040 31754 18068
rect 1104 17978 34868 18000
rect 1104 17926 5170 17978
rect 5222 17926 5234 17978
rect 5286 17926 5298 17978
rect 5350 17926 5362 17978
rect 5414 17926 5426 17978
rect 5478 17926 13611 17978
rect 13663 17926 13675 17978
rect 13727 17926 13739 17978
rect 13791 17926 13803 17978
rect 13855 17926 13867 17978
rect 13919 17926 22052 17978
rect 22104 17926 22116 17978
rect 22168 17926 22180 17978
rect 22232 17926 22244 17978
rect 22296 17926 22308 17978
rect 22360 17926 30493 17978
rect 30545 17926 30557 17978
rect 30609 17926 30621 17978
rect 30673 17926 30685 17978
rect 30737 17926 30749 17978
rect 30801 17926 34868 17978
rect 1104 17904 34868 17926
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17864 6515 17867
rect 6730 17864 6736 17876
rect 6503 17836 6736 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 27982 17864 27988 17876
rect 15436 17836 20484 17864
rect 27943 17836 27988 17864
rect 15436 17824 15442 17836
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 3510 17796 3516 17808
rect 3467 17768 3516 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3510 17756 3516 17768
rect 3568 17756 3574 17808
rect 11514 17688 11520 17740
rect 11572 17728 11578 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 11572 17700 13093 17728
rect 11572 17688 11578 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 18708 17700 19564 17728
rect 3234 17660 3240 17672
rect 3195 17632 3240 17660
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 6362 17660 6368 17672
rect 6323 17632 6368 17660
rect 6362 17620 6368 17632
rect 6420 17620 6426 17672
rect 6546 17660 6552 17672
rect 6507 17632 6552 17660
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 15194 17660 15200 17672
rect 15155 17632 15200 17660
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 18708 17669 18736 17700
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 17552 17632 17601 17660
rect 17552 17620 17558 17632
rect 17589 17629 17601 17632
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 17865 17663 17923 17669
rect 17865 17629 17877 17663
rect 17911 17660 17923 17663
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 17911 17632 18429 17660
rect 17911 17629 17923 17632
rect 17865 17623 17923 17629
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 2869 17595 2927 17601
rect 2869 17592 2881 17595
rect 2740 17564 2881 17592
rect 2740 17552 2746 17564
rect 2869 17561 2881 17564
rect 2915 17561 2927 17595
rect 2869 17555 2927 17561
rect 12158 17552 12164 17604
rect 12216 17552 12222 17604
rect 12805 17595 12863 17601
rect 12805 17561 12817 17595
rect 12851 17592 12863 17595
rect 12894 17592 12900 17604
rect 12851 17564 12900 17592
rect 12851 17561 12863 17564
rect 12805 17555 12863 17561
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 17310 17552 17316 17604
rect 17368 17592 17374 17604
rect 17880 17592 17908 17623
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19300 17632 19441 17660
rect 19300 17620 19306 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19536 17660 19564 17700
rect 20456 17660 20484 17836
rect 27982 17824 27988 17836
rect 28040 17824 28046 17876
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 32677 17867 32735 17873
rect 32677 17864 32689 17867
rect 29052 17836 32689 17864
rect 29052 17824 29058 17836
rect 32677 17833 32689 17836
rect 32723 17833 32735 17867
rect 32677 17827 32735 17833
rect 21542 17796 21548 17808
rect 21503 17768 21548 17796
rect 21542 17756 21548 17768
rect 21600 17796 21606 17808
rect 24762 17796 24768 17808
rect 21600 17768 24768 17796
rect 21600 17756 21606 17768
rect 24762 17756 24768 17768
rect 24820 17756 24826 17808
rect 27617 17731 27675 17737
rect 27617 17697 27629 17731
rect 27663 17728 27675 17731
rect 27890 17728 27896 17740
rect 27663 17700 27896 17728
rect 27663 17697 27675 17700
rect 27617 17691 27675 17697
rect 27890 17688 27896 17700
rect 27948 17728 27954 17740
rect 28445 17731 28503 17737
rect 28445 17728 28457 17731
rect 27948 17700 28457 17728
rect 27948 17688 27954 17700
rect 28445 17697 28457 17700
rect 28491 17697 28503 17731
rect 32306 17728 32312 17740
rect 28445 17691 28503 17697
rect 31772 17700 32312 17728
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 19536 17632 20392 17660
rect 20456 17632 21373 17660
rect 19429 17623 19487 17629
rect 17368 17564 17908 17592
rect 18877 17595 18935 17601
rect 17368 17552 17374 17564
rect 18877 17561 18889 17595
rect 18923 17592 18935 17595
rect 19674 17595 19732 17601
rect 19674 17592 19686 17595
rect 18923 17564 19686 17592
rect 18923 17561 18935 17564
rect 18877 17555 18935 17561
rect 19674 17561 19686 17564
rect 19720 17561 19732 17595
rect 20364 17592 20392 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 21361 17623 21419 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25041 17663 25099 17669
rect 25041 17629 25053 17663
rect 25087 17629 25099 17663
rect 25041 17623 25099 17629
rect 21542 17592 21548 17604
rect 20364 17564 21548 17592
rect 19674 17555 19732 17561
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 25056 17592 25084 17623
rect 25682 17620 25688 17672
rect 25740 17660 25746 17672
rect 27525 17663 27583 17669
rect 27525 17660 27537 17663
rect 25740 17632 27537 17660
rect 25740 17620 25746 17632
rect 27525 17629 27537 17632
rect 27571 17629 27583 17663
rect 27706 17660 27712 17672
rect 27667 17632 27712 17660
rect 27525 17623 27583 17629
rect 27706 17620 27712 17632
rect 27764 17620 27770 17672
rect 27798 17620 27804 17672
rect 27856 17660 27862 17672
rect 27856 17632 27901 17660
rect 27856 17620 27862 17632
rect 28534 17620 28540 17672
rect 28592 17660 28598 17672
rect 28629 17663 28687 17669
rect 28629 17660 28641 17663
rect 28592 17632 28641 17660
rect 28592 17620 28598 17632
rect 28629 17629 28641 17632
rect 28675 17629 28687 17663
rect 28902 17660 28908 17672
rect 28815 17632 28908 17660
rect 28629 17623 28687 17629
rect 28902 17620 28908 17632
rect 28960 17660 28966 17672
rect 30745 17663 30803 17669
rect 30745 17660 30757 17663
rect 28960 17632 30757 17660
rect 28960 17620 28966 17632
rect 30745 17629 30757 17632
rect 30791 17629 30803 17663
rect 30926 17660 30932 17672
rect 30839 17632 30932 17660
rect 30745 17623 30803 17629
rect 30926 17620 30932 17632
rect 30984 17660 30990 17672
rect 31772 17669 31800 17700
rect 32306 17688 32312 17700
rect 32364 17728 32370 17740
rect 33597 17731 33655 17737
rect 33597 17728 33609 17731
rect 32364 17700 33609 17728
rect 32364 17688 32370 17700
rect 33597 17697 33609 17700
rect 33643 17697 33655 17731
rect 33597 17691 33655 17697
rect 31757 17663 31815 17669
rect 31757 17660 31769 17663
rect 30984 17632 31769 17660
rect 30984 17620 30990 17632
rect 31757 17629 31769 17632
rect 31803 17629 31815 17663
rect 31757 17623 31815 17629
rect 31941 17663 31999 17669
rect 31941 17629 31953 17663
rect 31987 17660 31999 17663
rect 32585 17663 32643 17669
rect 31987 17632 32536 17660
rect 31987 17629 31999 17632
rect 31941 17623 31999 17629
rect 26602 17592 26608 17604
rect 25056 17564 26608 17592
rect 26602 17552 26608 17564
rect 26660 17552 26666 17604
rect 31110 17592 31116 17604
rect 31071 17564 31116 17592
rect 31110 17552 31116 17564
rect 31168 17552 31174 17604
rect 31849 17595 31907 17601
rect 31849 17561 31861 17595
rect 31895 17592 31907 17595
rect 32401 17595 32459 17601
rect 32401 17592 32413 17595
rect 31895 17564 32413 17592
rect 31895 17561 31907 17564
rect 31849 17555 31907 17561
rect 32401 17561 32413 17564
rect 32447 17561 32459 17595
rect 32508 17592 32536 17632
rect 32585 17629 32597 17663
rect 32631 17660 32643 17663
rect 32766 17660 32772 17672
rect 32631 17632 32772 17660
rect 32631 17629 32643 17632
rect 32585 17623 32643 17629
rect 32766 17620 32772 17632
rect 32824 17660 32830 17672
rect 33229 17663 33287 17669
rect 33229 17660 33241 17663
rect 32824 17632 33241 17660
rect 32824 17620 32830 17632
rect 33229 17629 33241 17632
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 33413 17663 33471 17669
rect 33413 17629 33425 17663
rect 33459 17629 33471 17663
rect 33413 17623 33471 17629
rect 33428 17592 33456 17623
rect 32508 17564 33456 17592
rect 32401 17555 32459 17561
rect 33244 17536 33272 17564
rect 3050 17524 3056 17536
rect 3011 17496 3056 17524
rect 3050 17484 3056 17496
rect 3108 17484 3114 17536
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 3200 17496 3245 17524
rect 3200 17484 3206 17496
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 9950 17524 9956 17536
rect 7156 17496 9956 17524
rect 7156 17484 7162 17496
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11333 17527 11391 17533
rect 11333 17524 11345 17527
rect 11020 17496 11345 17524
rect 11020 17484 11026 17496
rect 11333 17493 11345 17496
rect 11379 17493 11391 17527
rect 11333 17487 11391 17493
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 13044 17496 16497 17524
rect 13044 17484 13050 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 16485 17487 16543 17493
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 16632 17496 17417 17524
rect 16632 17484 16638 17496
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 17405 17487 17463 17493
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 17773 17527 17831 17533
rect 17773 17524 17785 17527
rect 17644 17496 17785 17524
rect 17644 17484 17650 17496
rect 17773 17493 17785 17496
rect 17819 17493 17831 17527
rect 17773 17487 17831 17493
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 20809 17527 20867 17533
rect 20809 17524 20821 17527
rect 18555 17496 20821 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 20809 17493 20821 17496
rect 20855 17524 20867 17527
rect 20898 17524 20904 17536
rect 20855 17496 20904 17524
rect 20855 17493 20867 17496
rect 20809 17487 20867 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 24581 17527 24639 17533
rect 24581 17493 24593 17527
rect 24627 17524 24639 17527
rect 24854 17524 24860 17536
rect 24627 17496 24860 17524
rect 24627 17493 24639 17496
rect 24581 17487 24639 17493
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 24949 17527 25007 17533
rect 24949 17493 24961 17527
rect 24995 17524 25007 17527
rect 25774 17524 25780 17536
rect 24995 17496 25780 17524
rect 24995 17493 25007 17496
rect 24949 17487 25007 17493
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 28810 17524 28816 17536
rect 28771 17496 28816 17524
rect 28810 17484 28816 17496
rect 28868 17484 28874 17536
rect 33226 17484 33232 17536
rect 33284 17484 33290 17536
rect 1104 17434 35027 17456
rect 1104 17382 9390 17434
rect 9442 17382 9454 17434
rect 9506 17382 9518 17434
rect 9570 17382 9582 17434
rect 9634 17382 9646 17434
rect 9698 17382 17831 17434
rect 17883 17382 17895 17434
rect 17947 17382 17959 17434
rect 18011 17382 18023 17434
rect 18075 17382 18087 17434
rect 18139 17382 26272 17434
rect 26324 17382 26336 17434
rect 26388 17382 26400 17434
rect 26452 17382 26464 17434
rect 26516 17382 26528 17434
rect 26580 17382 34713 17434
rect 34765 17382 34777 17434
rect 34829 17382 34841 17434
rect 34893 17382 34905 17434
rect 34957 17382 34969 17434
rect 35021 17382 35027 17434
rect 1104 17360 35027 17382
rect 4433 17323 4491 17329
rect 4433 17289 4445 17323
rect 4479 17320 4491 17323
rect 6914 17320 6920 17332
rect 4479 17292 6920 17320
rect 4479 17289 4491 17292
rect 4433 17283 4491 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 10318 17320 10324 17332
rect 9600 17292 10324 17320
rect 2958 17252 2964 17264
rect 2919 17224 2964 17252
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 6932 17252 6960 17280
rect 6932 17224 8248 17252
rect 4246 17184 4252 17196
rect 4094 17156 4252 17184
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 6730 17184 6736 17196
rect 6691 17156 6736 17184
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6880 17156 7113 17184
rect 6880 17144 6886 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7524 17156 7573 17184
rect 7524 17144 7530 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8220 17193 8248 17224
rect 9214 17212 9220 17264
rect 9272 17252 9278 17264
rect 9600 17261 9628 17292
rect 10318 17280 10324 17292
rect 10376 17320 10382 17332
rect 14366 17320 14372 17332
rect 10376 17292 14372 17320
rect 10376 17280 10382 17292
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 19484 17292 19533 17320
rect 19484 17280 19490 17292
rect 19521 17289 19533 17292
rect 19567 17289 19579 17323
rect 19521 17283 19579 17289
rect 19628 17292 22094 17320
rect 9585 17255 9643 17261
rect 9585 17252 9597 17255
rect 9272 17224 9597 17252
rect 9272 17212 9278 17224
rect 9585 17221 9597 17224
rect 9631 17221 9643 17255
rect 9585 17215 9643 17221
rect 12250 17212 12256 17264
rect 12308 17212 12314 17264
rect 13170 17212 13176 17264
rect 13228 17252 13234 17264
rect 13265 17255 13323 17261
rect 13265 17252 13277 17255
rect 13228 17224 13277 17252
rect 13228 17212 13234 17224
rect 13265 17221 13277 17224
rect 13311 17221 13323 17255
rect 16850 17252 16856 17264
rect 16811 17224 16856 17252
rect 13265 17215 13323 17221
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 18230 17252 18236 17264
rect 18191 17224 18236 17252
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 9858 17184 9864 17196
rect 9771 17156 9864 17184
rect 8205 17147 8263 17153
rect 9858 17144 9864 17156
rect 9916 17184 9922 17196
rect 10042 17184 10048 17196
rect 9916 17156 10048 17184
rect 9916 17144 9922 17156
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 15436 17156 16221 17184
rect 15436 17144 15442 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 17218 17144 17224 17196
rect 17276 17184 17282 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17276 17156 17693 17184
rect 17276 17144 17282 17156
rect 17681 17153 17693 17156
rect 17727 17184 17739 17187
rect 19628 17184 19656 17292
rect 20809 17255 20867 17261
rect 20809 17221 20821 17255
rect 20855 17252 20867 17255
rect 21174 17252 21180 17264
rect 20855 17224 21180 17252
rect 20855 17221 20867 17224
rect 20809 17215 20867 17221
rect 21174 17212 21180 17224
rect 21232 17212 21238 17264
rect 17727 17156 19656 17184
rect 20625 17187 20683 17193
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17184 20959 17187
rect 20990 17184 20996 17196
rect 20947 17156 20996 17184
rect 20947 17153 20959 17156
rect 20901 17147 20959 17153
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 6638 17116 6644 17128
rect 6599 17088 6644 17116
rect 6638 17076 6644 17088
rect 6696 17076 6702 17128
rect 9769 17119 9827 17125
rect 9769 17085 9781 17119
rect 9815 17116 9827 17119
rect 10134 17116 10140 17128
rect 9815 17088 10140 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 11514 17076 11520 17128
rect 11572 17116 11578 17128
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 11572 17088 13553 17116
rect 11572 17076 11578 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 15930 17116 15936 17128
rect 15891 17088 15936 17116
rect 13541 17079 13599 17085
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 20640 17116 20668 17147
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 22066 17184 22094 17292
rect 23198 17280 23204 17332
rect 23256 17320 23262 17332
rect 25682 17320 25688 17332
rect 23256 17292 25360 17320
rect 25643 17292 25688 17320
rect 23256 17280 23262 17292
rect 23376 17255 23434 17261
rect 23376 17221 23388 17255
rect 23422 17252 23434 17255
rect 23566 17252 23572 17264
rect 23422 17224 23572 17252
rect 23422 17221 23434 17224
rect 23376 17215 23434 17221
rect 23566 17212 23572 17224
rect 23624 17212 23630 17264
rect 23842 17184 23848 17196
rect 22066 17156 23848 17184
rect 23842 17144 23848 17156
rect 23900 17144 23906 17196
rect 25038 17184 25044 17196
rect 24999 17156 25044 17184
rect 25038 17144 25044 17156
rect 25096 17144 25102 17196
rect 25332 17193 25360 17292
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 27798 17280 27804 17332
rect 27856 17320 27862 17332
rect 28537 17323 28595 17329
rect 28537 17320 28549 17323
rect 27856 17292 28549 17320
rect 27856 17280 27862 17292
rect 28537 17289 28549 17292
rect 28583 17289 28595 17323
rect 28537 17283 28595 17289
rect 28810 17280 28816 17332
rect 28868 17280 28874 17332
rect 29086 17280 29092 17332
rect 29144 17320 29150 17332
rect 30745 17323 30803 17329
rect 30745 17320 30757 17323
rect 29144 17292 30757 17320
rect 29144 17280 29150 17292
rect 30745 17289 30757 17292
rect 30791 17289 30803 17323
rect 30926 17320 30932 17332
rect 30887 17292 30932 17320
rect 30745 17283 30803 17289
rect 30926 17280 30932 17292
rect 30984 17280 30990 17332
rect 32214 17320 32220 17332
rect 31496 17292 32220 17320
rect 25409 17255 25467 17261
rect 25409 17221 25421 17255
rect 25455 17252 25467 17255
rect 25774 17252 25780 17264
rect 25455 17224 25780 17252
rect 25455 17221 25467 17224
rect 25409 17215 25467 17221
rect 25774 17212 25780 17224
rect 25832 17212 25838 17264
rect 28629 17255 28687 17261
rect 28629 17221 28641 17255
rect 28675 17252 28687 17255
rect 28828 17252 28856 17280
rect 31496 17261 31524 17292
rect 32214 17280 32220 17292
rect 32272 17320 32278 17332
rect 32509 17323 32567 17329
rect 32509 17320 32521 17323
rect 32272 17292 32521 17320
rect 32272 17280 32278 17292
rect 32509 17289 32521 17292
rect 32555 17289 32567 17323
rect 32509 17283 32567 17289
rect 32677 17323 32735 17329
rect 32677 17289 32689 17323
rect 32723 17320 32735 17323
rect 32858 17320 32864 17332
rect 32723 17292 32864 17320
rect 32723 17289 32735 17292
rect 32677 17283 32735 17289
rect 32858 17280 32864 17292
rect 32916 17280 32922 17332
rect 33226 17320 33232 17332
rect 33187 17292 33232 17320
rect 33226 17280 33232 17292
rect 33284 17280 33290 17332
rect 29825 17255 29883 17261
rect 29825 17252 29837 17255
rect 28675 17224 29837 17252
rect 28675 17221 28687 17224
rect 28629 17215 28687 17221
rect 29825 17221 29837 17224
rect 29871 17221 29883 17255
rect 30837 17255 30895 17261
rect 30837 17252 30849 17255
rect 29825 17215 29883 17221
rect 29932 17224 30849 17252
rect 25590 17193 25596 17196
rect 25134 17187 25192 17193
rect 25134 17153 25146 17187
rect 25180 17153 25192 17187
rect 25134 17147 25192 17153
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 25547 17187 25596 17193
rect 25547 17153 25559 17187
rect 25593 17153 25596 17187
rect 25547 17147 25596 17153
rect 17552 17088 20668 17116
rect 17552 17076 17558 17088
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 23106 17116 23112 17128
rect 22612 17088 23112 17116
rect 22612 17076 22618 17088
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 10152 17048 10180 17076
rect 8168 17020 9720 17048
rect 10152 17020 11928 17048
rect 8168 17008 8174 17020
rect 8202 16980 8208 16992
rect 8163 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 9692 16989 9720 17020
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16949 9735 16983
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 9677 16943 9735 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11204 16952 11805 16980
rect 11204 16940 11210 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11900 16980 11928 17020
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 19518 17048 19524 17060
rect 19300 17020 19524 17048
rect 19300 17008 19306 17020
rect 19518 17008 19524 17020
rect 19576 17008 19582 17060
rect 25148 17048 25176 17147
rect 25590 17144 25596 17147
rect 25648 17144 25654 17196
rect 26050 17144 26056 17196
rect 26108 17184 26114 17196
rect 26145 17187 26203 17193
rect 26145 17184 26157 17187
rect 26108 17156 26157 17184
rect 26108 17144 26114 17156
rect 26145 17153 26157 17156
rect 26191 17153 26203 17187
rect 28534 17184 28540 17196
rect 28495 17156 28540 17184
rect 26145 17147 26203 17153
rect 28534 17144 28540 17156
rect 28592 17144 28598 17196
rect 28813 17187 28871 17193
rect 28813 17153 28825 17187
rect 28859 17184 28871 17187
rect 28902 17184 28908 17196
rect 28859 17156 28908 17184
rect 28859 17153 28871 17156
rect 28813 17147 28871 17153
rect 28902 17144 28908 17156
rect 28960 17144 28966 17196
rect 29932 17193 29960 17224
rect 30837 17221 30849 17224
rect 30883 17252 30895 17255
rect 31481 17255 31539 17261
rect 31481 17252 31493 17255
rect 30883 17224 31493 17252
rect 30883 17221 30895 17224
rect 30837 17215 30895 17221
rect 31481 17221 31493 17224
rect 31527 17221 31539 17255
rect 32309 17255 32367 17261
rect 32309 17252 32321 17255
rect 31481 17215 31539 17221
rect 31680 17224 32321 17252
rect 29733 17187 29791 17193
rect 29733 17153 29745 17187
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17153 29975 17187
rect 29917 17147 29975 17153
rect 30469 17187 30527 17193
rect 30469 17153 30481 17187
rect 30515 17153 30527 17187
rect 30469 17147 30527 17153
rect 30613 17187 30671 17193
rect 30613 17153 30625 17187
rect 30659 17184 30671 17187
rect 31386 17184 31392 17196
rect 30659 17156 31392 17184
rect 30659 17153 30671 17156
rect 30613 17147 30671 17153
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17116 26479 17119
rect 26602 17116 26608 17128
rect 26467 17088 26608 17116
rect 26467 17085 26479 17088
rect 26421 17079 26479 17085
rect 26602 17076 26608 17088
rect 26660 17076 26666 17128
rect 29748 17116 29776 17147
rect 30282 17116 30288 17128
rect 29748 17088 30288 17116
rect 30282 17076 30288 17088
rect 30340 17116 30346 17128
rect 30484 17116 30512 17147
rect 31386 17144 31392 17156
rect 31444 17144 31450 17196
rect 31570 17144 31576 17196
rect 31628 17184 31634 17196
rect 31680 17193 31708 17224
rect 32309 17221 32321 17224
rect 32355 17221 32367 17255
rect 32309 17215 32367 17221
rect 31665 17187 31723 17193
rect 31665 17184 31677 17187
rect 31628 17156 31677 17184
rect 31628 17144 31634 17156
rect 31665 17153 31677 17156
rect 31711 17153 31723 17187
rect 31665 17147 31723 17153
rect 31757 17187 31815 17193
rect 31757 17153 31769 17187
rect 31803 17184 31815 17187
rect 32398 17184 32404 17196
rect 31803 17156 32404 17184
rect 31803 17153 31815 17156
rect 31757 17147 31815 17153
rect 32398 17144 32404 17156
rect 32456 17184 32462 17196
rect 32766 17184 32772 17196
rect 32456 17156 32772 17184
rect 32456 17144 32462 17156
rect 32766 17144 32772 17156
rect 32824 17144 32830 17196
rect 32876 17184 32904 17280
rect 33137 17187 33195 17193
rect 33137 17184 33149 17187
rect 32876 17156 33149 17184
rect 33137 17153 33149 17156
rect 33183 17153 33195 17187
rect 33137 17147 33195 17153
rect 33321 17187 33379 17193
rect 33321 17153 33333 17187
rect 33367 17153 33379 17187
rect 33321 17147 33379 17153
rect 33336 17116 33364 17147
rect 30340 17088 30512 17116
rect 31726 17088 33364 17116
rect 30340 17076 30346 17088
rect 24044 17020 25176 17048
rect 31481 17051 31539 17057
rect 12618 16980 12624 16992
rect 11900 16952 12624 16980
rect 11793 16943 11851 16949
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 20438 16980 20444 16992
rect 20399 16952 20444 16980
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 24044 16980 24072 17020
rect 31481 17017 31493 17051
rect 31527 17048 31539 17051
rect 31726 17048 31754 17088
rect 31527 17020 31754 17048
rect 31527 17017 31539 17020
rect 31481 17011 31539 17017
rect 23440 16952 24072 16980
rect 23440 16940 23446 16952
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 24489 16983 24547 16989
rect 24489 16980 24501 16983
rect 24452 16952 24501 16980
rect 24452 16940 24458 16952
rect 24489 16949 24501 16952
rect 24535 16949 24547 16983
rect 24489 16943 24547 16949
rect 24762 16940 24768 16992
rect 24820 16980 24826 16992
rect 31294 16980 31300 16992
rect 24820 16952 31300 16980
rect 24820 16940 24826 16952
rect 31294 16940 31300 16952
rect 31352 16940 31358 16992
rect 32493 16983 32551 16989
rect 32493 16949 32505 16983
rect 32539 16980 32551 16983
rect 32766 16980 32772 16992
rect 32539 16952 32772 16980
rect 32539 16949 32551 16952
rect 32493 16943 32551 16949
rect 32766 16940 32772 16952
rect 32824 16940 32830 16992
rect 1104 16890 34868 16912
rect 1104 16838 5170 16890
rect 5222 16838 5234 16890
rect 5286 16838 5298 16890
rect 5350 16838 5362 16890
rect 5414 16838 5426 16890
rect 5478 16838 13611 16890
rect 13663 16838 13675 16890
rect 13727 16838 13739 16890
rect 13791 16838 13803 16890
rect 13855 16838 13867 16890
rect 13919 16838 22052 16890
rect 22104 16838 22116 16890
rect 22168 16838 22180 16890
rect 22232 16838 22244 16890
rect 22296 16838 22308 16890
rect 22360 16838 30493 16890
rect 30545 16838 30557 16890
rect 30609 16838 30621 16890
rect 30673 16838 30685 16890
rect 30737 16838 30749 16890
rect 30801 16838 34868 16890
rect 1104 16816 34868 16838
rect 2682 16736 2688 16788
rect 2740 16776 2746 16788
rect 3234 16776 3240 16788
rect 2740 16736 2774 16776
rect 3195 16748 3240 16776
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 6546 16736 6552 16788
rect 6604 16776 6610 16788
rect 6825 16779 6883 16785
rect 6825 16776 6837 16779
rect 6604 16748 6837 16776
rect 6604 16736 6610 16748
rect 6825 16745 6837 16748
rect 6871 16745 6883 16779
rect 11054 16776 11060 16788
rect 6825 16739 6883 16745
rect 7024 16748 11060 16776
rect 2746 16708 2774 16736
rect 3053 16711 3111 16717
rect 3053 16708 3065 16711
rect 2746 16680 3065 16708
rect 3053 16677 3065 16680
rect 3099 16677 3111 16711
rect 3053 16671 3111 16677
rect 5905 16711 5963 16717
rect 5905 16677 5917 16711
rect 5951 16708 5963 16711
rect 6638 16708 6644 16720
rect 5951 16680 6644 16708
rect 5951 16677 5963 16680
rect 5905 16671 5963 16677
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 7024 16640 7052 16748
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 12250 16776 12256 16788
rect 12211 16748 12256 16776
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 15930 16776 15936 16788
rect 15528 16748 15936 16776
rect 15528 16736 15534 16748
rect 15930 16736 15936 16748
rect 15988 16776 15994 16788
rect 19426 16776 19432 16788
rect 15988 16748 19432 16776
rect 15988 16736 15994 16748
rect 19426 16736 19432 16748
rect 19484 16776 19490 16788
rect 19484 16748 20944 16776
rect 19484 16736 19490 16748
rect 7190 16708 7196 16720
rect 7151 16680 7196 16708
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 8202 16668 8208 16720
rect 8260 16708 8266 16720
rect 9769 16711 9827 16717
rect 9769 16708 9781 16711
rect 8260 16680 9781 16708
rect 8260 16668 8266 16680
rect 9769 16677 9781 16680
rect 9815 16677 9827 16711
rect 10962 16708 10968 16720
rect 9769 16671 9827 16677
rect 9876 16680 10968 16708
rect 4264 16612 7052 16640
rect 7101 16643 7159 16649
rect 4264 16584 4292 16612
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7282 16640 7288 16652
rect 7340 16649 7346 16652
rect 7340 16643 7380 16649
rect 7232 16612 7288 16640
rect 7101 16603 7159 16609
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4246 16572 4252 16584
rect 4207 16544 4252 16572
rect 4065 16535 4123 16541
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 3108 16476 3433 16504
rect 3108 16464 3114 16476
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 4080 16504 4108 16535
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 6454 16532 6460 16584
rect 6512 16572 6518 16584
rect 7116 16572 7144 16603
rect 7282 16600 7288 16612
rect 7368 16640 7380 16643
rect 9876 16640 9904 16680
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 14829 16711 14887 16717
rect 14829 16677 14841 16711
rect 14875 16708 14887 16711
rect 15194 16708 15200 16720
rect 14875 16680 15200 16708
rect 14875 16677 14887 16680
rect 14829 16671 14887 16677
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 20916 16708 20944 16748
rect 20990 16736 20996 16788
rect 21048 16776 21054 16788
rect 21361 16779 21419 16785
rect 21361 16776 21373 16779
rect 21048 16748 21373 16776
rect 21048 16736 21054 16748
rect 21361 16745 21373 16748
rect 21407 16745 21419 16779
rect 26142 16776 26148 16788
rect 21361 16739 21419 16745
rect 22066 16748 26148 16776
rect 22066 16708 22094 16748
rect 26142 16736 26148 16748
rect 26200 16736 26206 16788
rect 31110 16736 31116 16788
rect 31168 16776 31174 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 31168 16748 31217 16776
rect 31168 16736 31174 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 31205 16739 31263 16745
rect 31294 16736 31300 16788
rect 31352 16776 31358 16788
rect 32214 16776 32220 16788
rect 31352 16748 31754 16776
rect 32175 16748 32220 16776
rect 31352 16736 31358 16748
rect 31570 16708 31576 16720
rect 20916 16680 22094 16708
rect 29840 16680 31576 16708
rect 7368 16612 9904 16640
rect 7368 16609 7380 16612
rect 7340 16603 7380 16609
rect 7340 16600 7346 16603
rect 12434 16600 12440 16652
rect 12492 16600 12498 16652
rect 14734 16600 14740 16652
rect 14792 16640 14798 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 14792 16612 15301 16640
rect 14792 16600 14798 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 17494 16640 17500 16652
rect 17455 16612 17500 16640
rect 15289 16603 15347 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 26108 16612 26556 16640
rect 26108 16600 26114 16612
rect 9677 16575 9735 16581
rect 9677 16572 9689 16575
rect 6512 16544 9689 16572
rect 6512 16532 6518 16544
rect 9677 16541 9689 16544
rect 9723 16541 9735 16575
rect 9950 16572 9956 16584
rect 9911 16544 9956 16572
rect 9677 16535 9735 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 10100 16544 10145 16572
rect 10100 16532 10106 16544
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 12066 16572 12072 16584
rect 11112 16544 12072 16572
rect 11112 16532 11118 16544
rect 12066 16532 12072 16544
rect 12124 16572 12130 16584
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 12124 16544 12173 16572
rect 12124 16532 12130 16544
rect 12161 16541 12173 16544
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16566 12403 16575
rect 12452 16566 12480 16600
rect 12391 16541 12480 16566
rect 12345 16538 12480 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 12345 16535 12403 16538
rect 14369 16535 14427 16541
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 15378 16572 15384 16584
rect 14691 16544 15384 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 5074 16504 5080 16516
rect 4080 16476 5080 16504
rect 3421 16467 3479 16473
rect 5074 16464 5080 16476
rect 5132 16464 5138 16516
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16504 5595 16507
rect 7469 16507 7527 16513
rect 5583 16476 6592 16504
rect 5583 16473 5595 16476
rect 5537 16467 5595 16473
rect 6564 16448 6592 16476
rect 7469 16473 7481 16507
rect 7515 16504 7527 16507
rect 11146 16504 11152 16516
rect 7515 16476 11152 16504
rect 7515 16473 7527 16476
rect 7469 16467 7527 16473
rect 3221 16439 3279 16445
rect 3221 16405 3233 16439
rect 3267 16436 3279 16439
rect 5997 16439 6055 16445
rect 5997 16436 6009 16439
rect 3267 16408 6009 16436
rect 3267 16405 3279 16408
rect 3221 16399 3279 16405
rect 5997 16405 6009 16408
rect 6043 16436 6055 16439
rect 6362 16436 6368 16448
rect 6043 16408 6368 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 6546 16396 6552 16448
rect 6604 16436 6610 16448
rect 7484 16436 7512 16467
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 14274 16464 14280 16516
rect 14332 16504 14338 16516
rect 14384 16504 14412 16535
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15556 16575 15614 16581
rect 15556 16541 15568 16575
rect 15602 16572 15614 16575
rect 16574 16572 16580 16584
rect 15602 16544 16580 16572
rect 15602 16541 15614 16544
rect 15556 16535 15614 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17218 16572 17224 16584
rect 17179 16544 17224 16572
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16572 19487 16575
rect 19518 16572 19524 16584
rect 19475 16544 19524 16572
rect 19475 16541 19487 16544
rect 19429 16535 19487 16541
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 19696 16575 19754 16581
rect 19696 16541 19708 16575
rect 19742 16572 19754 16575
rect 20438 16572 20444 16584
rect 19742 16544 20444 16572
rect 19742 16541 19754 16544
rect 19696 16535 19754 16541
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16541 21603 16575
rect 24578 16572 24584 16584
rect 24539 16544 24584 16572
rect 21545 16535 21603 16541
rect 17310 16504 17316 16516
rect 14332 16476 17316 16504
rect 14332 16464 14338 16476
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 19242 16464 19248 16516
rect 19300 16504 19306 16516
rect 21560 16504 21588 16535
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 26421 16575 26479 16581
rect 26421 16572 26433 16575
rect 24688 16544 26433 16572
rect 22462 16504 22468 16516
rect 19300 16476 22468 16504
rect 19300 16464 19306 16476
rect 22462 16464 22468 16476
rect 22520 16504 22526 16516
rect 24688 16504 24716 16544
rect 26421 16541 26433 16544
rect 26467 16541 26479 16575
rect 26528 16572 26556 16612
rect 28994 16600 29000 16652
rect 29052 16640 29058 16652
rect 29730 16640 29736 16652
rect 29052 16612 29736 16640
rect 29052 16600 29058 16612
rect 29730 16600 29736 16612
rect 29788 16600 29794 16652
rect 26528 16544 26740 16572
rect 26421 16535 26479 16541
rect 26712 16516 26740 16544
rect 22520 16476 24716 16504
rect 24848 16507 24906 16513
rect 22520 16464 22526 16476
rect 24848 16473 24860 16507
rect 24894 16504 24906 16507
rect 26050 16504 26056 16516
rect 24894 16476 26056 16504
rect 24894 16473 24906 16476
rect 24848 16467 24906 16473
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 26694 16504 26700 16516
rect 26655 16476 26700 16504
rect 26694 16464 26700 16476
rect 26752 16464 26758 16516
rect 29086 16464 29092 16516
rect 29144 16504 29150 16516
rect 29840 16504 29868 16680
rect 31386 16640 31392 16652
rect 31220 16612 31392 16640
rect 31220 16581 31248 16612
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 31496 16581 31524 16680
rect 31570 16668 31576 16680
rect 31628 16668 31634 16720
rect 31726 16708 31754 16748
rect 32214 16736 32220 16748
rect 32272 16736 32278 16788
rect 33686 16708 33692 16720
rect 31726 16680 33692 16708
rect 33686 16668 33692 16680
rect 33744 16668 33750 16720
rect 32582 16640 32588 16652
rect 31726 16612 32588 16640
rect 29917 16575 29975 16581
rect 29917 16541 29929 16575
rect 29963 16572 29975 16575
rect 31205 16575 31263 16581
rect 31205 16572 31217 16575
rect 29963 16544 31217 16572
rect 29963 16541 29975 16544
rect 29917 16535 29975 16541
rect 31205 16541 31217 16544
rect 31251 16541 31263 16575
rect 31205 16535 31263 16541
rect 31481 16575 31539 16581
rect 31481 16541 31493 16575
rect 31527 16541 31539 16575
rect 31481 16535 31539 16541
rect 31609 16575 31667 16581
rect 31609 16541 31621 16575
rect 31655 16572 31667 16575
rect 31726 16572 31754 16612
rect 32582 16600 32588 16612
rect 32640 16600 32646 16652
rect 31655 16544 31754 16572
rect 31655 16541 31667 16544
rect 31609 16535 31667 16541
rect 32030 16532 32036 16584
rect 32088 16572 32094 16584
rect 32401 16575 32459 16581
rect 32401 16572 32413 16575
rect 32088 16544 32413 16572
rect 32088 16532 32094 16544
rect 32401 16541 32413 16544
rect 32447 16541 32459 16575
rect 32401 16535 32459 16541
rect 30009 16507 30067 16513
rect 30009 16504 30021 16507
rect 29144 16476 30021 16504
rect 29144 16464 29150 16476
rect 30009 16473 30021 16476
rect 30055 16473 30067 16507
rect 31389 16507 31447 16513
rect 31389 16504 31401 16507
rect 30009 16467 30067 16473
rect 30116 16476 31401 16504
rect 30116 16448 30144 16476
rect 31389 16473 31401 16476
rect 31435 16473 31447 16507
rect 32048 16504 32076 16532
rect 31389 16467 31447 16473
rect 31726 16476 32076 16504
rect 6604 16408 7512 16436
rect 10229 16439 10287 16445
rect 6604 16396 6610 16408
rect 10229 16405 10241 16439
rect 10275 16436 10287 16439
rect 10410 16436 10416 16448
rect 10275 16408 10416 16436
rect 10275 16405 10287 16408
rect 10229 16399 10287 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 14458 16436 14464 16448
rect 14419 16408 14464 16436
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 16669 16439 16727 16445
rect 16669 16405 16681 16439
rect 16715 16436 16727 16439
rect 17586 16436 17592 16448
rect 16715 16408 17592 16436
rect 16715 16405 16727 16408
rect 16669 16399 16727 16405
rect 17586 16396 17592 16408
rect 17644 16396 17650 16448
rect 20809 16439 20867 16445
rect 20809 16405 20821 16439
rect 20855 16436 20867 16439
rect 21174 16436 21180 16448
rect 20855 16408 21180 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 25958 16436 25964 16448
rect 25919 16408 25964 16436
rect 25958 16396 25964 16408
rect 26016 16396 26022 16448
rect 30098 16396 30104 16448
rect 30156 16436 30162 16448
rect 30282 16436 30288 16448
rect 30156 16408 30201 16436
rect 30243 16408 30288 16436
rect 30156 16396 30162 16408
rect 30282 16396 30288 16408
rect 30340 16396 30346 16448
rect 31404 16436 31432 16467
rect 31726 16436 31754 16476
rect 31404 16408 31754 16436
rect 1104 16346 35027 16368
rect 1104 16294 9390 16346
rect 9442 16294 9454 16346
rect 9506 16294 9518 16346
rect 9570 16294 9582 16346
rect 9634 16294 9646 16346
rect 9698 16294 17831 16346
rect 17883 16294 17895 16346
rect 17947 16294 17959 16346
rect 18011 16294 18023 16346
rect 18075 16294 18087 16346
rect 18139 16294 26272 16346
rect 26324 16294 26336 16346
rect 26388 16294 26400 16346
rect 26452 16294 26464 16346
rect 26516 16294 26528 16346
rect 26580 16294 34713 16346
rect 34765 16294 34777 16346
rect 34829 16294 34841 16346
rect 34893 16294 34905 16346
rect 34957 16294 34969 16346
rect 35021 16294 35027 16346
rect 1104 16272 35027 16294
rect 5534 16232 5540 16244
rect 5447 16204 5540 16232
rect 5534 16192 5540 16204
rect 5592 16232 5598 16244
rect 6454 16232 6460 16244
rect 5592 16204 6460 16232
rect 5592 16192 5598 16204
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 6730 16232 6736 16244
rect 6691 16204 6736 16232
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 12250 16232 12256 16244
rect 11011 16204 12256 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13412 16204 13461 16232
rect 13412 16192 13418 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 19242 16232 19248 16244
rect 13449 16195 13507 16201
rect 14016 16204 19248 16232
rect 5552 16164 5580 16192
rect 5718 16164 5724 16176
rect 5460 16136 5580 16164
rect 5631 16136 5724 16164
rect 5460 16105 5488 16136
rect 5718 16124 5724 16136
rect 5776 16164 5782 16176
rect 6822 16164 6828 16176
rect 5776 16136 6828 16164
rect 5776 16124 5782 16136
rect 6822 16124 6828 16136
rect 6880 16124 6886 16176
rect 7282 16164 7288 16176
rect 7116 16136 7288 16164
rect 5445 16099 5503 16105
rect 5445 16065 5457 16099
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16065 5595 16099
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 5537 16059 5595 16065
rect 5552 16028 5580 16059
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 6733 16099 6791 16105
rect 6733 16096 6745 16099
rect 6696 16068 6745 16096
rect 6696 16056 6702 16068
rect 6733 16065 6745 16068
rect 6779 16096 6791 16099
rect 7116 16096 7144 16136
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 8849 16167 8907 16173
rect 8849 16133 8861 16167
rect 8895 16164 8907 16167
rect 11514 16164 11520 16176
rect 8895 16136 11520 16164
rect 8895 16133 8907 16136
rect 8849 16127 8907 16133
rect 11514 16124 11520 16136
rect 11572 16124 11578 16176
rect 6779 16068 7144 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7248 16068 7389 16096
rect 7248 16056 7254 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 7466 16056 7472 16108
rect 7524 16096 7530 16108
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 7524 16068 8769 16096
rect 7524 16056 7530 16068
rect 8757 16065 8769 16068
rect 8803 16065 8815 16099
rect 10410 16096 10416 16108
rect 10371 16068 10416 16096
rect 8757 16059 8815 16065
rect 10410 16056 10416 16068
rect 10468 16056 10474 16108
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11146 16096 11152 16108
rect 11107 16068 11152 16096
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 12406 16068 13277 16096
rect 7098 16028 7104 16040
rect 5552 16000 7104 16028
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 6454 15920 6460 15972
rect 6512 15960 6518 15972
rect 7668 15960 7696 15991
rect 6512 15932 7696 15960
rect 7929 15963 7987 15969
rect 6512 15920 6518 15932
rect 7929 15929 7941 15963
rect 7975 15960 7987 15963
rect 12406 15960 12434 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13464 16096 13492 16195
rect 14016 16105 14044 16204
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19518 16232 19524 16244
rect 19479 16204 19524 16232
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 20441 16235 20499 16241
rect 20441 16201 20453 16235
rect 20487 16232 20499 16235
rect 20530 16232 20536 16244
rect 20487 16204 20536 16232
rect 20487 16201 20499 16204
rect 20441 16195 20499 16201
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 22646 16232 22652 16244
rect 20732 16204 22508 16232
rect 22607 16204 22652 16232
rect 14274 16164 14280 16176
rect 14235 16136 14280 16164
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 15194 16173 15200 16176
rect 15188 16164 15200 16173
rect 15155 16136 15200 16164
rect 15188 16127 15200 16136
rect 15194 16124 15200 16127
rect 15252 16124 15258 16176
rect 18230 16164 18236 16176
rect 18191 16136 18236 16164
rect 18230 16124 18236 16136
rect 18288 16124 18294 16176
rect 20732 16173 20760 16204
rect 20717 16167 20775 16173
rect 20717 16133 20729 16167
rect 20763 16133 20775 16167
rect 20717 16127 20775 16133
rect 21174 16124 21180 16176
rect 21232 16164 21238 16176
rect 22480 16164 22508 16204
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 26050 16232 26056 16244
rect 26011 16204 26056 16232
rect 26050 16192 26056 16204
rect 26108 16192 26114 16244
rect 29086 16232 29092 16244
rect 28552 16204 29092 16232
rect 25958 16164 25964 16176
rect 21232 16136 22140 16164
rect 22480 16136 25964 16164
rect 21232 16124 21238 16136
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13464 16068 14013 16096
rect 13265 16059 13323 16065
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 17402 16096 17408 16108
rect 17363 16068 17408 16096
rect 14001 16059 14059 16065
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 17678 16096 17684 16108
rect 17639 16068 17684 16096
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 20530 16056 20536 16108
rect 20588 16105 20594 16108
rect 20588 16099 20637 16105
rect 20588 16065 20591 16099
rect 20625 16065 20637 16099
rect 20588 16059 20637 16065
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 20588 16056 20594 16059
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14792 16000 14933 16028
rect 14792 15988 14798 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 17773 16031 17831 16037
rect 17773 15997 17785 16031
rect 17819 16028 17831 16031
rect 19610 16028 19616 16040
rect 17819 16000 19616 16028
rect 17819 15997 17831 16000
rect 17773 15991 17831 15997
rect 19610 15988 19616 16000
rect 19668 16028 19674 16040
rect 20824 16028 20852 16059
rect 20898 16056 20904 16108
rect 20956 16105 20962 16108
rect 20956 16099 20995 16105
rect 20983 16065 20995 16099
rect 21082 16096 21088 16108
rect 21043 16068 21088 16096
rect 20956 16059 20995 16065
rect 20956 16056 20962 16059
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22112 16105 22140 16136
rect 25958 16124 25964 16136
rect 26016 16164 26022 16176
rect 26421 16167 26479 16173
rect 26421 16164 26433 16167
rect 26016 16136 26433 16164
rect 26016 16124 26022 16136
rect 26421 16133 26433 16136
rect 26467 16133 26479 16167
rect 26421 16127 26479 16133
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21968 16068 22017 16096
rect 21968 16056 21974 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22098 16099 22156 16105
rect 22098 16065 22110 16099
rect 22144 16065 22156 16099
rect 22098 16059 22156 16065
rect 22281 16099 22339 16105
rect 22281 16065 22293 16099
rect 22327 16065 22339 16099
rect 22281 16059 22339 16065
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 22511 16099 22569 16105
rect 22511 16065 22523 16099
rect 22557 16096 22569 16099
rect 23106 16096 23112 16108
rect 22557 16068 23112 16096
rect 22557 16065 22569 16068
rect 22511 16059 22569 16065
rect 19668 16000 20944 16028
rect 19668 15988 19674 16000
rect 7975 15932 12434 15960
rect 20916 15960 20944 16000
rect 22296 15960 22324 16059
rect 20916 15932 22324 15960
rect 22388 15960 22416 16059
rect 23106 16056 23112 16068
rect 23164 16056 23170 16108
rect 25130 16096 25136 16108
rect 25091 16068 25136 16096
rect 25130 16056 25136 16068
rect 25188 16056 25194 16108
rect 26234 16096 26240 16108
rect 26195 16068 26240 16096
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 26513 16099 26571 16105
rect 26513 16065 26525 16099
rect 26559 16096 26571 16099
rect 26602 16096 26608 16108
rect 26559 16068 26608 16096
rect 26559 16065 26571 16068
rect 26513 16059 26571 16065
rect 26602 16056 26608 16068
rect 26660 16056 26666 16108
rect 27706 16056 27712 16108
rect 27764 16096 27770 16108
rect 28552 16105 28580 16204
rect 29086 16192 29092 16204
rect 29144 16192 29150 16244
rect 32582 16192 32588 16244
rect 32640 16232 32646 16244
rect 33042 16232 33048 16244
rect 32640 16204 33048 16232
rect 32640 16192 32646 16204
rect 33042 16192 33048 16204
rect 33100 16232 33106 16244
rect 33689 16235 33747 16241
rect 33689 16232 33701 16235
rect 33100 16204 33701 16232
rect 33100 16192 33106 16204
rect 33689 16201 33701 16204
rect 33735 16201 33747 16235
rect 33689 16195 33747 16201
rect 28629 16167 28687 16173
rect 28629 16133 28641 16167
rect 28675 16164 28687 16167
rect 31386 16164 31392 16176
rect 28675 16136 31392 16164
rect 28675 16133 28687 16136
rect 28629 16127 28687 16133
rect 31386 16124 31392 16136
rect 31444 16164 31450 16176
rect 33226 16164 33232 16176
rect 31444 16136 33232 16164
rect 31444 16124 31450 16136
rect 33226 16124 33232 16136
rect 33284 16124 33290 16176
rect 28537 16099 28595 16105
rect 28537 16096 28549 16099
rect 27764 16068 28549 16096
rect 27764 16056 27770 16068
rect 28537 16065 28549 16068
rect 28583 16065 28595 16099
rect 28537 16059 28595 16065
rect 28721 16099 28779 16105
rect 28721 16065 28733 16099
rect 28767 16065 28779 16099
rect 28721 16059 28779 16065
rect 28905 16099 28963 16105
rect 28905 16065 28917 16099
rect 28951 16096 28963 16099
rect 28994 16096 29000 16108
rect 28951 16068 29000 16096
rect 28951 16065 28963 16068
rect 28905 16059 28963 16065
rect 24394 15988 24400 16040
rect 24452 16028 24458 16040
rect 28736 16028 28764 16059
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 29549 16099 29607 16105
rect 29549 16065 29561 16099
rect 29595 16096 29607 16099
rect 30282 16096 30288 16108
rect 29595 16068 30288 16096
rect 29595 16065 29607 16068
rect 29549 16059 29607 16065
rect 30282 16056 30288 16068
rect 30340 16056 30346 16108
rect 32576 16099 32634 16105
rect 32576 16065 32588 16099
rect 32622 16096 32634 16099
rect 33870 16096 33876 16108
rect 32622 16068 33876 16096
rect 32622 16065 32634 16068
rect 32576 16059 32634 16065
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 30098 16028 30104 16040
rect 24452 16000 30104 16028
rect 24452 15988 24458 16000
rect 30098 15988 30104 16000
rect 30156 15988 30162 16040
rect 32306 16028 32312 16040
rect 32267 16000 32312 16028
rect 32306 15988 32312 16000
rect 32364 15988 32370 16040
rect 32214 15960 32220 15972
rect 22388 15932 32220 15960
rect 7975 15929 7987 15932
rect 7929 15923 7987 15929
rect 32214 15920 32220 15932
rect 32272 15920 32278 15972
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 16301 15895 16359 15901
rect 16301 15892 16313 15895
rect 14516 15864 16313 15892
rect 14516 15852 14522 15864
rect 16301 15861 16313 15864
rect 16347 15892 16359 15895
rect 20070 15892 20076 15904
rect 16347 15864 20076 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 24578 15892 24584 15904
rect 23891 15864 24584 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 28353 15895 28411 15901
rect 28353 15892 28365 15895
rect 28224 15864 28365 15892
rect 28224 15852 28230 15864
rect 28353 15861 28365 15864
rect 28399 15861 28411 15895
rect 29454 15892 29460 15904
rect 29415 15864 29460 15892
rect 28353 15855 28411 15861
rect 29454 15852 29460 15864
rect 29512 15852 29518 15904
rect 1104 15802 34868 15824
rect 1104 15750 5170 15802
rect 5222 15750 5234 15802
rect 5286 15750 5298 15802
rect 5350 15750 5362 15802
rect 5414 15750 5426 15802
rect 5478 15750 13611 15802
rect 13663 15750 13675 15802
rect 13727 15750 13739 15802
rect 13791 15750 13803 15802
rect 13855 15750 13867 15802
rect 13919 15750 22052 15802
rect 22104 15750 22116 15802
rect 22168 15750 22180 15802
rect 22232 15750 22244 15802
rect 22296 15750 22308 15802
rect 22360 15750 30493 15802
rect 30545 15750 30557 15802
rect 30609 15750 30621 15802
rect 30673 15750 30685 15802
rect 30737 15750 30749 15802
rect 30801 15750 34868 15802
rect 1104 15728 34868 15750
rect 4982 15648 4988 15700
rect 5040 15688 5046 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 5040 15660 5273 15688
rect 5040 15648 5046 15660
rect 5261 15657 5273 15660
rect 5307 15688 5319 15691
rect 7742 15688 7748 15700
rect 5307 15660 7748 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 11054 15688 11060 15700
rect 10919 15660 11060 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 15120 15660 17908 15688
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 2958 15620 2964 15632
rect 2915 15592 2964 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 2958 15580 2964 15592
rect 3016 15580 3022 15632
rect 13633 15623 13691 15629
rect 13633 15589 13645 15623
rect 13679 15620 13691 15623
rect 14550 15620 14556 15632
rect 13679 15592 14556 15620
rect 13679 15589 13691 15592
rect 13633 15583 13691 15589
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 5074 15552 5080 15564
rect 2700 15524 5080 15552
rect 2700 15493 2728 15524
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 6546 15552 6552 15564
rect 6104 15524 6552 15552
rect 6104 15496 6132 15524
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 13446 15512 13452 15564
rect 13504 15552 13510 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 13504 15524 14933 15552
rect 13504 15512 13510 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 4246 15484 4252 15496
rect 3007 15456 4252 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 6086 15484 6092 15496
rect 5999 15456 6092 15484
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 6454 15484 6460 15496
rect 6319 15456 6460 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 12618 15484 12624 15496
rect 12579 15456 12624 15484
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 12713 15487 12771 15493
rect 12713 15453 12725 15487
rect 12759 15484 12771 15487
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 12759 15456 13369 15484
rect 12759 15453 12771 15456
rect 12713 15447 12771 15453
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 14274 15484 14280 15496
rect 13679 15456 14280 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 15120 15493 15148 15660
rect 16574 15620 16580 15632
rect 16040 15592 16580 15620
rect 15105 15487 15163 15493
rect 15105 15453 15117 15487
rect 15151 15453 15163 15487
rect 15105 15447 15163 15453
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15484 15347 15487
rect 15654 15484 15660 15496
rect 15335 15456 15660 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 16040 15493 16068 15592
rect 16574 15580 16580 15592
rect 16632 15620 16638 15632
rect 17402 15620 17408 15632
rect 16632 15592 17408 15620
rect 16632 15580 16638 15592
rect 17402 15580 17408 15592
rect 17460 15580 17466 15632
rect 16117 15555 16175 15561
rect 16117 15521 16129 15555
rect 16163 15552 16175 15555
rect 16390 15552 16396 15564
rect 16163 15524 16396 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 17880 15493 17908 15660
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 26050 15688 26056 15700
rect 25188 15660 26056 15688
rect 25188 15648 25194 15660
rect 26050 15648 26056 15660
rect 26108 15688 26114 15700
rect 26421 15691 26479 15697
rect 26421 15688 26433 15691
rect 26108 15660 26433 15688
rect 26108 15648 26114 15660
rect 26421 15657 26433 15660
rect 26467 15657 26479 15691
rect 26421 15651 26479 15657
rect 31665 15691 31723 15697
rect 31665 15657 31677 15691
rect 31711 15688 31723 15691
rect 31754 15688 31760 15700
rect 31711 15660 31760 15688
rect 31711 15657 31723 15660
rect 31665 15651 31723 15657
rect 31754 15648 31760 15660
rect 31812 15688 31818 15700
rect 32306 15688 32312 15700
rect 31812 15660 32312 15688
rect 31812 15648 31818 15660
rect 32306 15648 32312 15660
rect 32364 15648 32370 15700
rect 33870 15688 33876 15700
rect 33831 15660 33876 15688
rect 33870 15648 33876 15660
rect 33928 15648 33934 15700
rect 21910 15580 21916 15632
rect 21968 15620 21974 15632
rect 27985 15623 28043 15629
rect 27985 15620 27997 15623
rect 21968 15592 27997 15620
rect 21968 15580 21974 15592
rect 27985 15589 27997 15592
rect 28031 15589 28043 15623
rect 27985 15583 28043 15589
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 19978 15552 19984 15564
rect 18279 15524 19984 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 22554 15552 22560 15564
rect 22515 15524 22560 15552
rect 22554 15512 22560 15524
rect 22612 15512 22618 15564
rect 24762 15552 24768 15564
rect 23216 15524 24768 15552
rect 16301 15487 16359 15493
rect 16301 15484 16313 15487
rect 16264 15456 16313 15484
rect 16264 15444 16270 15456
rect 16301 15453 16313 15456
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15484 17923 15487
rect 18322 15484 18328 15496
rect 17911 15456 18328 15484
rect 17911 15453 17923 15456
rect 17865 15447 17923 15453
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 20806 15484 20812 15496
rect 20767 15456 20812 15484
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 23216 15493 23244 15524
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 28166 15552 28172 15564
rect 28127 15524 28172 15552
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 28353 15555 28411 15561
rect 28353 15521 28365 15555
rect 28399 15552 28411 15555
rect 29454 15552 29460 15564
rect 28399 15524 29460 15552
rect 28399 15521 28411 15524
rect 28353 15515 28411 15521
rect 29454 15512 29460 15524
rect 29512 15512 29518 15564
rect 23201 15487 23259 15493
rect 23201 15453 23213 15487
rect 23247 15453 23259 15487
rect 23474 15484 23480 15496
rect 23435 15456 23480 15484
rect 23201 15447 23259 15453
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 27798 15444 27804 15496
rect 27856 15484 27862 15496
rect 28261 15487 28319 15493
rect 28261 15484 28273 15487
rect 27856 15456 28273 15484
rect 27856 15444 27862 15456
rect 28261 15453 28273 15456
rect 28307 15453 28319 15487
rect 28442 15484 28448 15496
rect 28403 15456 28448 15484
rect 28261 15447 28319 15453
rect 28442 15444 28448 15456
rect 28500 15444 28506 15496
rect 33410 15484 33416 15496
rect 33371 15456 33416 15484
rect 33410 15444 33416 15456
rect 33468 15444 33474 15496
rect 33686 15484 33692 15496
rect 33647 15456 33692 15484
rect 33686 15444 33692 15456
rect 33744 15444 33750 15496
rect 5445 15419 5503 15425
rect 5445 15385 5457 15419
rect 5491 15416 5503 15419
rect 5534 15416 5540 15428
rect 5491 15388 5540 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 6181 15419 6239 15425
rect 6181 15385 6193 15419
rect 6227 15416 6239 15419
rect 7190 15416 7196 15428
rect 6227 15388 7196 15416
rect 6227 15385 6239 15388
rect 6181 15379 6239 15385
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 5077 15351 5135 15357
rect 5077 15348 5089 15351
rect 4488 15320 5089 15348
rect 4488 15308 4494 15320
rect 5077 15317 5089 15320
rect 5123 15317 5135 15351
rect 5077 15311 5135 15317
rect 5245 15351 5303 15357
rect 5245 15317 5257 15351
rect 5291 15348 5303 15351
rect 6196 15348 6224 15379
rect 7190 15376 7196 15388
rect 7248 15376 7254 15428
rect 12066 15376 12072 15428
rect 12124 15416 12130 15428
rect 12161 15419 12219 15425
rect 12161 15416 12173 15419
rect 12124 15388 12173 15416
rect 12124 15376 12130 15388
rect 12161 15385 12173 15388
rect 12207 15416 12219 15419
rect 17310 15416 17316 15428
rect 12207 15388 17316 15416
rect 12207 15385 12219 15388
rect 12161 15379 12219 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17678 15416 17684 15428
rect 17639 15388 17684 15416
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 22370 15376 22376 15428
rect 22428 15416 22434 15428
rect 23382 15416 23388 15428
rect 22428 15388 23388 15416
rect 22428 15376 22434 15388
rect 23382 15376 23388 15388
rect 23440 15376 23446 15428
rect 25130 15416 25136 15428
rect 25091 15388 25136 15416
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 32953 15419 33011 15425
rect 32953 15385 32965 15419
rect 32999 15416 33011 15419
rect 33594 15416 33600 15428
rect 32999 15388 33600 15416
rect 32999 15385 33011 15388
rect 32953 15379 33011 15385
rect 33594 15376 33600 15388
rect 33652 15376 33658 15428
rect 6822 15348 6828 15360
rect 5291 15320 6224 15348
rect 6783 15320 6828 15348
rect 5291 15317 5303 15320
rect 5245 15311 5303 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 23017 15351 23075 15357
rect 23017 15348 23029 15351
rect 21048 15320 23029 15348
rect 21048 15308 21054 15320
rect 23017 15317 23029 15320
rect 23063 15317 23075 15351
rect 23017 15311 23075 15317
rect 33042 15308 33048 15360
rect 33100 15348 33106 15360
rect 33505 15351 33563 15357
rect 33505 15348 33517 15351
rect 33100 15320 33517 15348
rect 33100 15308 33106 15320
rect 33505 15317 33517 15320
rect 33551 15317 33563 15351
rect 33505 15311 33563 15317
rect 1104 15258 35027 15280
rect 1104 15206 9390 15258
rect 9442 15206 9454 15258
rect 9506 15206 9518 15258
rect 9570 15206 9582 15258
rect 9634 15206 9646 15258
rect 9698 15206 17831 15258
rect 17883 15206 17895 15258
rect 17947 15206 17959 15258
rect 18011 15206 18023 15258
rect 18075 15206 18087 15258
rect 18139 15206 26272 15258
rect 26324 15206 26336 15258
rect 26388 15206 26400 15258
rect 26452 15206 26464 15258
rect 26516 15206 26528 15258
rect 26580 15206 34713 15258
rect 34765 15206 34777 15258
rect 34829 15206 34841 15258
rect 34893 15206 34905 15258
rect 34957 15206 34969 15258
rect 35021 15206 35027 15258
rect 1104 15184 35027 15206
rect 5436 15147 5494 15153
rect 5436 15113 5448 15147
rect 5482 15144 5494 15147
rect 5718 15144 5724 15156
rect 5482 15116 5724 15144
rect 5482 15113 5494 15116
rect 5436 15107 5494 15113
rect 5718 15104 5724 15116
rect 5776 15144 5782 15156
rect 6362 15144 6368 15156
rect 5776 15116 6368 15144
rect 5776 15104 5782 15116
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 18414 15144 18420 15156
rect 16071 15116 18420 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 21818 15144 21824 15156
rect 19260 15116 21824 15144
rect 2958 15036 2964 15088
rect 3016 15036 3022 15088
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6454 15076 6460 15088
rect 5859 15048 6460 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6454 15036 6460 15048
rect 6512 15036 6518 15088
rect 9677 15079 9735 15085
rect 9677 15045 9689 15079
rect 9723 15076 9735 15079
rect 11974 15076 11980 15088
rect 9723 15048 11980 15076
rect 9723 15045 9735 15048
rect 9677 15039 9735 15045
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 17405 15079 17463 15085
rect 16224 15048 17080 15076
rect 16224 15020 16252 15048
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4522 15008 4528 15020
rect 4203 14980 4528 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 1670 14940 1676 14952
rect 1631 14912 1676 14940
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2682 14940 2688 14952
rect 1995 14912 2688 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2682 14900 2688 14912
rect 2740 14940 2746 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 2740 14912 4077 14940
rect 2740 14900 2746 14912
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 3234 14832 3240 14884
rect 3292 14872 3298 14884
rect 3421 14875 3479 14881
rect 3421 14872 3433 14875
rect 3292 14844 3433 14872
rect 3292 14832 3298 14844
rect 3421 14841 3433 14844
rect 3467 14872 3479 14875
rect 4172 14872 4200 14971
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 9030 15008 9036 15020
rect 8991 14980 9036 15008
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 9766 15008 9772 15020
rect 9263 14980 9772 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 10376 14980 10425 15008
rect 10376 14968 10382 14980
rect 10413 14977 10425 14980
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 10505 15011 10563 15017
rect 10505 14977 10517 15011
rect 10551 14977 10563 15011
rect 10686 15008 10692 15020
rect 10647 14980 10692 15008
rect 10505 14971 10563 14977
rect 8938 14940 8944 14952
rect 8851 14912 8944 14940
rect 8938 14900 8944 14912
rect 8996 14940 9002 14952
rect 9858 14940 9864 14952
rect 8996 14912 9864 14940
rect 8996 14900 9002 14912
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 3467 14844 4200 14872
rect 10428 14872 10456 14971
rect 10520 14940 10548 14971
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 12158 15008 12164 15020
rect 10796 14980 12164 15008
rect 10796 14940 10824 14980
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 13446 15008 13452 15020
rect 12406 14980 13452 15008
rect 11146 14940 11152 14952
rect 10520 14912 10824 14940
rect 11107 14912 11152 14940
rect 11146 14900 11152 14912
rect 11204 14900 11210 14952
rect 12406 14872 12434 14980
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 15654 14968 15660 15020
rect 15712 15008 15718 15020
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15712 14980 16129 15008
rect 15712 14968 15718 14980
rect 16117 14977 16129 14980
rect 16163 15008 16175 15011
rect 16206 15008 16212 15020
rect 16163 14980 16212 15008
rect 16163 14977 16175 14980
rect 16117 14971 16175 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 17052 15017 17080 15048
rect 17405 15045 17417 15079
rect 17451 15076 17463 15079
rect 19260 15076 19288 15116
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22278 15144 22284 15156
rect 22191 15116 22284 15144
rect 22278 15104 22284 15116
rect 22336 15144 22342 15156
rect 23382 15144 23388 15156
rect 22336 15116 23388 15144
rect 22336 15104 22342 15116
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 23477 15147 23535 15153
rect 23477 15113 23489 15147
rect 23523 15144 23535 15147
rect 25130 15144 25136 15156
rect 23523 15116 25136 15144
rect 23523 15113 23535 15116
rect 23477 15107 23535 15113
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 33594 15144 33600 15156
rect 33555 15116 33600 15144
rect 33594 15104 33600 15116
rect 33652 15104 33658 15156
rect 17451 15048 19288 15076
rect 17451 15045 17463 15048
rect 17405 15039 17463 15045
rect 19334 15036 19340 15088
rect 19392 15076 19398 15088
rect 21910 15076 21916 15088
rect 19392 15048 21916 15076
rect 19392 15036 19398 15048
rect 21910 15036 21916 15048
rect 21968 15076 21974 15088
rect 23109 15079 23167 15085
rect 23109 15076 23121 15079
rect 21968 15048 23121 15076
rect 21968 15036 21974 15048
rect 23109 15045 23121 15048
rect 23155 15045 23167 15079
rect 23109 15039 23167 15045
rect 23293 15079 23351 15085
rect 23293 15045 23305 15079
rect 23339 15076 23351 15079
rect 23339 15048 23428 15076
rect 23339 15045 23351 15048
rect 23293 15039 23351 15045
rect 23400 15020 23428 15048
rect 26694 15036 26700 15088
rect 26752 15076 26758 15088
rect 29825 15079 29883 15085
rect 29825 15076 29837 15079
rect 26752 15048 29837 15076
rect 26752 15036 26758 15048
rect 29825 15045 29837 15048
rect 29871 15045 29883 15079
rect 29825 15039 29883 15045
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 17037 15011 17095 15017
rect 16899 14980 16988 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 16316 14940 16344 14971
rect 16960 14940 16988 14980
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 18230 15008 18236 15020
rect 18191 14980 18236 15008
rect 17037 14971 17095 14977
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 20346 14968 20352 15020
rect 20404 15008 20410 15020
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 20404 14980 20637 15008
rect 20404 14968 20410 14980
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20806 15008 20812 15020
rect 20767 14980 20812 15008
rect 20625 14971 20683 14977
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 22373 15011 22431 15017
rect 20956 14980 21001 15008
rect 20956 14968 20962 14980
rect 22373 14977 22385 15011
rect 22419 15008 22431 15011
rect 22462 15008 22468 15020
rect 22419 14980 22468 15008
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 23382 14968 23388 15020
rect 23440 14968 23446 15020
rect 25130 15008 25136 15020
rect 25188 15017 25194 15020
rect 25100 14980 25136 15008
rect 25130 14968 25136 14980
rect 25188 14971 25200 15017
rect 25188 14968 25194 14971
rect 29914 14968 29920 15020
rect 29972 15008 29978 15020
rect 32309 15011 32367 15017
rect 32309 15008 32321 15011
rect 29972 14980 32321 15008
rect 29972 14968 29978 14980
rect 32309 14977 32321 14980
rect 32355 14977 32367 15011
rect 32309 14971 32367 14977
rect 18138 14940 18144 14952
rect 16316 14912 16896 14940
rect 16960 14912 18144 14940
rect 16868 14884 16896 14912
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 25409 14943 25467 14949
rect 25409 14909 25421 14943
rect 25455 14940 25467 14943
rect 26418 14940 26424 14952
rect 25455 14912 26424 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 10428 14844 12434 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 16850 14832 16856 14884
rect 16908 14832 16914 14884
rect 19610 14832 19616 14884
rect 19668 14872 19674 14884
rect 22462 14872 22468 14884
rect 19668 14844 22468 14872
rect 19668 14832 19674 14844
rect 22462 14832 22468 14844
rect 22520 14872 22526 14884
rect 23198 14872 23204 14884
rect 22520 14844 23204 14872
rect 22520 14832 22526 14844
rect 23198 14832 23204 14844
rect 23256 14832 23262 14884
rect 29638 14872 29644 14884
rect 29599 14844 29644 14872
rect 29638 14832 29644 14844
rect 29696 14832 29702 14884
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 5261 14807 5319 14813
rect 5261 14804 5273 14807
rect 4304 14776 5273 14804
rect 4304 14764 4310 14776
rect 5261 14773 5273 14776
rect 5307 14773 5319 14807
rect 5261 14767 5319 14773
rect 5445 14807 5503 14813
rect 5445 14773 5457 14807
rect 5491 14804 5503 14807
rect 6086 14804 6092 14816
rect 5491 14776 6092 14804
rect 5491 14773 5503 14776
rect 5445 14767 5503 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 19702 14804 19708 14816
rect 19663 14776 19708 14804
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 20438 14804 20444 14816
rect 20399 14776 20444 14804
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 22278 14804 22284 14816
rect 20956 14776 22284 14804
rect 20956 14764 20962 14776
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 23290 14804 23296 14816
rect 23251 14776 23296 14804
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 24026 14804 24032 14816
rect 23987 14776 24032 14804
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 1104 14714 34868 14736
rect 1104 14662 5170 14714
rect 5222 14662 5234 14714
rect 5286 14662 5298 14714
rect 5350 14662 5362 14714
rect 5414 14662 5426 14714
rect 5478 14662 13611 14714
rect 13663 14662 13675 14714
rect 13727 14662 13739 14714
rect 13791 14662 13803 14714
rect 13855 14662 13867 14714
rect 13919 14662 22052 14714
rect 22104 14662 22116 14714
rect 22168 14662 22180 14714
rect 22232 14662 22244 14714
rect 22296 14662 22308 14714
rect 22360 14662 30493 14714
rect 30545 14662 30557 14714
rect 30609 14662 30621 14714
rect 30673 14662 30685 14714
rect 30737 14662 30749 14714
rect 30801 14662 34868 14714
rect 1104 14640 34868 14662
rect 6181 14603 6239 14609
rect 6181 14569 6193 14603
rect 6227 14600 6239 14603
rect 6822 14600 6828 14612
rect 6227 14572 6828 14600
rect 6227 14569 6239 14572
rect 6181 14563 6239 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7190 14600 7196 14612
rect 7151 14572 7196 14600
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 19484 14572 19625 14600
rect 19484 14560 19490 14572
rect 19613 14569 19625 14572
rect 19659 14600 19671 14603
rect 22097 14603 22155 14609
rect 19659 14572 21680 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 7377 14535 7435 14541
rect 7377 14501 7389 14535
rect 7423 14532 7435 14535
rect 8294 14532 8300 14544
rect 7423 14504 8300 14532
rect 7423 14501 7435 14504
rect 7377 14495 7435 14501
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 8478 14532 8484 14544
rect 8439 14504 8484 14532
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 9217 14535 9275 14541
rect 9217 14501 9229 14535
rect 9263 14532 9275 14535
rect 9306 14532 9312 14544
rect 9263 14504 9312 14532
rect 9263 14501 9275 14504
rect 9217 14495 9275 14501
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 20714 14492 20720 14544
rect 20772 14492 20778 14544
rect 21652 14532 21680 14572
rect 22097 14569 22109 14603
rect 22143 14600 22155 14603
rect 22370 14600 22376 14612
rect 22143 14572 22376 14600
rect 22143 14569 22155 14572
rect 22097 14563 22155 14569
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 25774 14560 25780 14612
rect 25832 14600 25838 14612
rect 25961 14603 26019 14609
rect 25961 14600 25973 14603
rect 25832 14572 25973 14600
rect 25832 14560 25838 14572
rect 25961 14569 25973 14572
rect 26007 14569 26019 14603
rect 25961 14563 26019 14569
rect 26602 14560 26608 14612
rect 26660 14600 26666 14612
rect 33226 14600 33232 14612
rect 26660 14572 28304 14600
rect 33187 14572 33232 14600
rect 26660 14560 26666 14572
rect 23290 14532 23296 14544
rect 21652 14504 23296 14532
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 1394 14424 1400 14476
rect 1452 14464 1458 14476
rect 17310 14464 17316 14476
rect 1452 14436 15608 14464
rect 17223 14436 17316 14464
rect 1452 14424 1458 14436
rect 2682 14396 2688 14408
rect 2643 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 3050 14396 3056 14408
rect 2915 14368 3056 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 6362 14396 6368 14408
rect 6323 14368 6368 14396
rect 6089 14359 6147 14365
rect 2958 14328 2964 14340
rect 2919 14300 2964 14328
rect 2958 14288 2964 14300
rect 3016 14288 3022 14340
rect 6104 14328 6132 14359
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 7190 14396 7196 14408
rect 6472 14368 7196 14396
rect 6472 14328 6500 14368
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7926 14396 7932 14408
rect 7839 14368 7932 14396
rect 7926 14356 7932 14368
rect 7984 14396 7990 14408
rect 7984 14368 9812 14396
rect 7984 14356 7990 14368
rect 9784 14340 9812 14368
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 12802 14396 12808 14408
rect 11112 14368 12808 14396
rect 11112 14356 11118 14368
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 13722 14396 13728 14408
rect 12943 14368 13728 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 6104 14300 6500 14328
rect 6638 14288 6644 14340
rect 6696 14328 6702 14340
rect 7009 14331 7067 14337
rect 7009 14328 7021 14331
rect 6696 14300 7021 14328
rect 6696 14288 6702 14300
rect 7009 14297 7021 14300
rect 7055 14297 7067 14331
rect 7009 14291 7067 14297
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8021 14331 8079 14337
rect 8021 14328 8033 14331
rect 7892 14300 8033 14328
rect 7892 14288 7898 14300
rect 8021 14297 8033 14300
rect 8067 14297 8079 14331
rect 8202 14328 8208 14340
rect 8163 14300 8208 14328
rect 8021 14291 8079 14297
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14297 9551 14331
rect 9766 14328 9772 14340
rect 9679 14300 9772 14328
rect 9493 14291 9551 14297
rect 6549 14263 6607 14269
rect 6549 14229 6561 14263
rect 6595 14260 6607 14263
rect 6914 14260 6920 14272
rect 6595 14232 6920 14260
rect 6595 14229 6607 14232
rect 6549 14223 6607 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 7219 14263 7277 14269
rect 7219 14229 7231 14263
rect 7265 14260 7277 14263
rect 7466 14260 7472 14272
rect 7265 14232 7472 14260
rect 7265 14229 7277 14232
rect 7219 14223 7277 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 9508 14260 9536 14291
rect 9766 14288 9772 14300
rect 9824 14328 9830 14340
rect 10686 14328 10692 14340
rect 9824 14300 10692 14328
rect 9824 14288 9830 14300
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12912 14328 12940 14359
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 15580 14405 15608 14436
rect 17310 14424 17316 14436
rect 17368 14464 17374 14476
rect 20732 14464 20760 14492
rect 24578 14464 24584 14476
rect 17368 14436 20760 14464
rect 24539 14436 24584 14464
rect 17368 14424 17374 14436
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 17678 14356 17684 14408
rect 17736 14396 17742 14408
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17736 14368 17785 14396
rect 17736 14356 17742 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 18196 14368 18245 14396
rect 18196 14356 18202 14368
rect 18233 14365 18245 14368
rect 18279 14396 18291 14399
rect 18414 14396 18420 14408
rect 18279 14368 18420 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18555 14368 19656 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 13078 14328 13084 14340
rect 12492 14300 12940 14328
rect 13039 14300 13084 14328
rect 12492 14288 12498 14300
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 19392 14300 19441 14328
rect 19392 14288 19398 14300
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19628 14328 19656 14368
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20990 14405 20996 14408
rect 20717 14399 20775 14405
rect 20717 14396 20729 14399
rect 19760 14368 20729 14396
rect 19760 14356 19766 14368
rect 20717 14365 20729 14368
rect 20763 14365 20775 14399
rect 20984 14396 20996 14405
rect 20951 14368 20996 14396
rect 20717 14359 20775 14365
rect 20984 14359 20996 14368
rect 20990 14356 20996 14359
rect 21048 14356 21054 14408
rect 24854 14405 24860 14408
rect 24848 14396 24860 14405
rect 24815 14368 24860 14396
rect 24848 14359 24860 14368
rect 24854 14356 24860 14359
rect 24912 14356 24918 14408
rect 26418 14396 26424 14408
rect 26331 14368 26424 14396
rect 26418 14356 26424 14368
rect 26476 14396 26482 14408
rect 26970 14396 26976 14408
rect 26476 14368 26976 14396
rect 26476 14356 26482 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 28276 14405 28304 14572
rect 33226 14560 33232 14572
rect 33284 14560 33290 14612
rect 31389 14467 31447 14473
rect 31389 14433 31401 14467
rect 31435 14464 31447 14467
rect 31754 14464 31760 14476
rect 31435 14436 31760 14464
rect 31435 14433 31447 14436
rect 31389 14427 31447 14433
rect 31754 14424 31760 14436
rect 31812 14424 31818 14476
rect 31849 14467 31907 14473
rect 31849 14433 31861 14467
rect 31895 14464 31907 14467
rect 32306 14464 32312 14476
rect 31895 14436 32312 14464
rect 31895 14433 31907 14436
rect 31849 14427 31907 14433
rect 32306 14424 32312 14436
rect 32364 14424 32370 14476
rect 28261 14399 28319 14405
rect 28261 14365 28273 14399
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28537 14399 28595 14405
rect 28537 14365 28549 14399
rect 28583 14396 28595 14399
rect 28810 14396 28816 14408
rect 28583 14368 28816 14396
rect 28583 14365 28595 14368
rect 28537 14359 28595 14365
rect 28810 14356 28816 14368
rect 28868 14356 28874 14408
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 31113 14399 31171 14405
rect 31113 14396 31125 14399
rect 30156 14368 31125 14396
rect 30156 14356 30162 14368
rect 31113 14365 31125 14368
rect 31159 14365 31171 14399
rect 32122 14396 32128 14408
rect 32083 14368 32128 14396
rect 31113 14359 31171 14365
rect 32122 14356 32128 14368
rect 32180 14356 32186 14408
rect 22094 14328 22100 14340
rect 19628 14300 22100 14328
rect 19429 14291 19487 14297
rect 22094 14288 22100 14300
rect 22152 14288 22158 14340
rect 22186 14288 22192 14340
rect 22244 14328 22250 14340
rect 23382 14328 23388 14340
rect 22244 14300 23388 14328
rect 22244 14288 22250 14300
rect 23382 14288 23388 14300
rect 23440 14328 23446 14340
rect 26688 14331 26746 14337
rect 23440 14300 24900 14328
rect 23440 14288 23446 14300
rect 8168 14232 9536 14260
rect 9677 14263 9735 14269
rect 8168 14220 8174 14232
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 10226 14260 10232 14272
rect 9723 14232 10232 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 19610 14260 19616 14272
rect 19571 14232 19616 14260
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 19794 14260 19800 14272
rect 19755 14232 19800 14260
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 21174 14220 21180 14272
rect 21232 14260 21238 14272
rect 24762 14260 24768 14272
rect 21232 14232 24768 14260
rect 21232 14220 21238 14232
rect 24762 14220 24768 14232
rect 24820 14220 24826 14272
rect 24872 14260 24900 14300
rect 26688 14297 26700 14331
rect 26734 14328 26746 14331
rect 28721 14331 28779 14337
rect 28721 14328 28733 14331
rect 26734 14300 28733 14328
rect 26734 14297 26746 14300
rect 26688 14291 26746 14297
rect 28721 14297 28733 14300
rect 28767 14297 28779 14331
rect 28721 14291 28779 14297
rect 28994 14288 29000 14340
rect 29052 14328 29058 14340
rect 29733 14331 29791 14337
rect 29733 14328 29745 14331
rect 29052 14300 29745 14328
rect 29052 14288 29058 14300
rect 29733 14297 29745 14300
rect 29779 14297 29791 14331
rect 29733 14291 29791 14297
rect 25590 14260 25596 14272
rect 24872 14232 25596 14260
rect 25590 14220 25596 14232
rect 25648 14260 25654 14272
rect 27522 14260 27528 14272
rect 25648 14232 27528 14260
rect 25648 14220 25654 14232
rect 27522 14220 27528 14232
rect 27580 14220 27586 14272
rect 27614 14220 27620 14272
rect 27672 14260 27678 14272
rect 27801 14263 27859 14269
rect 27801 14260 27813 14263
rect 27672 14232 27813 14260
rect 27672 14220 27678 14232
rect 27801 14229 27813 14232
rect 27847 14260 27859 14263
rect 28353 14263 28411 14269
rect 28353 14260 28365 14263
rect 27847 14232 28365 14260
rect 27847 14229 27859 14232
rect 27801 14223 27859 14229
rect 28353 14229 28365 14232
rect 28399 14229 28411 14263
rect 28353 14223 28411 14229
rect 31938 14220 31944 14272
rect 31996 14260 32002 14272
rect 32766 14260 32772 14272
rect 31996 14232 32772 14260
rect 31996 14220 32002 14232
rect 32766 14220 32772 14232
rect 32824 14220 32830 14272
rect 1104 14170 35027 14192
rect 1104 14118 9390 14170
rect 9442 14118 9454 14170
rect 9506 14118 9518 14170
rect 9570 14118 9582 14170
rect 9634 14118 9646 14170
rect 9698 14118 17831 14170
rect 17883 14118 17895 14170
rect 17947 14118 17959 14170
rect 18011 14118 18023 14170
rect 18075 14118 18087 14170
rect 18139 14118 26272 14170
rect 26324 14118 26336 14170
rect 26388 14118 26400 14170
rect 26452 14118 26464 14170
rect 26516 14118 26528 14170
rect 26580 14118 34713 14170
rect 34765 14118 34777 14170
rect 34829 14118 34841 14170
rect 34893 14118 34905 14170
rect 34957 14118 34969 14170
rect 35021 14118 35027 14170
rect 1104 14096 35027 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 1728 14028 2605 14056
rect 1728 14016 1734 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3694 14056 3700 14068
rect 3016 14028 3700 14056
rect 3016 14016 3022 14028
rect 3694 14016 3700 14028
rect 3752 14056 3758 14068
rect 5905 14059 5963 14065
rect 3752 14028 5764 14056
rect 3752 14016 3758 14028
rect 4430 13988 4436 14000
rect 4391 13960 4436 13988
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3050 13920 3056 13932
rect 2731 13892 3056 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3050 13880 3056 13892
rect 3108 13920 3114 13932
rect 3602 13920 3608 13932
rect 3108 13892 3608 13920
rect 3108 13880 3114 13892
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 5736 13920 5764 14028
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 7926 14056 7932 14068
rect 5951 14028 7932 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9950 14056 9956 14068
rect 8260 14028 9956 14056
rect 8260 14016 8266 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 12434 14056 12440 14068
rect 11164 14028 12440 14056
rect 6362 13948 6368 14000
rect 6420 13988 6426 14000
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6420 13960 6561 13988
rect 6420 13948 6426 13960
rect 6549 13957 6561 13960
rect 6595 13988 6607 13991
rect 6638 13988 6644 14000
rect 6595 13960 6644 13988
rect 6595 13957 6607 13960
rect 6549 13951 6607 13957
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 6733 13991 6791 13997
rect 6733 13957 6745 13991
rect 6779 13988 6791 13991
rect 7466 13988 7472 14000
rect 6779 13960 7472 13988
rect 6779 13957 6791 13960
rect 6733 13951 6791 13957
rect 6748 13920 6776 13951
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 11054 13988 11060 14000
rect 9600 13960 11060 13988
rect 5736 13892 6776 13920
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 8386 13920 8392 13932
rect 7055 13892 8392 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 9600 13929 9628 13960
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13889 9643 13923
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9585 13883 9643 13889
rect 9692 13892 9781 13920
rect 4154 13852 4160 13864
rect 4115 13824 4160 13852
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 9692 13852 9720 13892
rect 9769 13889 9781 13892
rect 9815 13920 9827 13923
rect 11164 13920 11192 14028
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 12860 14028 14412 14056
rect 12860 14016 12866 14028
rect 11974 13948 11980 14000
rect 12032 13988 12038 14000
rect 12069 13991 12127 13997
rect 12069 13988 12081 13991
rect 12032 13960 12081 13988
rect 12032 13948 12038 13960
rect 12069 13957 12081 13960
rect 12115 13957 12127 13991
rect 12069 13951 12127 13957
rect 13078 13948 13084 14000
rect 13136 13948 13142 14000
rect 9815 13892 11192 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14384 13929 14412 14028
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 20162 14056 20168 14068
rect 17000 14028 20168 14056
rect 17000 14016 17006 14028
rect 17604 13997 17632 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 22005 14059 22063 14065
rect 22005 14056 22017 14059
rect 20680 14028 22017 14056
rect 20680 14016 20686 14028
rect 22005 14025 22017 14028
rect 22051 14025 22063 14059
rect 28994 14056 29000 14068
rect 22005 14019 22063 14025
rect 27724 14028 29000 14056
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13957 17647 13991
rect 17589 13951 17647 13957
rect 19061 13991 19119 13997
rect 19061 13957 19073 13991
rect 19107 13988 19119 13991
rect 19426 13988 19432 14000
rect 19107 13960 19432 13988
rect 19107 13957 19119 13960
rect 19061 13951 19119 13957
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 19972 13991 20030 13997
rect 19972 13957 19984 13991
rect 20018 13988 20030 13991
rect 20438 13988 20444 14000
rect 20018 13960 20444 13988
rect 20018 13957 20030 13960
rect 19972 13951 20030 13957
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 22281 13991 22339 13997
rect 22281 13957 22293 13991
rect 22327 13988 22339 13991
rect 24026 13988 24032 14000
rect 22327 13960 24032 13988
rect 22327 13957 22339 13960
rect 22281 13951 22339 13957
rect 24026 13948 24032 13960
rect 24084 13988 24090 14000
rect 24673 13991 24731 13997
rect 24673 13988 24685 13991
rect 24084 13960 24685 13988
rect 24084 13948 24090 13960
rect 24673 13957 24685 13960
rect 24719 13957 24731 13991
rect 24673 13951 24731 13957
rect 24762 13948 24768 14000
rect 24820 13988 24826 14000
rect 27479 13991 27537 13997
rect 27479 13988 27491 13991
rect 24820 13960 27491 13988
rect 24820 13948 24826 13960
rect 27479 13957 27491 13960
rect 27525 13957 27537 13991
rect 27479 13951 27537 13957
rect 27617 13991 27675 13997
rect 27617 13957 27629 13991
rect 27663 13988 27675 13991
rect 27724 13988 27752 14028
rect 28994 14016 29000 14028
rect 29052 14016 29058 14068
rect 29089 14059 29147 14065
rect 29089 14025 29101 14059
rect 29135 14056 29147 14059
rect 29914 14056 29920 14068
rect 29135 14028 29920 14056
rect 29135 14025 29147 14028
rect 29089 14019 29147 14025
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 30098 14056 30104 14068
rect 30059 14028 30104 14056
rect 30098 14016 30104 14028
rect 30156 14016 30162 14068
rect 31389 14059 31447 14065
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 31938 14056 31944 14068
rect 31435 14028 31944 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 31938 14016 31944 14028
rect 31996 14016 32002 14068
rect 32030 14016 32036 14068
rect 32088 14056 32094 14068
rect 33686 14056 33692 14068
rect 32088 14028 33692 14056
rect 32088 14016 32094 14028
rect 33686 14016 33692 14028
rect 33744 14016 33750 14068
rect 28718 13988 28724 14000
rect 27663 13960 27752 13988
rect 28679 13960 28724 13988
rect 27663 13957 27675 13960
rect 27617 13951 27675 13957
rect 28718 13948 28724 13960
rect 28776 13948 28782 14000
rect 28902 13988 28908 14000
rect 28863 13960 28908 13988
rect 28902 13948 28908 13960
rect 28960 13948 28966 14000
rect 29012 13988 29040 14016
rect 29733 13991 29791 13997
rect 29733 13988 29745 13991
rect 29012 13960 29745 13988
rect 29733 13957 29745 13960
rect 29779 13957 29791 13991
rect 29733 13951 29791 13957
rect 31220 13960 31616 13988
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13780 13892 14197 13920
rect 13780 13880 13786 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 15378 13920 15384 13932
rect 15339 13892 15384 13920
rect 14369 13883 14427 13889
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 16850 13920 16856 13932
rect 16811 13892 16856 13920
rect 16301 13883 16359 13889
rect 9858 13852 9864 13864
rect 5132 13824 9720 13852
rect 9819 13824 9864 13852
rect 5132 13812 5138 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 11790 13852 11796 13864
rect 11751 13824 11796 13852
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 13262 13812 13268 13864
rect 13320 13852 13326 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13320 13824 13553 13852
rect 13320 13812 13326 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 14090 13852 14096 13864
rect 14051 13824 14096 13852
rect 13541 13815 13599 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 16316 13852 16344 13883
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17678 13920 17684 13932
rect 17359 13892 17684 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 15252 13824 16344 13852
rect 15252 13812 15258 13824
rect 16025 13787 16083 13793
rect 16025 13753 16037 13787
rect 16071 13784 16083 13787
rect 17328 13784 17356 13883
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 18782 13920 18788 13932
rect 18743 13892 18788 13920
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 19702 13920 19708 13932
rect 19663 13892 19708 13920
rect 19702 13880 19708 13892
rect 19760 13880 19766 13932
rect 22186 13920 22192 13932
rect 22147 13892 22192 13920
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22373 13923 22431 13929
rect 22373 13889 22385 13923
rect 22419 13920 22431 13923
rect 22462 13920 22468 13932
rect 22419 13892 22468 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 24578 13920 24584 13932
rect 24539 13892 24584 13920
rect 22557 13883 22615 13889
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 22572 13852 22600 13883
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13920 24915 13923
rect 25038 13920 25044 13932
rect 24903 13892 25044 13920
rect 24903 13889 24915 13892
rect 24857 13883 24915 13889
rect 25038 13880 25044 13892
rect 25096 13920 25102 13932
rect 27706 13920 27712 13932
rect 25096 13892 27476 13920
rect 27667 13892 27712 13920
rect 25096 13880 25102 13892
rect 20864 13824 22600 13852
rect 24596 13852 24624 13880
rect 26602 13852 26608 13864
rect 24596 13824 26608 13852
rect 20864 13812 20870 13824
rect 21100 13793 21128 13824
rect 26602 13812 26608 13824
rect 26660 13812 26666 13864
rect 27338 13852 27344 13864
rect 27299 13824 27344 13852
rect 27338 13812 27344 13824
rect 27396 13812 27402 13864
rect 27448 13852 27476 13892
rect 27706 13880 27712 13892
rect 27764 13880 27770 13932
rect 27798 13880 27804 13932
rect 27856 13920 27862 13932
rect 29638 13920 29644 13932
rect 27856 13892 27901 13920
rect 29599 13892 29644 13920
rect 27856 13880 27862 13892
rect 29638 13880 29644 13892
rect 29696 13880 29702 13932
rect 29917 13923 29975 13929
rect 29917 13889 29929 13923
rect 29963 13920 29975 13923
rect 30374 13920 30380 13932
rect 29963 13892 30380 13920
rect 29963 13889 29975 13892
rect 29917 13883 29975 13889
rect 30374 13880 30380 13892
rect 30432 13880 30438 13932
rect 27985 13855 28043 13861
rect 27448 13824 27660 13852
rect 16071 13756 17356 13784
rect 21085 13787 21143 13793
rect 16071 13753 16083 13756
rect 16025 13747 16083 13753
rect 21085 13753 21097 13787
rect 21131 13753 21143 13787
rect 21085 13747 21143 13753
rect 25041 13787 25099 13793
rect 25041 13753 25053 13787
rect 25087 13784 25099 13787
rect 25130 13784 25136 13796
rect 25087 13756 25136 13784
rect 25087 13753 25099 13756
rect 25041 13747 25099 13753
rect 25130 13744 25136 13756
rect 25188 13744 25194 13796
rect 6733 13719 6791 13725
rect 6733 13685 6745 13719
rect 6779 13716 6791 13719
rect 6822 13716 6828 13728
rect 6779 13688 6828 13716
rect 6779 13685 6791 13688
rect 6733 13679 6791 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 27632 13716 27660 13824
rect 27985 13821 27997 13855
rect 28031 13852 28043 13855
rect 28626 13852 28632 13864
rect 28031 13824 28632 13852
rect 28031 13821 28043 13824
rect 27985 13815 28043 13821
rect 28626 13812 28632 13824
rect 28684 13812 28690 13864
rect 31220 13852 31248 13960
rect 31588 13929 31616 13960
rect 31772 13960 32260 13988
rect 31772 13929 31800 13960
rect 31573 13923 31631 13929
rect 31313 13913 31371 13919
rect 31313 13879 31325 13913
rect 31359 13910 31371 13913
rect 31359 13882 31432 13910
rect 31573 13889 31585 13923
rect 31619 13889 31631 13923
rect 31573 13883 31631 13889
rect 31757 13923 31815 13929
rect 31757 13889 31769 13923
rect 31803 13889 31815 13923
rect 32232 13920 32260 13960
rect 32585 13923 32643 13929
rect 32585 13920 32597 13923
rect 32232 13892 32597 13920
rect 31757 13883 31815 13889
rect 32585 13889 32597 13892
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 31359 13879 31371 13882
rect 31313 13873 31371 13879
rect 28828 13824 31248 13852
rect 28828 13784 28856 13824
rect 28736 13756 28856 13784
rect 28736 13716 28764 13756
rect 28902 13716 28908 13728
rect 27632 13688 28764 13716
rect 28863 13688 28908 13716
rect 28902 13676 28908 13688
rect 28960 13676 28966 13728
rect 29638 13676 29644 13728
rect 29696 13716 29702 13728
rect 31404 13716 31432 13882
rect 31588 13852 31616 13883
rect 32030 13852 32036 13864
rect 31588 13824 32036 13852
rect 32030 13812 32036 13824
rect 32088 13812 32094 13864
rect 32306 13852 32312 13864
rect 32267 13824 32312 13852
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 32766 13812 32772 13864
rect 32824 13852 32830 13864
rect 33689 13855 33747 13861
rect 33689 13852 33701 13855
rect 32824 13824 33701 13852
rect 32824 13812 32830 13824
rect 33689 13821 33701 13824
rect 33735 13821 33747 13855
rect 33689 13815 33747 13821
rect 33410 13716 33416 13728
rect 29696 13688 33416 13716
rect 29696 13676 29702 13688
rect 33410 13676 33416 13688
rect 33468 13676 33474 13728
rect 1104 13626 34868 13648
rect 1104 13574 5170 13626
rect 5222 13574 5234 13626
rect 5286 13574 5298 13626
rect 5350 13574 5362 13626
rect 5414 13574 5426 13626
rect 5478 13574 13611 13626
rect 13663 13574 13675 13626
rect 13727 13574 13739 13626
rect 13791 13574 13803 13626
rect 13855 13574 13867 13626
rect 13919 13574 22052 13626
rect 22104 13574 22116 13626
rect 22168 13574 22180 13626
rect 22232 13574 22244 13626
rect 22296 13574 22308 13626
rect 22360 13574 30493 13626
rect 30545 13574 30557 13626
rect 30609 13574 30621 13626
rect 30673 13574 30685 13626
rect 30737 13574 30749 13626
rect 30801 13574 34868 13626
rect 1104 13552 34868 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4154 13512 4160 13524
rect 3467 13484 4160 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 5534 13512 5540 13524
rect 5495 13484 5540 13512
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 10502 13512 10508 13524
rect 5644 13484 10508 13512
rect 4246 13444 4252 13456
rect 2976 13416 4252 13444
rect 2976 13385 3004 13416
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 5644 13444 5672 13484
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 15378 13512 15384 13524
rect 10888 13484 15384 13512
rect 4632 13416 5672 13444
rect 2961 13379 3019 13385
rect 2961 13376 2973 13379
rect 2516 13348 2973 13376
rect 2516 13317 2544 13348
rect 2961 13345 2973 13348
rect 3007 13345 3019 13379
rect 2961 13339 3019 13345
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3878 13308 3884 13320
rect 3283 13280 3884 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 2332 13240 2360 13271
rect 3068 13240 3096 13271
rect 3878 13268 3884 13280
rect 3936 13268 3942 13320
rect 4632 13317 4660 13416
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 8352 13416 9168 13444
rect 8352 13404 8358 13416
rect 9140 13388 9168 13416
rect 9122 13376 9128 13388
rect 5552 13348 8432 13376
rect 9035 13348 9128 13376
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5132 13280 5365 13308
rect 5132 13268 5138 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 3970 13240 3976 13252
rect 2332 13212 3976 13240
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4062 13200 4068 13252
rect 4120 13240 4126 13252
rect 4249 13243 4307 13249
rect 4249 13240 4261 13243
rect 4120 13212 4261 13240
rect 4120 13200 4126 13212
rect 4249 13209 4261 13212
rect 4295 13240 4307 13243
rect 5552 13240 5580 13348
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13308 5687 13311
rect 8294 13308 8300 13320
rect 5675 13280 8300 13308
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 4295 13212 5580 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 5644 13172 5672 13271
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 8404 13317 8432 13348
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8573 13243 8631 13249
rect 8573 13209 8585 13243
rect 8619 13240 8631 13243
rect 8662 13240 8668 13252
rect 8619 13212 8668 13240
rect 8619 13209 8631 13212
rect 8573 13203 8631 13209
rect 8662 13200 8668 13212
rect 8720 13200 8726 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 8772 13212 9413 13240
rect 3200 13144 5672 13172
rect 3200 13132 3206 13144
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8478 13172 8484 13184
rect 7524 13144 8484 13172
rect 7524 13132 7530 13144
rect 8478 13132 8484 13144
rect 8536 13172 8542 13184
rect 8772 13172 8800 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 9858 13200 9864 13252
rect 9916 13200 9922 13252
rect 8536 13144 8800 13172
rect 8536 13132 8542 13144
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 10888 13181 10916 13484
rect 15378 13472 15384 13484
rect 15436 13512 15442 13524
rect 15654 13512 15660 13524
rect 15436 13484 15516 13512
rect 15615 13484 15660 13512
rect 15436 13472 15442 13484
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11514 13376 11520 13388
rect 11204 13348 11520 13376
rect 11204 13336 11210 13348
rect 11514 13336 11520 13348
rect 11572 13376 11578 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11572 13348 12081 13376
rect 11572 13336 11578 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13136 13348 13553 13376
rect 13136 13336 13142 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 13556 13308 13584 13339
rect 15102 13308 15108 13320
rect 13556 13280 15108 13308
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 15488 13317 15516 13484
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 26970 13472 26976 13524
rect 27028 13512 27034 13524
rect 27341 13515 27399 13521
rect 27341 13512 27353 13515
rect 27028 13484 27353 13512
rect 27028 13472 27034 13484
rect 27341 13481 27353 13484
rect 27387 13481 27399 13515
rect 27341 13475 27399 13481
rect 31665 13515 31723 13521
rect 31665 13481 31677 13515
rect 31711 13512 31723 13515
rect 32306 13512 32312 13524
rect 31711 13484 32312 13512
rect 31711 13481 31723 13484
rect 31665 13475 31723 13481
rect 32306 13472 32312 13484
rect 32364 13472 32370 13524
rect 18322 13404 18328 13456
rect 18380 13404 18386 13456
rect 18340 13376 18368 13404
rect 18509 13379 18567 13385
rect 18064 13348 18460 13376
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13308 15531 13311
rect 15746 13308 15752 13320
rect 15519 13280 15752 13308
rect 15519 13277 15531 13280
rect 15473 13271 15531 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16390 13308 16396 13320
rect 16351 13280 16396 13308
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 18064 13317 18092 13348
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18322 13308 18328 13320
rect 18283 13280 18328 13308
rect 18049 13271 18107 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 14090 13240 14096 13252
rect 13294 13212 14096 13240
rect 14090 13200 14096 13212
rect 14148 13200 14154 13252
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15620 13212 16221 13240
rect 15620 13200 15626 13212
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 16761 13243 16819 13249
rect 16761 13209 16773 13243
rect 16807 13240 16819 13243
rect 16850 13240 16856 13252
rect 16807 13212 16856 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 16850 13200 16856 13212
rect 16908 13240 16914 13252
rect 17494 13240 17500 13252
rect 16908 13212 17500 13240
rect 16908 13200 16914 13212
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18432 13240 18460 13348
rect 18509 13345 18521 13379
rect 18555 13376 18567 13379
rect 20530 13376 20536 13388
rect 18555 13348 20536 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 20530 13336 20536 13348
rect 20588 13376 20594 13388
rect 22370 13376 22376 13388
rect 20588 13348 22376 13376
rect 20588 13336 20594 13348
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 20257 13311 20315 13317
rect 20257 13308 20269 13311
rect 19852 13280 20269 13308
rect 19852 13268 19858 13280
rect 20257 13277 20269 13280
rect 20303 13277 20315 13311
rect 26050 13308 26056 13320
rect 26011 13280 26056 13308
rect 20257 13271 20315 13277
rect 26050 13268 26056 13280
rect 26108 13268 26114 13320
rect 32953 13311 33011 13317
rect 32953 13277 32965 13311
rect 32999 13308 33011 13311
rect 33594 13308 33600 13320
rect 32999 13280 33600 13308
rect 32999 13277 33011 13280
rect 32953 13271 33011 13277
rect 33594 13268 33600 13280
rect 33652 13268 33658 13320
rect 18506 13240 18512 13252
rect 18432 13212 18512 13240
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 9088 13144 10885 13172
rect 9088 13132 9094 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 18230 13132 18236 13184
rect 18288 13172 18294 13184
rect 21545 13175 21603 13181
rect 21545 13172 21557 13175
rect 18288 13144 21557 13172
rect 18288 13132 18294 13144
rect 21545 13141 21557 13144
rect 21591 13141 21603 13175
rect 21545 13135 21603 13141
rect 1104 13082 35027 13104
rect 1104 13030 9390 13082
rect 9442 13030 9454 13082
rect 9506 13030 9518 13082
rect 9570 13030 9582 13082
rect 9634 13030 9646 13082
rect 9698 13030 17831 13082
rect 17883 13030 17895 13082
rect 17947 13030 17959 13082
rect 18011 13030 18023 13082
rect 18075 13030 18087 13082
rect 18139 13030 26272 13082
rect 26324 13030 26336 13082
rect 26388 13030 26400 13082
rect 26452 13030 26464 13082
rect 26516 13030 26528 13082
rect 26580 13030 34713 13082
rect 34765 13030 34777 13082
rect 34829 13030 34841 13082
rect 34893 13030 34905 13082
rect 34957 13030 34969 13082
rect 35021 13030 35027 13082
rect 1104 13008 35027 13030
rect 3878 12968 3884 12980
rect 3839 12940 3884 12968
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 4028 12940 4353 12968
rect 4028 12928 4034 12940
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 4341 12931 4399 12937
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 11790 12968 11796 12980
rect 9180 12940 11796 12968
rect 9180 12928 9186 12940
rect 2406 12900 2412 12912
rect 2367 12872 2412 12900
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 3050 12860 3056 12912
rect 3108 12860 3114 12912
rect 8662 12860 8668 12912
rect 8720 12860 8726 12912
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 9401 12903 9459 12909
rect 9401 12900 9413 12903
rect 9364 12872 9413 12900
rect 9364 12860 9370 12872
rect 9401 12869 9413 12872
rect 9447 12869 9459 12903
rect 9401 12863 9459 12869
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12801 2191 12835
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 2133 12795 2191 12801
rect 3620 12804 4353 12832
rect 2148 12764 2176 12795
rect 3620 12776 3648 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4522 12832 4528 12844
rect 4483 12804 4528 12832
rect 4341 12795 4399 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 9692 12841 9720 12940
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 22922 12968 22928 12980
rect 17644 12940 22416 12968
rect 22883 12940 22928 12968
rect 17644 12928 17650 12940
rect 12986 12900 12992 12912
rect 12947 12872 12992 12900
rect 12986 12860 12992 12872
rect 13044 12860 13050 12912
rect 14734 12900 14740 12912
rect 14695 12872 14740 12900
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 18322 12900 18328 12912
rect 18064 12872 18328 12900
rect 18064 12844 18092 12872
rect 18322 12860 18328 12872
rect 18380 12900 18386 12912
rect 19153 12903 19211 12909
rect 18380 12872 19012 12900
rect 18380 12860 18386 12872
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15252 12804 15393 12832
rect 15252 12792 15258 12804
rect 15381 12801 15393 12804
rect 15427 12832 15439 12835
rect 15562 12832 15568 12844
rect 15427 12804 15568 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16390 12832 16396 12844
rect 16071 12804 16396 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 3142 12764 3148 12776
rect 2148 12736 3148 12764
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 3602 12724 3608 12776
rect 3660 12724 3666 12776
rect 16040 12764 16068 12795
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 18046 12832 18052 12844
rect 18007 12804 18052 12832
rect 17589 12795 17647 12801
rect 14568 12736 16068 12764
rect 16117 12767 16175 12773
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 13170 12696 13176 12708
rect 10560 12668 13176 12696
rect 10560 12656 10566 12668
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 14568 12640 14596 12736
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16574 12764 16580 12776
rect 16163 12736 16580 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16574 12724 16580 12736
rect 16632 12764 16638 12776
rect 17604 12764 17632 12795
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 18690 12832 18696 12844
rect 18472 12804 18696 12832
rect 18472 12792 18478 12804
rect 18690 12792 18696 12804
rect 18748 12832 18754 12844
rect 18984 12841 19012 12872
rect 19153 12869 19165 12903
rect 19199 12900 19211 12903
rect 19610 12900 19616 12912
rect 19199 12872 19616 12900
rect 19199 12869 19211 12872
rect 19153 12863 19211 12869
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 18748 12804 18797 12832
rect 18748 12792 18754 12804
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 19961 12835 20019 12841
rect 19961 12832 19973 12835
rect 19852 12804 19973 12832
rect 19852 12792 19858 12804
rect 19961 12801 19973 12804
rect 20007 12801 20019 12835
rect 22278 12832 22284 12844
rect 22239 12804 22284 12832
rect 19961 12795 20019 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 22388 12841 22416 12940
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 27893 12971 27951 12977
rect 27893 12937 27905 12971
rect 27939 12968 27951 12971
rect 28442 12968 28448 12980
rect 27939 12940 28448 12968
rect 27939 12937 27951 12940
rect 27893 12931 27951 12937
rect 28442 12928 28448 12940
rect 28500 12928 28506 12980
rect 28534 12928 28540 12980
rect 28592 12968 28598 12980
rect 28721 12971 28779 12977
rect 28721 12968 28733 12971
rect 28592 12940 28733 12968
rect 28592 12928 28598 12940
rect 28721 12937 28733 12940
rect 28767 12937 28779 12971
rect 28721 12931 28779 12937
rect 32122 12928 32128 12980
rect 32180 12968 32186 12980
rect 32309 12971 32367 12977
rect 32309 12968 32321 12971
rect 32180 12940 32321 12968
rect 32180 12928 32186 12940
rect 32309 12937 32321 12940
rect 32355 12937 32367 12971
rect 32309 12931 32367 12937
rect 32677 12971 32735 12977
rect 32677 12937 32689 12971
rect 32723 12968 32735 12971
rect 33226 12968 33232 12980
rect 32723 12940 33232 12968
rect 32723 12937 32735 12940
rect 32677 12931 32735 12937
rect 33226 12928 33232 12940
rect 33284 12928 33290 12980
rect 22649 12903 22707 12909
rect 22649 12869 22661 12903
rect 22695 12900 22707 12903
rect 24762 12900 24768 12912
rect 22695 12872 24768 12900
rect 22695 12869 22707 12872
rect 22649 12863 22707 12869
rect 24762 12860 24768 12872
rect 24820 12860 24826 12912
rect 27522 12900 27528 12912
rect 27483 12872 27528 12900
rect 27522 12860 27528 12872
rect 27580 12860 27586 12912
rect 27617 12903 27675 12909
rect 27617 12869 27629 12903
rect 27663 12900 27675 12903
rect 28258 12900 28264 12912
rect 27663 12872 28264 12900
rect 27663 12869 27675 12872
rect 27617 12863 27675 12869
rect 28258 12860 28264 12872
rect 28316 12860 28322 12912
rect 30282 12900 30288 12912
rect 28736 12872 30288 12900
rect 22374 12835 22432 12841
rect 22374 12801 22386 12835
rect 22420 12801 22432 12835
rect 22554 12832 22560 12844
rect 22515 12804 22560 12832
rect 22374 12795 22432 12801
rect 22554 12792 22560 12804
rect 22612 12792 22618 12844
rect 22787 12835 22845 12841
rect 22787 12801 22799 12835
rect 22833 12832 22845 12835
rect 22922 12832 22928 12844
rect 22833 12804 22928 12832
rect 22833 12801 22845 12804
rect 22787 12795 22845 12801
rect 22922 12792 22928 12804
rect 22980 12792 22986 12844
rect 27246 12832 27252 12844
rect 27207 12804 27252 12832
rect 27246 12792 27252 12804
rect 27304 12792 27310 12844
rect 27397 12835 27455 12841
rect 27397 12801 27409 12835
rect 27443 12832 27455 12835
rect 27755 12835 27813 12841
rect 27443 12804 27660 12832
rect 27443 12801 27455 12804
rect 27397 12795 27455 12801
rect 27632 12776 27660 12804
rect 27755 12801 27767 12835
rect 27801 12832 27813 12835
rect 27982 12832 27988 12844
rect 27801 12804 27988 12832
rect 27801 12801 27813 12804
rect 27755 12795 27813 12801
rect 27982 12792 27988 12804
rect 28040 12792 28046 12844
rect 28537 12835 28595 12841
rect 28537 12801 28549 12835
rect 28583 12832 28595 12835
rect 28736 12832 28764 12872
rect 30282 12860 30288 12872
rect 30340 12860 30346 12912
rect 28583 12804 28764 12832
rect 28813 12835 28871 12841
rect 28583 12801 28595 12804
rect 28537 12795 28595 12801
rect 28813 12801 28825 12835
rect 28859 12801 28871 12835
rect 28813 12795 28871 12801
rect 18322 12764 18328 12776
rect 16632 12736 17632 12764
rect 18283 12736 18328 12764
rect 16632 12724 16638 12736
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 7558 12588 7564 12640
rect 7616 12628 7622 12640
rect 7929 12631 7987 12637
rect 7929 12628 7941 12631
rect 7616 12600 7941 12628
rect 7616 12588 7622 12600
rect 7929 12597 7941 12600
rect 7975 12628 7987 12631
rect 14550 12628 14556 12640
rect 7975 12600 14556 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 19720 12628 19748 12727
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 23014 12764 23020 12776
rect 21140 12736 23020 12764
rect 21140 12724 21146 12736
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 27614 12724 27620 12776
rect 27672 12724 27678 12776
rect 28828 12764 28856 12795
rect 29638 12792 29644 12844
rect 29696 12832 29702 12844
rect 29733 12835 29791 12841
rect 29733 12832 29745 12835
rect 29696 12804 29745 12832
rect 29696 12792 29702 12804
rect 29733 12801 29745 12804
rect 29779 12801 29791 12835
rect 32490 12832 32496 12844
rect 32451 12804 32496 12832
rect 29733 12795 29791 12801
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 32769 12835 32827 12841
rect 32769 12801 32781 12835
rect 32815 12832 32827 12835
rect 33410 12832 33416 12844
rect 32815 12804 33416 12832
rect 32815 12801 32827 12804
rect 32769 12795 32827 12801
rect 33410 12792 33416 12804
rect 33468 12792 33474 12844
rect 29549 12767 29607 12773
rect 29549 12764 29561 12767
rect 28828 12736 29561 12764
rect 29549 12733 29561 12736
rect 29595 12764 29607 12767
rect 30190 12764 30196 12776
rect 29595 12736 30196 12764
rect 29595 12733 29607 12736
rect 29549 12727 29607 12733
rect 30190 12724 30196 12736
rect 30248 12724 30254 12776
rect 23290 12696 23296 12708
rect 22066 12668 23296 12696
rect 19978 12628 19984 12640
rect 19720 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 21082 12628 21088 12640
rect 21043 12600 21088 12628
rect 21082 12588 21088 12600
rect 21140 12628 21146 12640
rect 22066 12628 22094 12668
rect 23290 12656 23296 12668
rect 23348 12656 23354 12708
rect 28074 12656 28080 12708
rect 28132 12696 28138 12708
rect 28902 12696 28908 12708
rect 28132 12668 28908 12696
rect 28132 12656 28138 12668
rect 28902 12656 28908 12668
rect 28960 12696 28966 12708
rect 31018 12696 31024 12708
rect 28960 12668 31024 12696
rect 28960 12656 28966 12668
rect 31018 12656 31024 12668
rect 31076 12656 31082 12708
rect 28350 12628 28356 12640
rect 21140 12600 22094 12628
rect 28311 12600 28356 12628
rect 21140 12588 21146 12600
rect 28350 12588 28356 12600
rect 28408 12588 28414 12640
rect 1104 12538 34868 12560
rect 1104 12486 5170 12538
rect 5222 12486 5234 12538
rect 5286 12486 5298 12538
rect 5350 12486 5362 12538
rect 5414 12486 5426 12538
rect 5478 12486 13611 12538
rect 13663 12486 13675 12538
rect 13727 12486 13739 12538
rect 13791 12486 13803 12538
rect 13855 12486 13867 12538
rect 13919 12486 22052 12538
rect 22104 12486 22116 12538
rect 22168 12486 22180 12538
rect 22232 12486 22244 12538
rect 22296 12486 22308 12538
rect 22360 12486 30493 12538
rect 30545 12486 30557 12538
rect 30609 12486 30621 12538
rect 30673 12486 30685 12538
rect 30737 12486 30749 12538
rect 30801 12486 34868 12538
rect 1104 12464 34868 12486
rect 3050 12424 3056 12436
rect 3011 12396 3056 12424
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 19794 12384 19800 12436
rect 19852 12424 19858 12436
rect 19889 12427 19947 12433
rect 19889 12424 19901 12427
rect 19852 12396 19901 12424
rect 19852 12384 19858 12396
rect 19889 12393 19901 12396
rect 19935 12393 19947 12427
rect 19889 12387 19947 12393
rect 20254 12384 20260 12436
rect 20312 12424 20318 12436
rect 20806 12424 20812 12436
rect 20312 12396 20812 12424
rect 20312 12384 20318 12396
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 21910 12384 21916 12436
rect 21968 12424 21974 12436
rect 22097 12427 22155 12433
rect 22097 12424 22109 12427
rect 21968 12396 22109 12424
rect 21968 12384 21974 12396
rect 22097 12393 22109 12396
rect 22143 12424 22155 12427
rect 22738 12424 22744 12436
rect 22143 12396 22744 12424
rect 22143 12393 22155 12396
rect 22097 12387 22155 12393
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 23014 12424 23020 12436
rect 22975 12396 23020 12424
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 23382 12384 23388 12436
rect 23440 12424 23446 12436
rect 24854 12424 24860 12436
rect 23440 12396 24860 12424
rect 23440 12384 23446 12396
rect 24854 12384 24860 12396
rect 24912 12424 24918 12436
rect 24912 12396 28856 12424
rect 24912 12384 24918 12396
rect 28828 12368 28856 12396
rect 18322 12316 18328 12368
rect 18380 12356 18386 12368
rect 23106 12356 23112 12368
rect 18380 12328 23112 12356
rect 18380 12316 18386 12328
rect 23106 12316 23112 12328
rect 23164 12356 23170 12368
rect 23164 12328 27016 12356
rect 23164 12316 23170 12328
rect 16669 12291 16727 12297
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 18046 12288 18052 12300
rect 16715 12260 18052 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12220 3203 12223
rect 4062 12220 4068 12232
rect 3191 12192 4068 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 2958 12112 2964 12164
rect 3016 12152 3022 12164
rect 3160 12152 3188 12183
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 14550 12220 14556 12232
rect 14511 12192 14556 12220
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 15194 12220 15200 12232
rect 15155 12192 15200 12220
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15804 12192 15945 12220
rect 15804 12180 15810 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16540 12192 16589 12220
rect 16540 12180 16546 12192
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 17494 12220 17500 12232
rect 17455 12192 17500 12220
rect 16577 12183 16635 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17972 12229 18000 12260
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 21082 12288 21088 12300
rect 19536 12260 21088 12288
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18782 12220 18788 12232
rect 18279 12192 18788 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 18782 12180 18788 12192
rect 18840 12180 18846 12232
rect 19536 12229 19564 12260
rect 21082 12248 21088 12260
rect 21140 12248 21146 12300
rect 22066 12260 23612 12288
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 3016 12124 3188 12152
rect 15013 12155 15071 12161
rect 3016 12112 3022 12124
rect 15013 12121 15025 12155
rect 15059 12152 15071 12155
rect 16942 12152 16948 12164
rect 15059 12124 16948 12152
rect 15059 12121 15071 12124
rect 15013 12115 15071 12121
rect 16942 12112 16948 12124
rect 17000 12152 17006 12164
rect 18690 12152 18696 12164
rect 17000 12124 18696 12152
rect 17000 12112 17006 12124
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 19444 12152 19472 12183
rect 19610 12180 19616 12232
rect 19668 12220 19674 12232
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19668 12192 19717 12220
rect 19668 12180 19674 12192
rect 19705 12189 19717 12192
rect 19751 12220 19763 12223
rect 20346 12220 20352 12232
rect 19751 12192 20352 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 22066 12220 22094 12260
rect 20588 12192 22094 12220
rect 20588 12180 20594 12192
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 22520 12192 23213 12220
rect 22520 12180 22526 12192
rect 23201 12189 23213 12192
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 23290 12180 23296 12232
rect 23348 12220 23354 12232
rect 23584 12229 23612 12260
rect 24670 12248 24676 12300
rect 24728 12288 24734 12300
rect 24728 12260 25084 12288
rect 24728 12248 24734 12260
rect 23477 12223 23535 12229
rect 23348 12192 23393 12220
rect 23348 12180 23354 12192
rect 23477 12189 23489 12223
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 24854 12220 24860 12232
rect 24811 12192 24860 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 20254 12152 20260 12164
rect 19444 12124 20260 12152
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 20714 12112 20720 12164
rect 20772 12152 20778 12164
rect 20809 12155 20867 12161
rect 20809 12152 20821 12155
rect 20772 12124 20821 12152
rect 20772 12112 20778 12124
rect 20809 12121 20821 12124
rect 20855 12121 20867 12155
rect 20809 12115 20867 12121
rect 21266 12112 21272 12164
rect 21324 12152 21330 12164
rect 22094 12152 22100 12164
rect 21324 12124 22100 12152
rect 21324 12112 21330 12124
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 22186 12112 22192 12164
rect 22244 12152 22250 12164
rect 22922 12152 22928 12164
rect 22244 12124 22928 12152
rect 22244 12112 22250 12124
rect 22922 12112 22928 12124
rect 22980 12112 22986 12164
rect 23492 12152 23520 12183
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 25056 12229 25084 12260
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12189 25099 12223
rect 26988 12220 27016 12328
rect 28810 12316 28816 12368
rect 28868 12356 28874 12368
rect 32122 12356 32128 12368
rect 28868 12328 32128 12356
rect 28868 12316 28874 12328
rect 32122 12316 32128 12328
rect 32180 12316 32186 12368
rect 27798 12220 27804 12232
rect 26988 12192 27804 12220
rect 25041 12183 25099 12189
rect 27798 12180 27804 12192
rect 27856 12220 27862 12232
rect 28123 12223 28181 12229
rect 28123 12220 28135 12223
rect 27856 12192 28135 12220
rect 27856 12180 27862 12192
rect 28123 12189 28135 12192
rect 28169 12189 28181 12223
rect 28534 12220 28540 12232
rect 28495 12192 28540 12220
rect 28123 12183 28181 12189
rect 28534 12180 28540 12192
rect 28592 12180 28598 12232
rect 28626 12180 28632 12232
rect 28684 12220 28690 12232
rect 28684 12192 28729 12220
rect 28684 12180 28690 12192
rect 28261 12155 28319 12161
rect 23492 12124 28028 12152
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 22646 12084 22652 12096
rect 20220 12056 22652 12084
rect 20220 12044 20226 12056
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 24578 12084 24584 12096
rect 24539 12056 24584 12084
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 24762 12044 24768 12096
rect 24820 12084 24826 12096
rect 28000 12093 28028 12124
rect 28261 12121 28273 12155
rect 28307 12121 28319 12155
rect 28261 12115 28319 12121
rect 28353 12155 28411 12161
rect 28353 12121 28365 12155
rect 28399 12152 28411 12155
rect 28442 12152 28448 12164
rect 28399 12124 28448 12152
rect 28399 12121 28411 12124
rect 28353 12115 28411 12121
rect 24949 12087 25007 12093
rect 24949 12084 24961 12087
rect 24820 12056 24961 12084
rect 24820 12044 24826 12056
rect 24949 12053 24961 12056
rect 24995 12053 25007 12087
rect 24949 12047 25007 12053
rect 27985 12087 28043 12093
rect 27985 12053 27997 12087
rect 28031 12053 28043 12087
rect 28276 12084 28304 12115
rect 28442 12112 28448 12124
rect 28500 12112 28506 12164
rect 31202 12084 31208 12096
rect 28276 12056 31208 12084
rect 27985 12047 28043 12053
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 1104 11994 35027 12016
rect 1104 11942 9390 11994
rect 9442 11942 9454 11994
rect 9506 11942 9518 11994
rect 9570 11942 9582 11994
rect 9634 11942 9646 11994
rect 9698 11942 17831 11994
rect 17883 11942 17895 11994
rect 17947 11942 17959 11994
rect 18011 11942 18023 11994
rect 18075 11942 18087 11994
rect 18139 11942 26272 11994
rect 26324 11942 26336 11994
rect 26388 11942 26400 11994
rect 26452 11942 26464 11994
rect 26516 11942 26528 11994
rect 26580 11942 34713 11994
rect 34765 11942 34777 11994
rect 34829 11942 34841 11994
rect 34893 11942 34905 11994
rect 34957 11942 34969 11994
rect 35021 11942 35027 11994
rect 1104 11920 35027 11942
rect 17129 11883 17187 11889
rect 17129 11849 17141 11883
rect 17175 11880 17187 11883
rect 22186 11880 22192 11892
rect 17175 11852 22192 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 22370 11880 22376 11892
rect 22331 11852 22376 11880
rect 22370 11840 22376 11852
rect 22428 11840 22434 11892
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 22888 11852 24716 11880
rect 22888 11840 22894 11852
rect 15194 11812 15200 11824
rect 14200 11784 15200 11812
rect 13262 11704 13268 11756
rect 13320 11744 13326 11756
rect 14200 11753 14228 11784
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 15746 11812 15752 11824
rect 15707 11784 15752 11812
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 16301 11815 16359 11821
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 16758 11812 16764 11824
rect 16347 11784 16764 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 16758 11772 16764 11784
rect 16816 11812 16822 11824
rect 16816 11784 18184 11812
rect 16816 11772 16822 11784
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13320 11716 14197 11744
rect 13320 11704 13326 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14185 11707 14243 11713
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 14737 11747 14795 11753
rect 14737 11744 14749 11747
rect 14608 11716 14749 11744
rect 14608 11704 14614 11716
rect 14737 11713 14749 11716
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15344 11716 15945 11744
rect 15344 11704 15350 11716
rect 15933 11713 15945 11716
rect 15979 11744 15991 11747
rect 16482 11744 16488 11756
rect 15979 11716 16488 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 17052 11753 17080 11784
rect 18156 11753 18184 11784
rect 22462 11772 22468 11824
rect 22520 11812 22526 11824
rect 22741 11815 22799 11821
rect 22741 11812 22753 11815
rect 22520 11784 22753 11812
rect 22520 11772 22526 11784
rect 22741 11781 22753 11784
rect 22787 11781 22799 11815
rect 22741 11775 22799 11781
rect 24112 11815 24170 11821
rect 24112 11781 24124 11815
rect 24158 11812 24170 11815
rect 24578 11812 24584 11824
rect 24158 11784 24584 11812
rect 24158 11781 24170 11784
rect 24112 11775 24170 11781
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 24688 11812 24716 11852
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 25225 11883 25283 11889
rect 25225 11880 25237 11883
rect 24820 11852 25237 11880
rect 24820 11840 24826 11852
rect 25225 11849 25237 11852
rect 25271 11849 25283 11883
rect 28718 11880 28724 11892
rect 25225 11843 25283 11849
rect 25700 11852 28724 11880
rect 25700 11821 25728 11852
rect 28718 11840 28724 11852
rect 28776 11880 28782 11892
rect 30834 11880 30840 11892
rect 28776 11852 30840 11880
rect 28776 11840 28782 11852
rect 30834 11840 30840 11852
rect 30892 11840 30898 11892
rect 31202 11880 31208 11892
rect 31163 11852 31208 11880
rect 31202 11840 31208 11852
rect 31260 11840 31266 11892
rect 32214 11840 32220 11892
rect 32272 11880 32278 11892
rect 32677 11883 32735 11889
rect 32677 11880 32689 11883
rect 32272 11852 32689 11880
rect 32272 11840 32278 11852
rect 32677 11849 32689 11852
rect 32723 11880 32735 11883
rect 33594 11880 33600 11892
rect 32723 11852 33600 11880
rect 32723 11849 32735 11852
rect 32677 11843 32735 11849
rect 33594 11840 33600 11852
rect 33652 11840 33658 11892
rect 25685 11815 25743 11821
rect 25685 11812 25697 11815
rect 24688 11784 25697 11812
rect 25685 11781 25697 11784
rect 25731 11781 25743 11815
rect 25685 11775 25743 11781
rect 25869 11815 25927 11821
rect 25869 11781 25881 11815
rect 25915 11781 25927 11815
rect 25869 11775 25927 11781
rect 27700 11815 27758 11821
rect 27700 11781 27712 11815
rect 27746 11812 27758 11815
rect 28350 11812 28356 11824
rect 27746 11784 28356 11812
rect 27746 11781 27758 11784
rect 27700 11775 27758 11781
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16632 11716 16865 11744
rect 16632 11704 16638 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 20340 11747 20398 11753
rect 20340 11713 20352 11747
rect 20386 11744 20398 11747
rect 20898 11744 20904 11756
rect 20386 11716 20904 11744
rect 20386 11713 20398 11716
rect 20340 11707 20398 11713
rect 14277 11611 14335 11617
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 17696 11608 17724 11707
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 21082 11704 21088 11756
rect 21140 11744 21146 11756
rect 22554 11744 22560 11756
rect 21140 11716 22560 11744
rect 21140 11704 21146 11716
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 22646 11704 22652 11756
rect 22704 11744 22710 11756
rect 22925 11747 22983 11753
rect 22704 11716 22749 11744
rect 22704 11704 22710 11716
rect 22925 11713 22937 11747
rect 22971 11713 22983 11747
rect 22925 11707 22983 11713
rect 18414 11676 18420 11688
rect 18375 11648 18420 11676
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 20036 11648 20085 11676
rect 20036 11636 20042 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 22940 11676 22968 11707
rect 23014 11704 23020 11756
rect 23072 11744 23078 11756
rect 25884 11744 25912 11775
rect 28350 11772 28356 11784
rect 28408 11772 28414 11824
rect 30374 11772 30380 11824
rect 30432 11812 30438 11824
rect 30432 11784 31432 11812
rect 30432 11772 30438 11784
rect 25958 11744 25964 11756
rect 23072 11716 25964 11744
rect 23072 11704 23078 11716
rect 25958 11704 25964 11716
rect 26016 11704 26022 11756
rect 28074 11744 28080 11756
rect 26068 11716 28080 11744
rect 23842 11676 23848 11688
rect 20073 11639 20131 11645
rect 22066 11648 22968 11676
rect 23803 11648 23848 11676
rect 18506 11608 18512 11620
rect 14323 11580 18512 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 18506 11568 18512 11580
rect 18564 11568 18570 11620
rect 21358 11568 21364 11620
rect 21416 11608 21422 11620
rect 21453 11611 21511 11617
rect 21453 11608 21465 11611
rect 21416 11580 21465 11608
rect 21416 11568 21422 11580
rect 21453 11577 21465 11580
rect 21499 11608 21511 11611
rect 22066 11608 22094 11648
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 26068 11608 26096 11716
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 30190 11704 30196 11756
rect 30248 11744 30254 11756
rect 31404 11753 31432 11784
rect 31113 11747 31171 11753
rect 31113 11744 31125 11747
rect 30248 11716 31125 11744
rect 30248 11704 30254 11716
rect 31113 11713 31125 11716
rect 31159 11713 31171 11747
rect 31113 11707 31171 11713
rect 31389 11747 31447 11753
rect 31389 11713 31401 11747
rect 31435 11713 31447 11747
rect 31389 11707 31447 11713
rect 27433 11679 27491 11685
rect 27433 11645 27445 11679
rect 27479 11645 27491 11679
rect 31128 11676 31156 11707
rect 32122 11704 32128 11756
rect 32180 11744 32186 11756
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 32180 11716 32505 11744
rect 32180 11704 32186 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 32769 11747 32827 11753
rect 32769 11713 32781 11747
rect 32815 11713 32827 11747
rect 32769 11707 32827 11713
rect 32784 11676 32812 11707
rect 33410 11676 33416 11688
rect 31128 11648 33416 11676
rect 27433 11639 27491 11645
rect 21499 11580 22094 11608
rect 25884 11580 26096 11608
rect 21499 11577 21511 11580
rect 21453 11571 21511 11577
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22370 11540 22376 11552
rect 22152 11512 22376 11540
rect 22152 11500 22158 11512
rect 22370 11500 22376 11512
rect 22428 11540 22434 11552
rect 23382 11540 23388 11552
rect 22428 11512 23388 11540
rect 22428 11500 22434 11512
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 25884 11549 25912 11580
rect 25869 11543 25927 11549
rect 25869 11509 25881 11543
rect 25915 11509 25927 11543
rect 26050 11540 26056 11552
rect 26011 11512 26056 11540
rect 25869 11503 25927 11509
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 27448 11540 27476 11639
rect 33410 11636 33416 11648
rect 33468 11636 33474 11688
rect 28534 11568 28540 11620
rect 28592 11608 28598 11620
rect 28813 11611 28871 11617
rect 28813 11608 28825 11611
rect 28592 11580 28825 11608
rect 28592 11568 28598 11580
rect 28813 11577 28825 11580
rect 28859 11577 28871 11611
rect 28813 11571 28871 11577
rect 28718 11540 28724 11552
rect 27448 11512 28724 11540
rect 28718 11500 28724 11512
rect 28776 11500 28782 11552
rect 31570 11540 31576 11552
rect 31531 11512 31576 11540
rect 31570 11500 31576 11512
rect 31628 11500 31634 11552
rect 32306 11540 32312 11552
rect 32267 11512 32312 11540
rect 32306 11500 32312 11512
rect 32364 11500 32370 11552
rect 1104 11450 34868 11472
rect 1104 11398 5170 11450
rect 5222 11398 5234 11450
rect 5286 11398 5298 11450
rect 5350 11398 5362 11450
rect 5414 11398 5426 11450
rect 5478 11398 13611 11450
rect 13663 11398 13675 11450
rect 13727 11398 13739 11450
rect 13791 11398 13803 11450
rect 13855 11398 13867 11450
rect 13919 11398 22052 11450
rect 22104 11398 22116 11450
rect 22168 11398 22180 11450
rect 22232 11398 22244 11450
rect 22296 11398 22308 11450
rect 22360 11398 30493 11450
rect 30545 11398 30557 11450
rect 30609 11398 30621 11450
rect 30673 11398 30685 11450
rect 30737 11398 30749 11450
rect 30801 11398 34868 11450
rect 1104 11376 34868 11398
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 4522 11336 4528 11348
rect 4203 11308 4528 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 12250 11336 12256 11348
rect 11296 11308 12256 11336
rect 11296 11296 11302 11308
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 20530 11336 20536 11348
rect 20491 11308 20536 11336
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20956 11308 21005 11336
rect 20956 11296 20962 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 27982 11336 27988 11348
rect 20993 11299 21051 11305
rect 22066 11308 27988 11336
rect 13633 11271 13691 11277
rect 13633 11237 13645 11271
rect 13679 11268 13691 11271
rect 15838 11268 15844 11280
rect 13679 11240 15844 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 19518 11268 19524 11280
rect 18248 11240 19524 11268
rect 12164 11212 12216 11218
rect 18248 11209 18276 11240
rect 19518 11228 19524 11240
rect 19576 11268 19582 11280
rect 21082 11268 21088 11280
rect 19576 11240 21088 11268
rect 19576 11228 19582 11240
rect 21082 11228 21088 11240
rect 21140 11228 21146 11280
rect 18233 11203 18291 11209
rect 12164 11154 12216 11160
rect 16776 11172 18000 11200
rect 16776 11144 16804 11172
rect 4522 11092 4528 11144
rect 4580 11132 4586 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 4580 11104 5549 11132
rect 4580 11092 4586 11104
rect 5537 11101 5549 11104
rect 5583 11132 5595 11135
rect 7190 11132 7196 11144
rect 5583 11104 7196 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 7190 11092 7196 11104
rect 7248 11132 7254 11144
rect 10318 11132 10324 11144
rect 7248 11104 10324 11132
rect 7248 11092 7254 11104
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 10588 11135 10646 11141
rect 10588 11101 10600 11135
rect 10634 11132 10646 11135
rect 11054 11132 11060 11144
rect 10634 11104 11060 11132
rect 10634 11101 10646 11104
rect 10588 11095 10646 11101
rect 11054 11092 11060 11104
rect 11112 11132 11118 11144
rect 11974 11132 11980 11144
rect 11112 11104 11980 11132
rect 11112 11092 11118 11104
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12584 11104 12725 11132
rect 12584 11092 12590 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 12894 11132 12900 11144
rect 12759 11104 12900 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 16758 11132 16764 11144
rect 16719 11104 16764 11132
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16942 11132 16948 11144
rect 16903 11104 16948 11132
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17494 11132 17500 11144
rect 17455 11104 17500 11132
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 17972 11141 18000 11172
rect 18233 11169 18245 11203
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 18414 11160 18420 11212
rect 18472 11200 18478 11212
rect 22066 11200 22094 11308
rect 27982 11296 27988 11308
rect 28040 11336 28046 11348
rect 28350 11336 28356 11348
rect 28040 11308 28356 11336
rect 28040 11296 28046 11308
rect 28350 11296 28356 11308
rect 28408 11296 28414 11348
rect 31202 11296 31208 11348
rect 31260 11336 31266 11348
rect 31481 11339 31539 11345
rect 31481 11336 31493 11339
rect 31260 11308 31493 11336
rect 31260 11296 31266 11308
rect 31481 11305 31493 11308
rect 31527 11305 31539 11339
rect 31481 11299 31539 11305
rect 25038 11268 25044 11280
rect 18472 11172 22094 11200
rect 23768 11240 25044 11268
rect 18472 11160 18478 11172
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11101 18015 11135
rect 19886 11132 19892 11144
rect 19847 11104 19892 11132
rect 17957 11095 18015 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20070 11141 20076 11144
rect 20037 11135 20076 11141
rect 20037 11101 20049 11135
rect 20037 11095 20076 11101
rect 20070 11092 20076 11095
rect 20128 11092 20134 11144
rect 20162 11092 20168 11144
rect 20220 11132 20226 11144
rect 20364 11141 20392 11172
rect 20354 11135 20412 11141
rect 20220 11104 20265 11132
rect 20220 11092 20226 11104
rect 20354 11101 20366 11135
rect 20400 11101 20412 11135
rect 21174 11132 21180 11144
rect 21135 11104 21180 11132
rect 20354 11095 20412 11101
rect 21174 11092 21180 11104
rect 21232 11092 21238 11144
rect 21358 11132 21364 11144
rect 21319 11104 21364 11132
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 23768 11141 23796 11240
rect 25038 11228 25044 11240
rect 25096 11268 25102 11280
rect 25774 11268 25780 11280
rect 25096 11240 25780 11268
rect 25096 11228 25102 11240
rect 25774 11228 25780 11240
rect 25832 11228 25838 11280
rect 26142 11200 26148 11212
rect 23952 11172 26148 11200
rect 23952 11141 23980 11172
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 30926 11200 30932 11212
rect 29932 11172 30932 11200
rect 21453 11135 21511 11141
rect 21453 11101 21465 11135
rect 21499 11101 21511 11135
rect 23753 11135 23811 11141
rect 23753 11132 23765 11135
rect 21453 11095 21511 11101
rect 23492 11104 23765 11132
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 3973 11067 4031 11073
rect 3973 11064 3985 11067
rect 3844 11036 3985 11064
rect 3844 11024 3850 11036
rect 3973 11033 3985 11036
rect 4019 11033 4031 11067
rect 3973 11027 4031 11033
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 5804 11067 5862 11073
rect 5804 11064 5816 11067
rect 5684 11036 5816 11064
rect 5684 11024 5690 11036
rect 5804 11033 5816 11036
rect 5850 11064 5862 11067
rect 9306 11064 9312 11076
rect 5850 11036 9312 11064
rect 5850 11033 5862 11036
rect 5804 11027 5862 11033
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 12434 11064 12440 11076
rect 11716 11036 12440 11064
rect 4154 10956 4160 11008
rect 4212 11005 4218 11008
rect 4212 10999 4231 11005
rect 4219 10965 4231 10999
rect 4338 10996 4344 11008
rect 4299 10968 4344 10996
rect 4212 10959 4231 10965
rect 4212 10956 4218 10959
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 6914 10996 6920 11008
rect 6875 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 7374 10956 7380 11008
rect 7432 10996 7438 11008
rect 9766 10996 9772 11008
rect 7432 10968 9772 10996
rect 7432 10956 7438 10968
rect 9766 10956 9772 10968
rect 9824 10996 9830 11008
rect 11238 10996 11244 11008
rect 9824 10968 11244 10996
rect 9824 10956 9830 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 11716 11005 11744 11036
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 12618 11064 12624 11076
rect 12579 11036 12624 11064
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 13446 11064 13452 11076
rect 13407 11036 13452 11064
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 16666 11064 16672 11076
rect 16627 11036 16672 11064
rect 16666 11024 16672 11036
rect 16724 11024 16730 11076
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 20530 11064 20536 11076
rect 20303 11036 20536 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 20898 11024 20904 11076
rect 20956 11064 20962 11076
rect 21468 11064 21496 11095
rect 23492 11064 23520 11104
rect 23753 11101 23765 11104
rect 23799 11101 23811 11135
rect 23753 11095 23811 11101
rect 23937 11135 23995 11141
rect 23937 11101 23949 11135
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 24029 11135 24087 11141
rect 24029 11101 24041 11135
rect 24075 11132 24087 11135
rect 24578 11132 24584 11144
rect 24075 11104 24584 11132
rect 24075 11101 24087 11104
rect 24029 11095 24087 11101
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 26050 11132 26056 11144
rect 26011 11104 26056 11132
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 29362 11092 29368 11144
rect 29420 11132 29426 11144
rect 29932 11141 29960 11172
rect 30926 11160 30932 11172
rect 30984 11160 30990 11212
rect 29917 11135 29975 11141
rect 29917 11132 29929 11135
rect 29420 11104 29929 11132
rect 29420 11092 29426 11104
rect 29917 11101 29929 11104
rect 29963 11101 29975 11135
rect 30190 11132 30196 11144
rect 30151 11104 30196 11132
rect 29917 11095 29975 11101
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 32214 11092 32220 11144
rect 32272 11132 32278 11144
rect 32861 11135 32919 11141
rect 32861 11132 32873 11135
rect 32272 11104 32873 11132
rect 32272 11092 32278 11104
rect 32861 11101 32873 11104
rect 32907 11101 32919 11135
rect 32861 11095 32919 11101
rect 20956 11036 21496 11064
rect 22066 11036 23520 11064
rect 23569 11067 23627 11073
rect 20956 11024 20962 11036
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 12345 10999 12403 11005
rect 12345 10965 12357 10999
rect 12391 10996 12403 10999
rect 12710 10996 12716 11008
rect 12391 10968 12716 10996
rect 12391 10965 12403 10968
rect 12345 10959 12403 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 20438 10956 20444 11008
rect 20496 10996 20502 11008
rect 22066 10996 22094 11036
rect 23569 11033 23581 11067
rect 23615 11064 23627 11067
rect 24854 11064 24860 11076
rect 23615 11036 24860 11064
rect 23615 11033 23627 11036
rect 23569 11027 23627 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 27706 11024 27712 11076
rect 27764 11064 27770 11076
rect 30101 11067 30159 11073
rect 30101 11064 30113 11067
rect 27764 11036 30113 11064
rect 27764 11024 27770 11036
rect 30101 11033 30113 11036
rect 30147 11033 30159 11067
rect 30101 11027 30159 11033
rect 31570 11024 31576 11076
rect 31628 11064 31634 11076
rect 32594 11067 32652 11073
rect 32594 11064 32606 11067
rect 31628 11036 32606 11064
rect 31628 11024 31634 11036
rect 32594 11033 32606 11036
rect 32640 11033 32652 11067
rect 32594 11027 32652 11033
rect 27338 10996 27344 11008
rect 20496 10968 22094 10996
rect 27299 10968 27344 10996
rect 20496 10956 20502 10968
rect 27338 10956 27344 10968
rect 27396 10956 27402 11008
rect 29730 10996 29736 11008
rect 29691 10968 29736 10996
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 1104 10906 35027 10928
rect 1104 10854 9390 10906
rect 9442 10854 9454 10906
rect 9506 10854 9518 10906
rect 9570 10854 9582 10906
rect 9634 10854 9646 10906
rect 9698 10854 17831 10906
rect 17883 10854 17895 10906
rect 17947 10854 17959 10906
rect 18011 10854 18023 10906
rect 18075 10854 18087 10906
rect 18139 10854 26272 10906
rect 26324 10854 26336 10906
rect 26388 10854 26400 10906
rect 26452 10854 26464 10906
rect 26516 10854 26528 10906
rect 26580 10854 34713 10906
rect 34765 10854 34777 10906
rect 34829 10854 34841 10906
rect 34893 10854 34905 10906
rect 34957 10854 34969 10906
rect 35021 10854 35027 10906
rect 1104 10832 35027 10854
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8110 10792 8116 10804
rect 7975 10764 8116 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 9766 10792 9772 10804
rect 8720 10764 8984 10792
rect 8720 10752 8726 10764
rect 2958 10684 2964 10736
rect 3016 10724 3022 10736
rect 3016 10696 3464 10724
rect 3016 10684 3022 10696
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 3436 10665 3464 10696
rect 6730 10684 6736 10736
rect 6788 10724 6794 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 6788 10696 6837 10724
rect 6788 10684 6794 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7101 10727 7159 10733
rect 7101 10724 7113 10727
rect 6972 10696 7113 10724
rect 6972 10684 6978 10696
rect 7101 10693 7113 10696
rect 7147 10693 7159 10727
rect 7101 10687 7159 10693
rect 7193 10727 7251 10733
rect 7193 10693 7205 10727
rect 7239 10724 7251 10727
rect 7374 10724 7380 10736
rect 7239 10696 7380 10724
rect 7239 10693 7251 10696
rect 7193 10687 7251 10693
rect 7374 10684 7380 10696
rect 7432 10684 7438 10736
rect 7558 10724 7564 10736
rect 7519 10696 7564 10724
rect 7558 10684 7564 10696
rect 7616 10684 7622 10736
rect 8570 10684 8576 10736
rect 8628 10724 8634 10736
rect 8849 10727 8907 10733
rect 8849 10724 8861 10727
rect 8628 10696 8861 10724
rect 8628 10684 8634 10696
rect 8849 10693 8861 10696
rect 8895 10693 8907 10727
rect 8956 10724 8984 10764
rect 9232 10764 9772 10792
rect 9232 10733 9260 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 9950 10792 9956 10804
rect 9911 10764 9956 10792
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 10100 10764 13645 10792
rect 10100 10752 10106 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 25498 10752 25504 10804
rect 25556 10792 25562 10804
rect 25593 10795 25651 10801
rect 25593 10792 25605 10795
rect 25556 10764 25605 10792
rect 25556 10752 25562 10764
rect 25593 10761 25605 10764
rect 25639 10761 25651 10795
rect 28166 10792 28172 10804
rect 28127 10764 28172 10792
rect 25593 10755 25651 10761
rect 28166 10752 28172 10764
rect 28224 10752 28230 10804
rect 28718 10752 28724 10804
rect 28776 10792 28782 10804
rect 29917 10795 29975 10801
rect 29917 10792 29929 10795
rect 28776 10764 29929 10792
rect 28776 10752 28782 10764
rect 29917 10761 29929 10764
rect 29963 10761 29975 10795
rect 29917 10755 29975 10761
rect 33594 10752 33600 10804
rect 33652 10792 33658 10804
rect 33689 10795 33747 10801
rect 33689 10792 33701 10795
rect 33652 10764 33701 10792
rect 33652 10752 33658 10764
rect 33689 10761 33701 10764
rect 33735 10761 33747 10795
rect 33689 10755 33747 10761
rect 9084 10727 9142 10733
rect 9084 10724 9096 10727
rect 8956 10696 9096 10724
rect 8849 10687 8907 10693
rect 9084 10693 9096 10696
rect 9130 10693 9142 10727
rect 9084 10687 9142 10693
rect 9217 10727 9275 10733
rect 9217 10693 9229 10727
rect 9263 10693 9275 10727
rect 9217 10687 9275 10693
rect 9398 10684 9404 10736
rect 9456 10724 9462 10736
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 9456 10696 9597 10724
rect 9456 10684 9462 10696
rect 9585 10693 9597 10696
rect 9631 10693 9643 10727
rect 12526 10724 12532 10736
rect 12487 10696 12532 10724
rect 9585 10687 9643 10693
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 12894 10724 12900 10736
rect 12855 10696 12900 10724
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 13262 10724 13268 10736
rect 13223 10696 13268 10724
rect 13262 10684 13268 10696
rect 13320 10684 13326 10736
rect 18230 10724 18236 10736
rect 18191 10696 18236 10724
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 19978 10724 19984 10736
rect 19939 10696 19984 10724
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 25133 10727 25191 10733
rect 25133 10693 25145 10727
rect 25179 10724 25191 10727
rect 27338 10724 27344 10736
rect 25179 10696 27344 10724
rect 25179 10693 25191 10696
rect 25133 10687 25191 10693
rect 27338 10684 27344 10696
rect 27396 10724 27402 10736
rect 28629 10727 28687 10733
rect 28629 10724 28641 10727
rect 27396 10696 28641 10724
rect 27396 10684 27402 10696
rect 28629 10693 28641 10696
rect 28675 10693 28687 10727
rect 30834 10724 30840 10736
rect 30795 10696 30840 10724
rect 28629 10687 28687 10693
rect 30834 10684 30840 10696
rect 30892 10684 30898 10736
rect 31021 10727 31079 10733
rect 31021 10693 31033 10727
rect 31067 10693 31079 10727
rect 31021 10687 31079 10693
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 3108 10628 3249 10656
rect 3108 10616 3114 10628
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10625 3479 10659
rect 3421 10619 3479 10625
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3936 10628 3985 10656
rect 3936 10616 3942 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4246 10656 4252 10668
rect 4203 10628 4252 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 12158 10656 12164 10668
rect 6840 10654 9168 10656
rect 9232 10654 12164 10656
rect 6840 10628 12164 10654
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10557 3203 10591
rect 3326 10588 3332 10600
rect 3287 10560 3332 10588
rect 3145 10551 3203 10557
rect 3160 10520 3188 10551
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6604 10574 6670 10588
rect 6604 10560 6684 10574
rect 6604 10548 6610 10560
rect 3510 10520 3516 10532
rect 3160 10492 3516 10520
rect 3510 10480 3516 10492
rect 3568 10520 3574 10532
rect 4065 10523 4123 10529
rect 4065 10520 4077 10523
rect 3568 10492 4077 10520
rect 3568 10480 3574 10492
rect 4065 10489 4077 10492
rect 4111 10489 4123 10523
rect 6656 10520 6684 10560
rect 6840 10520 6868 10628
rect 8680 10574 8708 10628
rect 9140 10626 9260 10628
rect 12158 10616 12164 10628
rect 12216 10656 12222 10668
rect 12216 10628 12388 10656
rect 12216 10616 12222 10628
rect 12360 10574 12388 10628
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12492 10628 12817 10656
rect 12492 10616 12498 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 25682 10616 25688 10668
rect 25740 10665 25746 10668
rect 25740 10659 25789 10665
rect 25740 10625 25743 10659
rect 25777 10625 25789 10659
rect 25866 10656 25872 10668
rect 25827 10628 25872 10656
rect 25740 10619 25789 10625
rect 25740 10616 25746 10619
rect 25866 10616 25872 10628
rect 25924 10616 25930 10668
rect 25958 10616 25964 10668
rect 26016 10656 26022 10668
rect 26142 10656 26148 10668
rect 26016 10628 26061 10656
rect 26103 10628 26148 10656
rect 26016 10616 26022 10628
rect 26142 10616 26148 10628
rect 26200 10616 26206 10668
rect 26234 10616 26240 10668
rect 26292 10656 26298 10668
rect 27706 10665 27712 10668
rect 27525 10659 27583 10665
rect 26292 10628 26337 10656
rect 26292 10616 26298 10628
rect 27525 10625 27537 10659
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 27673 10659 27712 10665
rect 27673 10625 27685 10659
rect 27673 10619 27712 10625
rect 6656 10492 6868 10520
rect 27540 10520 27568 10619
rect 27706 10616 27712 10619
rect 27764 10616 27770 10668
rect 27801 10659 27859 10665
rect 27801 10625 27813 10659
rect 27847 10625 27859 10659
rect 27801 10619 27859 10625
rect 27816 10588 27844 10619
rect 27890 10616 27896 10668
rect 27948 10656 27954 10668
rect 28031 10659 28089 10665
rect 27948 10628 27993 10656
rect 27948 10616 27954 10628
rect 28031 10625 28043 10659
rect 28077 10656 28089 10659
rect 28350 10656 28356 10668
rect 28077 10628 28356 10656
rect 28077 10625 28089 10628
rect 28031 10619 28089 10625
rect 28350 10616 28356 10628
rect 28408 10656 28414 10668
rect 28902 10656 28908 10668
rect 28408 10628 28908 10656
rect 28408 10616 28414 10628
rect 28902 10616 28908 10628
rect 28960 10616 28966 10668
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 31036 10656 31064 10687
rect 32306 10684 32312 10736
rect 32364 10724 32370 10736
rect 32554 10727 32612 10733
rect 32554 10724 32566 10727
rect 32364 10696 32566 10724
rect 32364 10684 32370 10696
rect 32554 10693 32566 10696
rect 32600 10693 32612 10727
rect 32554 10687 32612 10693
rect 29972 10628 31064 10656
rect 29972 10616 29978 10628
rect 28442 10588 28448 10600
rect 27816 10560 28448 10588
rect 27706 10520 27712 10532
rect 27540 10492 27712 10520
rect 4065 10483 4123 10489
rect 27706 10480 27712 10492
rect 27764 10480 27770 10532
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2961 10455 3019 10461
rect 2961 10452 2973 10455
rect 2832 10424 2973 10452
rect 2832 10412 2838 10424
rect 2961 10421 2973 10424
rect 3007 10421 3019 10455
rect 8110 10452 8116 10464
rect 8071 10424 8116 10452
rect 2961 10415 3019 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 10134 10452 10140 10464
rect 10095 10424 10140 10452
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 13817 10455 13875 10461
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 14366 10452 14372 10464
rect 13863 10424 14372 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 23842 10452 23848 10464
rect 23803 10424 23848 10452
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 25958 10412 25964 10464
rect 26016 10452 26022 10464
rect 27816 10452 27844 10560
rect 28442 10548 28448 10560
rect 28500 10548 28506 10600
rect 32214 10548 32220 10600
rect 32272 10588 32278 10600
rect 32309 10591 32367 10597
rect 32309 10588 32321 10591
rect 32272 10560 32321 10588
rect 32272 10548 32278 10560
rect 32309 10557 32321 10560
rect 32355 10557 32367 10591
rect 32309 10551 32367 10557
rect 31018 10452 31024 10464
rect 26016 10424 27844 10452
rect 30979 10424 31024 10452
rect 26016 10412 26022 10424
rect 31018 10412 31024 10424
rect 31076 10412 31082 10464
rect 31205 10455 31263 10461
rect 31205 10421 31217 10455
rect 31251 10452 31263 10455
rect 32306 10452 32312 10464
rect 31251 10424 32312 10452
rect 31251 10421 31263 10424
rect 31205 10415 31263 10421
rect 32306 10412 32312 10424
rect 32364 10412 32370 10464
rect 1104 10362 34868 10384
rect 1104 10310 5170 10362
rect 5222 10310 5234 10362
rect 5286 10310 5298 10362
rect 5350 10310 5362 10362
rect 5414 10310 5426 10362
rect 5478 10310 13611 10362
rect 13663 10310 13675 10362
rect 13727 10310 13739 10362
rect 13791 10310 13803 10362
rect 13855 10310 13867 10362
rect 13919 10310 22052 10362
rect 22104 10310 22116 10362
rect 22168 10310 22180 10362
rect 22232 10310 22244 10362
rect 22296 10310 22308 10362
rect 22360 10310 30493 10362
rect 30545 10310 30557 10362
rect 30609 10310 30621 10362
rect 30673 10310 30685 10362
rect 30737 10310 30749 10362
rect 30801 10310 34868 10362
rect 1104 10288 34868 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 4062 10248 4068 10260
rect 3108 10220 4068 10248
rect 3108 10208 3114 10220
rect 4062 10208 4068 10220
rect 4120 10248 4126 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4120 10220 4169 10248
rect 4120 10208 4126 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 6730 10248 6736 10260
rect 6691 10220 6736 10248
rect 4157 10211 4215 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 8110 10248 8116 10260
rect 7616 10220 8116 10248
rect 7616 10208 7622 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8662 10248 8668 10260
rect 8619 10220 8668 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 12618 10248 12624 10260
rect 12579 10220 12624 10248
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 25314 10248 25320 10260
rect 21315 10220 25320 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 25314 10208 25320 10220
rect 25372 10208 25378 10260
rect 25961 10251 26019 10257
rect 25961 10217 25973 10251
rect 26007 10248 26019 10251
rect 26142 10248 26148 10260
rect 26007 10220 26148 10248
rect 26007 10217 26019 10220
rect 25961 10211 26019 10217
rect 26142 10208 26148 10220
rect 26200 10208 26206 10260
rect 26234 10208 26240 10260
rect 26292 10248 26298 10260
rect 29733 10251 29791 10257
rect 29733 10248 29745 10251
rect 26292 10220 29745 10248
rect 26292 10208 26298 10220
rect 29733 10217 29745 10220
rect 29779 10217 29791 10251
rect 29733 10211 29791 10217
rect 31665 10251 31723 10257
rect 31665 10217 31677 10251
rect 31711 10248 31723 10251
rect 32214 10248 32220 10260
rect 31711 10220 32220 10248
rect 31711 10217 31723 10220
rect 31665 10211 31723 10217
rect 32214 10208 32220 10220
rect 32272 10208 32278 10260
rect 4341 10183 4399 10189
rect 4341 10149 4353 10183
rect 4387 10149 4399 10183
rect 4341 10143 4399 10149
rect 3237 10115 3295 10121
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3878 10112 3884 10124
rect 3283 10084 3884 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 4356 10112 4384 10143
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 10042 10180 10048 10192
rect 8996 10152 10048 10180
rect 8996 10140 9002 10152
rect 10042 10140 10048 10152
rect 10100 10140 10106 10192
rect 27341 10183 27399 10189
rect 27341 10149 27353 10183
rect 27387 10180 27399 10183
rect 27614 10180 27620 10192
rect 27387 10152 27620 10180
rect 27387 10149 27399 10152
rect 27341 10143 27399 10149
rect 27614 10140 27620 10152
rect 27672 10140 27678 10192
rect 5353 10115 5411 10121
rect 5353 10112 5365 10115
rect 4356 10084 5365 10112
rect 5353 10081 5365 10084
rect 5399 10081 5411 10115
rect 7190 10112 7196 10124
rect 7151 10084 7196 10112
rect 5353 10075 5411 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2685 10047 2743 10053
rect 2685 10044 2697 10047
rect 2271 10016 2697 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2685 10013 2697 10016
rect 2731 10013 2743 10047
rect 2685 10007 2743 10013
rect 2130 9908 2136 9920
rect 2091 9880 2136 9908
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 2700 9908 2728 10007
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2832 10016 2881 10044
rect 2832 10004 2838 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 2961 10007 3019 10013
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 4264 10044 4292 10072
rect 3375 10016 4292 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 2976 9976 3004 10007
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 5368 10044 5396 10075
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 10318 10072 10324 10124
rect 10376 10112 10382 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10376 10084 11253 10112
rect 10376 10072 10382 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 19242 10072 19248 10124
rect 19300 10112 19306 10124
rect 19300 10084 20944 10112
rect 19300 10072 19306 10084
rect 6822 10044 6828 10056
rect 5368 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7466 10053 7472 10056
rect 7460 10044 7472 10053
rect 7427 10016 7472 10044
rect 7460 10007 7472 10016
rect 7466 10004 7472 10007
rect 7524 10004 7530 10056
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10013 17095 10047
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 17037 10007 17095 10013
rect 3970 9976 3976 9988
rect 2976 9948 3976 9976
rect 3344 9920 3372 9948
rect 3970 9936 3976 9948
rect 4028 9936 4034 9988
rect 4189 9979 4247 9985
rect 4189 9945 4201 9979
rect 4235 9976 4247 9979
rect 4356 9976 4384 10004
rect 5626 9985 5632 9988
rect 5620 9976 5632 9985
rect 4235 9948 4384 9976
rect 5587 9948 5632 9976
rect 4235 9945 4247 9948
rect 4189 9939 4247 9945
rect 5620 9939 5632 9948
rect 5626 9936 5632 9939
rect 5684 9936 5690 9988
rect 11514 9985 11520 9988
rect 11508 9976 11520 9985
rect 11427 9948 11520 9976
rect 11508 9939 11520 9948
rect 11572 9976 11578 9988
rect 11790 9976 11796 9988
rect 11572 9948 11796 9976
rect 11514 9936 11520 9939
rect 11572 9936 11578 9948
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 3053 9911 3111 9917
rect 3053 9908 3065 9911
rect 2700 9880 3065 9908
rect 3053 9877 3065 9880
rect 3099 9877 3111 9911
rect 3053 9871 3111 9877
rect 3326 9868 3332 9920
rect 3384 9868 3390 9920
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 13354 9908 13360 9920
rect 8168 9880 13360 9908
rect 8168 9868 8174 9880
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 16632 9880 16865 9908
rect 16632 9868 16638 9880
rect 16853 9877 16865 9880
rect 16899 9877 16911 9911
rect 17052 9908 17080 10007
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 20622 10044 20628 10056
rect 20583 10016 20628 10044
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 20916 10053 20944 10084
rect 23842 10072 23848 10124
rect 23900 10112 23906 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 23900 10084 24593 10112
rect 23900 10072 23906 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 28718 10112 28724 10124
rect 28679 10084 28724 10112
rect 24581 10075 24639 10081
rect 28718 10072 28724 10084
rect 28776 10072 28782 10124
rect 28902 10072 28908 10124
rect 28960 10112 28966 10124
rect 28960 10084 30144 10112
rect 28960 10072 28966 10084
rect 20718 10047 20776 10053
rect 20718 10013 20730 10047
rect 20764 10013 20776 10047
rect 20718 10007 20776 10013
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 17218 9976 17224 9988
rect 17131 9948 17224 9976
rect 17218 9936 17224 9948
rect 17276 9976 17282 9988
rect 20732 9976 20760 10007
rect 21082 10004 21088 10056
rect 21140 10053 21146 10056
rect 24854 10053 24860 10056
rect 21140 10044 21148 10053
rect 24848 10044 24860 10053
rect 21140 10016 21185 10044
rect 24815 10016 24860 10044
rect 21140 10007 21148 10016
rect 24848 10007 24860 10016
rect 21140 10004 21146 10007
rect 24854 10004 24860 10007
rect 24912 10004 24918 10056
rect 28465 10047 28523 10053
rect 28465 10013 28477 10047
rect 28511 10044 28523 10047
rect 29730 10044 29736 10056
rect 28511 10016 29736 10044
rect 28511 10013 28523 10016
rect 28465 10007 28523 10013
rect 29730 10004 29736 10016
rect 29788 10004 29794 10056
rect 29914 10004 29920 10056
rect 29972 10044 29978 10056
rect 30116 10053 30144 10084
rect 30101 10047 30159 10053
rect 29972 10016 30065 10044
rect 29972 10004 29978 10016
rect 30101 10013 30113 10047
rect 30147 10013 30159 10047
rect 30282 10044 30288 10056
rect 30243 10016 30288 10044
rect 30101 10007 30159 10013
rect 30282 10004 30288 10016
rect 30340 10004 30346 10056
rect 33410 10044 33416 10056
rect 33371 10016 33416 10044
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33686 10044 33692 10056
rect 33647 10016 33692 10044
rect 33686 10004 33692 10016
rect 33744 10004 33750 10056
rect 17276 9948 20760 9976
rect 20993 9979 21051 9985
rect 17276 9936 17282 9948
rect 20993 9945 21005 9979
rect 21039 9945 21051 9979
rect 20993 9939 21051 9945
rect 20438 9908 20444 9920
rect 17052 9880 20444 9908
rect 16853 9871 16911 9877
rect 20438 9868 20444 9880
rect 20496 9908 20502 9920
rect 20622 9908 20628 9920
rect 20496 9880 20628 9908
rect 20496 9868 20502 9880
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 20806 9868 20812 9920
rect 20864 9908 20870 9920
rect 21008 9908 21036 9939
rect 28994 9936 29000 9988
rect 29052 9976 29058 9988
rect 29932 9976 29960 10004
rect 29052 9948 29960 9976
rect 30009 9979 30067 9985
rect 29052 9936 29058 9948
rect 30009 9945 30021 9979
rect 30055 9945 30067 9979
rect 30009 9939 30067 9945
rect 32953 9979 33011 9985
rect 32953 9945 32965 9979
rect 32999 9976 33011 9979
rect 32999 9948 33732 9976
rect 32999 9945 33011 9948
rect 32953 9939 33011 9945
rect 20864 9880 21036 9908
rect 30024 9908 30052 9939
rect 33704 9920 33732 9948
rect 32214 9908 32220 9920
rect 30024 9880 32220 9908
rect 20864 9868 20870 9880
rect 32214 9868 32220 9880
rect 32272 9908 32278 9920
rect 33505 9911 33563 9917
rect 33505 9908 33517 9911
rect 32272 9880 33517 9908
rect 32272 9868 32278 9880
rect 33505 9877 33517 9880
rect 33551 9877 33563 9911
rect 33505 9871 33563 9877
rect 33686 9868 33692 9920
rect 33744 9868 33750 9920
rect 33870 9908 33876 9920
rect 33831 9880 33876 9908
rect 33870 9868 33876 9880
rect 33928 9868 33934 9920
rect 1104 9818 35027 9840
rect 1104 9766 9390 9818
rect 9442 9766 9454 9818
rect 9506 9766 9518 9818
rect 9570 9766 9582 9818
rect 9634 9766 9646 9818
rect 9698 9766 17831 9818
rect 17883 9766 17895 9818
rect 17947 9766 17959 9818
rect 18011 9766 18023 9818
rect 18075 9766 18087 9818
rect 18139 9766 26272 9818
rect 26324 9766 26336 9818
rect 26388 9766 26400 9818
rect 26452 9766 26464 9818
rect 26516 9766 26528 9818
rect 26580 9766 34713 9818
rect 34765 9766 34777 9818
rect 34829 9766 34841 9818
rect 34893 9766 34905 9818
rect 34957 9766 34969 9818
rect 35021 9766 35027 9818
rect 1104 9744 35027 9766
rect 4249 9707 4307 9713
rect 4249 9673 4261 9707
rect 4295 9704 4307 9707
rect 4338 9704 4344 9716
rect 4295 9676 4344 9704
rect 4295 9673 4307 9676
rect 4249 9667 4307 9673
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 8570 9704 8576 9716
rect 8531 9676 8576 9704
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 10134 9664 10140 9716
rect 10192 9704 10198 9716
rect 17126 9704 17132 9716
rect 10192 9676 17132 9704
rect 10192 9664 10198 9676
rect 17126 9664 17132 9676
rect 17184 9664 17190 9716
rect 27706 9704 27712 9716
rect 27667 9676 27712 9704
rect 27706 9664 27712 9676
rect 27764 9664 27770 9716
rect 2317 9639 2375 9645
rect 2317 9605 2329 9639
rect 2363 9636 2375 9639
rect 2498 9636 2504 9648
rect 2363 9608 2504 9636
rect 2363 9605 2375 9608
rect 2317 9599 2375 9605
rect 2498 9596 2504 9608
rect 2556 9636 2562 9648
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2556 9608 3341 9636
rect 2556 9596 2562 9608
rect 3329 9605 3341 9608
rect 3375 9605 3387 9639
rect 3329 9599 3387 9605
rect 3602 9596 3608 9648
rect 3660 9636 3666 9648
rect 3970 9636 3976 9648
rect 3660 9608 3976 9636
rect 3660 9596 3666 9608
rect 3970 9596 3976 9608
rect 4028 9636 4034 9648
rect 7466 9645 7472 9648
rect 4065 9639 4123 9645
rect 4065 9636 4077 9639
rect 4028 9608 4077 9636
rect 4028 9596 4034 9608
rect 4065 9605 4077 9608
rect 4111 9605 4123 9639
rect 7460 9636 7472 9645
rect 7427 9608 7472 9636
rect 4065 9599 4123 9605
rect 7460 9599 7472 9608
rect 7466 9596 7472 9599
rect 7524 9596 7530 9648
rect 17494 9596 17500 9648
rect 17552 9636 17558 9648
rect 17552 9608 19472 9636
rect 17552 9596 17558 9608
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 3142 9568 3148 9580
rect 2455 9540 3148 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2148 9500 2176 9531
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 4522 9568 4528 9580
rect 4483 9540 4528 9568
rect 3237 9531 3295 9537
rect 3050 9500 3056 9512
rect 2148 9472 3056 9500
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9364 2007 9367
rect 2590 9364 2596 9376
rect 1995 9336 2596 9364
rect 1995 9333 2007 9336
rect 1949 9327 2007 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 2866 9364 2872 9376
rect 2827 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 3252 9364 3280 9531
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 3510 9500 3516 9512
rect 3471 9472 3516 9500
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 5000 9500 5028 9531
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 6880 9540 7205 9568
rect 6880 9528 6886 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 11957 9571 12015 9577
rect 11957 9568 11969 9571
rect 11848 9540 11969 9568
rect 11848 9528 11854 9540
rect 11957 9537 11969 9540
rect 12003 9537 12015 9571
rect 11957 9531 12015 9537
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 17589 9571 17647 9577
rect 17589 9568 17601 9571
rect 17460 9540 17601 9568
rect 17460 9528 17466 9540
rect 17589 9537 17601 9540
rect 17635 9537 17647 9571
rect 17770 9568 17776 9580
rect 17731 9540 17776 9568
rect 17589 9531 17647 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18325 9571 18383 9577
rect 17920 9540 17965 9568
rect 17920 9528 17926 9540
rect 18325 9537 18337 9571
rect 18371 9537 18383 9571
rect 18506 9568 18512 9580
rect 18467 9540 18512 9568
rect 18325 9531 18383 9537
rect 4120 9472 5028 9500
rect 4120 9460 4126 9472
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 10836 9472 11713 9500
rect 10836 9460 10842 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 17678 9460 17684 9512
rect 17736 9500 17742 9512
rect 18340 9500 18368 9531
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 18782 9568 18788 9580
rect 18739 9540 18788 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 17736 9472 18368 9500
rect 17736 9460 17742 9472
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4264 9404 5089 9432
rect 4264 9373 4292 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 5077 9395 5135 9401
rect 12710 9392 12716 9444
rect 12768 9432 12774 9444
rect 13081 9435 13139 9441
rect 13081 9432 13093 9435
rect 12768 9404 13093 9432
rect 12768 9392 12774 9404
rect 13081 9401 13093 9404
rect 13127 9401 13139 9435
rect 13081 9395 13139 9401
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 18616 9432 18644 9531
rect 18782 9528 18788 9540
rect 18840 9568 18846 9580
rect 19334 9568 19340 9580
rect 18840 9540 19340 9568
rect 18840 9528 18846 9540
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19444 9577 19472 9608
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 19576 9608 19840 9636
rect 19576 9596 19582 9608
rect 19812 9577 19840 9608
rect 20346 9596 20352 9648
rect 20404 9636 20410 9648
rect 20990 9636 20996 9648
rect 20404 9608 20996 9636
rect 20404 9596 20410 9608
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 25682 9596 25688 9648
rect 25740 9636 25746 9648
rect 27341 9639 27399 9645
rect 27341 9636 27353 9639
rect 25740 9608 27353 9636
rect 25740 9596 25746 9608
rect 27341 9605 27353 9608
rect 27387 9605 27399 9639
rect 27341 9599 27399 9605
rect 27433 9639 27491 9645
rect 27433 9605 27445 9639
rect 27479 9636 27491 9639
rect 31386 9636 31392 9648
rect 27479 9608 31392 9636
rect 27479 9605 27491 9608
rect 27433 9599 27491 9605
rect 31386 9596 31392 9608
rect 31444 9596 31450 9648
rect 32306 9636 32312 9648
rect 32267 9608 32312 9636
rect 32306 9596 32312 9608
rect 32364 9596 32370 9648
rect 19429 9571 19487 9577
rect 19429 9537 19441 9571
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 19797 9531 19855 9537
rect 19242 9500 19248 9512
rect 18380 9404 18644 9432
rect 18800 9472 19248 9500
rect 18380 9392 18386 9404
rect 4249 9367 4307 9373
rect 4249 9364 4261 9367
rect 3252 9336 4261 9364
rect 4249 9333 4261 9336
rect 4295 9333 4307 9367
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 4249 9327 4307 9333
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 18800 9364 18828 9472
rect 19242 9460 19248 9472
rect 19300 9500 19306 9512
rect 19628 9500 19656 9531
rect 19300 9472 19656 9500
rect 19720 9500 19748 9531
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 20806 9568 20812 9580
rect 20767 9540 20812 9568
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 20956 9540 21001 9568
rect 20956 9528 20962 9540
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26016 9540 27169 9568
rect 26016 9528 26022 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9568 27583 9571
rect 27798 9568 27804 9580
rect 27571 9540 27804 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 27798 9528 27804 9540
rect 27856 9568 27862 9580
rect 28902 9568 28908 9580
rect 27856 9540 28908 9568
rect 27856 9528 27862 9540
rect 28902 9528 28908 9540
rect 28960 9528 28966 9580
rect 30190 9528 30196 9580
rect 30248 9568 30254 9580
rect 31297 9571 31355 9577
rect 31297 9568 31309 9571
rect 30248 9540 31309 9568
rect 30248 9528 30254 9540
rect 31297 9537 31309 9540
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 31573 9571 31631 9577
rect 31573 9537 31585 9571
rect 31619 9537 31631 9571
rect 31573 9531 31631 9537
rect 23658 9500 23664 9512
rect 19720 9472 23664 9500
rect 19300 9460 19306 9472
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 29362 9460 29368 9512
rect 29420 9500 29426 9512
rect 31588 9500 31616 9531
rect 29420 9472 31616 9500
rect 29420 9460 29426 9472
rect 18877 9435 18935 9441
rect 18877 9401 18889 9435
rect 18923 9432 18935 9435
rect 19794 9432 19800 9444
rect 18923 9404 19800 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 19886 9392 19892 9444
rect 19944 9432 19950 9444
rect 19981 9435 20039 9441
rect 19981 9432 19993 9435
rect 19944 9404 19993 9432
rect 19944 9392 19950 9404
rect 19981 9401 19993 9404
rect 20027 9401 20039 9435
rect 21082 9432 21088 9444
rect 19981 9395 20039 9401
rect 20272 9404 21088 9432
rect 18564 9336 18828 9364
rect 18564 9324 18570 9336
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 20272 9364 20300 9404
rect 21082 9392 21088 9404
rect 21140 9392 21146 9444
rect 21174 9392 21180 9444
rect 21232 9432 21238 9444
rect 27246 9432 27252 9444
rect 21232 9404 27252 9432
rect 21232 9392 21238 9404
rect 27246 9392 27252 9404
rect 27304 9392 27310 9444
rect 20438 9364 20444 9376
rect 19392 9336 20300 9364
rect 20399 9336 20444 9364
rect 19392 9324 19398 9336
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 28810 9364 28816 9376
rect 20588 9336 28816 9364
rect 20588 9324 20594 9336
rect 28810 9324 28816 9336
rect 28868 9324 28874 9376
rect 31754 9364 31760 9376
rect 31715 9336 31760 9364
rect 31754 9324 31760 9336
rect 31812 9324 31818 9376
rect 33597 9367 33655 9373
rect 33597 9333 33609 9367
rect 33643 9364 33655 9367
rect 33686 9364 33692 9376
rect 33643 9336 33692 9364
rect 33643 9333 33655 9336
rect 33597 9327 33655 9333
rect 33686 9324 33692 9336
rect 33744 9324 33750 9376
rect 1104 9274 34868 9296
rect 1104 9222 5170 9274
rect 5222 9222 5234 9274
rect 5286 9222 5298 9274
rect 5350 9222 5362 9274
rect 5414 9222 5426 9274
rect 5478 9222 13611 9274
rect 13663 9222 13675 9274
rect 13727 9222 13739 9274
rect 13791 9222 13803 9274
rect 13855 9222 13867 9274
rect 13919 9222 22052 9274
rect 22104 9222 22116 9274
rect 22168 9222 22180 9274
rect 22232 9222 22244 9274
rect 22296 9222 22308 9274
rect 22360 9222 30493 9274
rect 30545 9222 30557 9274
rect 30609 9222 30621 9274
rect 30673 9222 30685 9274
rect 30737 9222 30749 9274
rect 30801 9222 34868 9274
rect 1104 9200 34868 9222
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2682 9160 2688 9172
rect 2188 9132 2688 9160
rect 2188 9120 2194 9132
rect 2682 9120 2688 9132
rect 2740 9160 2746 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2740 9132 2973 9160
rect 2740 9120 2746 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12526 9160 12532 9172
rect 12207 9132 12532 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 16393 9163 16451 9169
rect 16393 9129 16405 9163
rect 16439 9160 16451 9163
rect 17218 9160 17224 9172
rect 16439 9132 17224 9160
rect 16439 9129 16451 9132
rect 16393 9123 16451 9129
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 20806 9120 20812 9172
rect 20864 9160 20870 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 20864 9132 21281 9160
rect 20864 9120 20870 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 27430 9160 27436 9172
rect 22888 9132 27436 9160
rect 22888 9120 22894 9132
rect 27430 9120 27436 9132
rect 27488 9120 27494 9172
rect 32214 9120 32220 9172
rect 32272 9160 32278 9172
rect 32309 9163 32367 9169
rect 32309 9160 32321 9163
rect 32272 9132 32321 9160
rect 32272 9120 32278 9132
rect 32309 9129 32321 9132
rect 32355 9129 32367 9163
rect 32309 9123 32367 9129
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2777 9095 2835 9101
rect 2777 9092 2789 9095
rect 2556 9064 2789 9092
rect 2556 9052 2562 9064
rect 2777 9061 2789 9064
rect 2823 9092 2835 9095
rect 3694 9092 3700 9104
rect 2823 9064 3700 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 3694 9052 3700 9064
rect 3752 9092 3758 9104
rect 30374 9092 30380 9104
rect 3752 9064 4016 9092
rect 3752 9052 3758 9064
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3988 9033 4016 9064
rect 24964 9064 30380 9092
rect 3973 9027 4031 9033
rect 3016 8996 3372 9024
rect 3016 8984 3022 8996
rect 3344 8965 3372 8996
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 10778 9024 10784 9036
rect 6880 8996 10784 9024
rect 6880 8984 6886 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 20990 8984 20996 9036
rect 21048 9024 21054 9036
rect 24964 9024 24992 9064
rect 21048 8996 24992 9024
rect 21048 8984 21054 8996
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4338 8956 4344 8968
rect 4203 8928 4344 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 11054 8965 11060 8968
rect 11048 8956 11060 8965
rect 11015 8928 11060 8956
rect 11048 8919 11060 8928
rect 11054 8916 11060 8919
rect 11112 8916 11118 8968
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8956 15071 8959
rect 15102 8956 15108 8968
rect 15059 8928 15108 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16356 8928 16865 8956
rect 16356 8916 16362 8928
rect 16853 8925 16865 8928
rect 16899 8956 16911 8959
rect 19518 8956 19524 8968
rect 16899 8928 19524 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 19886 8956 19892 8968
rect 19847 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 20156 8959 20214 8965
rect 20156 8925 20168 8959
rect 20202 8956 20214 8959
rect 20438 8956 20444 8968
rect 20202 8928 20444 8956
rect 20202 8925 20214 8928
rect 20156 8919 20214 8925
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 22664 8965 22692 8996
rect 22649 8959 22707 8965
rect 22649 8925 22661 8959
rect 22695 8925 22707 8959
rect 22830 8956 22836 8968
rect 22791 8928 22836 8956
rect 22649 8919 22707 8925
rect 22830 8916 22836 8928
rect 22888 8916 22894 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8925 22983 8959
rect 24578 8956 24584 8968
rect 24539 8928 24584 8956
rect 22925 8919 22983 8925
rect 2866 8848 2872 8900
rect 2924 8897 2930 8900
rect 2924 8891 2973 8897
rect 2924 8857 2927 8891
rect 2961 8857 2973 8891
rect 2924 8851 2973 8857
rect 15280 8891 15338 8897
rect 15280 8857 15292 8891
rect 15326 8888 15338 8891
rect 16574 8888 16580 8900
rect 15326 8860 16580 8888
rect 15326 8857 15338 8860
rect 15280 8851 15338 8857
rect 2924 8848 2930 8851
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 17120 8891 17178 8897
rect 17120 8857 17132 8891
rect 17166 8888 17178 8891
rect 17402 8888 17408 8900
rect 17166 8860 17408 8888
rect 17166 8857 17178 8860
rect 17120 8851 17178 8857
rect 17402 8848 17408 8860
rect 17460 8848 17466 8900
rect 17862 8888 17868 8900
rect 17696 8860 17868 8888
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17696 8820 17724 8860
rect 17862 8848 17868 8860
rect 17920 8888 17926 8900
rect 22940 8888 22968 8919
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 24964 8956 24992 8996
rect 24903 8928 24992 8956
rect 28721 8959 28779 8965
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 28721 8925 28733 8959
rect 28767 8925 28779 8959
rect 28721 8919 28779 8925
rect 17920 8860 22968 8888
rect 17920 8848 17926 8860
rect 23658 8848 23664 8900
rect 23716 8888 23722 8900
rect 24673 8891 24731 8897
rect 24673 8888 24685 8891
rect 23716 8860 24685 8888
rect 23716 8848 23722 8860
rect 24673 8857 24685 8860
rect 24719 8857 24731 8891
rect 28736 8888 28764 8919
rect 28810 8916 28816 8968
rect 28868 8956 28874 8968
rect 29012 8965 29040 9064
rect 30374 9052 30380 9064
rect 30432 9052 30438 9104
rect 28997 8959 29055 8965
rect 28868 8928 28913 8956
rect 28868 8916 28874 8928
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29086 8916 29092 8968
rect 29144 8956 29150 8968
rect 29917 8959 29975 8965
rect 29917 8956 29929 8959
rect 29144 8928 29929 8956
rect 29144 8916 29150 8928
rect 29917 8925 29929 8928
rect 29963 8925 29975 8959
rect 30190 8956 30196 8968
rect 29917 8919 29975 8925
rect 30024 8928 30196 8956
rect 30024 8888 30052 8928
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 32306 8916 32312 8968
rect 32364 8956 32370 8968
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 32364 8928 33701 8956
rect 32364 8916 32370 8928
rect 33689 8925 33701 8928
rect 33735 8925 33747 8959
rect 33689 8919 33747 8925
rect 28736 8860 30052 8888
rect 30101 8891 30159 8897
rect 24673 8851 24731 8857
rect 29012 8832 29040 8860
rect 30101 8857 30113 8891
rect 30147 8888 30159 8891
rect 30282 8888 30288 8900
rect 30147 8860 30288 8888
rect 30147 8857 30159 8860
rect 30101 8851 30159 8857
rect 30282 8848 30288 8860
rect 30340 8848 30346 8900
rect 33444 8891 33502 8897
rect 33444 8857 33456 8891
rect 33490 8888 33502 8891
rect 33870 8888 33876 8900
rect 33490 8860 33876 8888
rect 33490 8857 33502 8860
rect 33444 8851 33502 8857
rect 33870 8848 33876 8860
rect 33928 8848 33934 8900
rect 17276 8792 17724 8820
rect 17276 8780 17282 8792
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 18233 8823 18291 8829
rect 18233 8820 18245 8823
rect 17828 8792 18245 8820
rect 17828 8780 17834 8792
rect 18233 8789 18245 8792
rect 18279 8820 18291 8823
rect 20438 8820 20444 8832
rect 18279 8792 20444 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 21818 8780 21824 8832
rect 21876 8820 21882 8832
rect 22465 8823 22523 8829
rect 22465 8820 22477 8823
rect 21876 8792 22477 8820
rect 21876 8780 21882 8792
rect 22465 8789 22477 8792
rect 22511 8789 22523 8823
rect 25038 8820 25044 8832
rect 24999 8792 25044 8820
rect 22465 8783 22523 8789
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 25774 8780 25780 8832
rect 25832 8820 25838 8832
rect 28902 8820 28908 8832
rect 25832 8792 28908 8820
rect 25832 8780 25838 8792
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 28994 8780 29000 8832
rect 29052 8780 29058 8832
rect 29178 8820 29184 8832
rect 29139 8792 29184 8820
rect 29178 8780 29184 8792
rect 29236 8780 29242 8832
rect 29730 8820 29736 8832
rect 29691 8792 29736 8820
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 1104 8730 35027 8752
rect 1104 8678 9390 8730
rect 9442 8678 9454 8730
rect 9506 8678 9518 8730
rect 9570 8678 9582 8730
rect 9634 8678 9646 8730
rect 9698 8678 17831 8730
rect 17883 8678 17895 8730
rect 17947 8678 17959 8730
rect 18011 8678 18023 8730
rect 18075 8678 18087 8730
rect 18139 8678 26272 8730
rect 26324 8678 26336 8730
rect 26388 8678 26400 8730
rect 26452 8678 26464 8730
rect 26516 8678 26528 8730
rect 26580 8678 34713 8730
rect 34765 8678 34777 8730
rect 34829 8678 34841 8730
rect 34893 8678 34905 8730
rect 34957 8678 34969 8730
rect 35021 8678 35027 8730
rect 1104 8656 35027 8678
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3602 8616 3608 8628
rect 3563 8588 3608 8616
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 14921 8619 14979 8625
rect 14921 8585 14933 8619
rect 14967 8616 14979 8619
rect 17678 8616 17684 8628
rect 14967 8588 17684 8616
rect 14967 8585 14979 8588
rect 14921 8579 14979 8585
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 20898 8616 20904 8628
rect 17788 8588 20904 8616
rect 9585 8551 9643 8557
rect 9585 8517 9597 8551
rect 9631 8548 9643 8551
rect 12066 8548 12072 8560
rect 9631 8520 12072 8548
rect 9631 8517 9643 8520
rect 9585 8511 9643 8517
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 16056 8551 16114 8557
rect 16056 8517 16068 8551
rect 16102 8548 16114 8551
rect 17310 8548 17316 8560
rect 16102 8520 17316 8548
rect 16102 8517 16114 8520
rect 16056 8511 16114 8517
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 2590 8480 2596 8492
rect 2551 8452 2596 8480
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2869 8483 2927 8489
rect 2869 8480 2881 8483
rect 2832 8452 2881 8480
rect 2832 8440 2838 8452
rect 2869 8449 2881 8452
rect 2915 8449 2927 8483
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 2869 8443 2927 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 16298 8480 16304 8492
rect 16259 8452 16304 8480
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 17034 8440 17040 8492
rect 17092 8480 17098 8492
rect 17788 8489 17816 8588
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 22554 8576 22560 8628
rect 22612 8616 22618 8628
rect 23658 8616 23664 8628
rect 22612 8588 22968 8616
rect 23619 8588 23664 8616
rect 22612 8576 22618 8588
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 20625 8551 20683 8557
rect 20625 8548 20637 8551
rect 18564 8520 20637 8548
rect 18564 8508 18570 8520
rect 20625 8517 20637 8520
rect 20671 8517 20683 8551
rect 20625 8511 20683 8517
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 20990 8548 20996 8560
rect 20763 8520 20996 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 20990 8508 20996 8520
rect 21048 8508 21054 8560
rect 22738 8548 22744 8560
rect 22699 8520 22744 8548
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 22940 8557 22968 8588
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 25682 8616 25688 8628
rect 24136 8588 25688 8616
rect 22925 8551 22983 8557
rect 22925 8517 22937 8551
rect 22971 8548 22983 8551
rect 24136 8548 24164 8588
rect 25682 8576 25688 8588
rect 25740 8576 25746 8628
rect 25866 8616 25872 8628
rect 25827 8588 25872 8616
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 30009 8619 30067 8625
rect 28960 8588 29224 8616
rect 28960 8576 28966 8588
rect 22971 8520 24164 8548
rect 24796 8551 24854 8557
rect 22971 8517 22983 8520
rect 22925 8511 22983 8517
rect 24796 8517 24808 8551
rect 24842 8548 24854 8551
rect 25038 8548 25044 8560
rect 24842 8520 25044 8548
rect 24842 8517 24854 8520
rect 24796 8511 24854 8517
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 29086 8548 29092 8560
rect 28644 8520 29092 8548
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 17092 8452 17509 8480
rect 17092 8440 17098 8452
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 18230 8480 18236 8492
rect 18191 8452 18236 8480
rect 17773 8443 17831 8449
rect 17696 8412 17724 8443
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 20438 8480 20444 8492
rect 20399 8452 20444 8480
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20530 8440 20536 8492
rect 20588 8480 20594 8492
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20588 8452 20821 8480
rect 20588 8440 20594 8452
rect 20809 8449 20821 8452
rect 20855 8480 20867 8483
rect 21082 8480 21088 8492
rect 20855 8452 21088 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 24946 8440 24952 8492
rect 25004 8480 25010 8492
rect 25501 8483 25559 8489
rect 25501 8480 25513 8483
rect 25004 8452 25513 8480
rect 25004 8440 25010 8452
rect 25501 8449 25513 8452
rect 25547 8449 25559 8483
rect 25501 8443 25559 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8480 25743 8483
rect 25774 8480 25780 8492
rect 25731 8452 25780 8480
rect 25731 8449 25743 8452
rect 25685 8443 25743 8449
rect 25774 8440 25780 8452
rect 25832 8440 25838 8492
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8480 26019 8483
rect 26050 8480 26056 8492
rect 26007 8452 26056 8480
rect 26007 8449 26019 8452
rect 25961 8443 26019 8449
rect 26050 8440 26056 8452
rect 26108 8440 26114 8492
rect 28644 8489 28672 8520
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 29196 8548 29224 8588
rect 30009 8585 30021 8619
rect 30055 8616 30067 8619
rect 30282 8616 30288 8628
rect 30055 8588 30288 8616
rect 30055 8585 30067 8588
rect 30009 8579 30067 8585
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 31386 8576 31392 8628
rect 31444 8616 31450 8628
rect 33689 8619 33747 8625
rect 33689 8616 33701 8619
rect 31444 8588 33701 8616
rect 31444 8576 31450 8588
rect 33689 8585 33701 8588
rect 33735 8585 33747 8619
rect 33689 8579 33747 8585
rect 30469 8551 30527 8557
rect 30469 8548 30481 8551
rect 29196 8520 30481 8548
rect 30469 8517 30481 8520
rect 30515 8517 30527 8551
rect 30469 8511 30527 8517
rect 30576 8520 30972 8548
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8449 28687 8483
rect 28629 8443 28687 8449
rect 28896 8483 28954 8489
rect 28896 8449 28908 8483
rect 28942 8480 28954 8483
rect 29730 8480 29736 8492
rect 28942 8452 29736 8480
rect 28942 8449 28954 8452
rect 28896 8443 28954 8449
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 30190 8440 30196 8492
rect 30248 8480 30254 8492
rect 30576 8480 30604 8520
rect 30248 8452 30604 8480
rect 30653 8483 30711 8489
rect 30248 8440 30254 8452
rect 30653 8449 30665 8483
rect 30699 8449 30711 8483
rect 30834 8480 30840 8492
rect 30795 8452 30840 8480
rect 30653 8443 30711 8449
rect 18322 8412 18328 8424
rect 17696 8384 18328 8412
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 19886 8372 19892 8424
rect 19944 8412 19950 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19944 8384 19993 8412
rect 19944 8372 19950 8384
rect 19981 8381 19993 8384
rect 20027 8412 20039 8415
rect 21266 8412 21272 8424
rect 20027 8384 21272 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 25038 8412 25044 8424
rect 24999 8384 25044 8412
rect 25038 8372 25044 8384
rect 25096 8372 25102 8424
rect 30668 8412 30696 8443
rect 30834 8440 30840 8452
rect 30892 8440 30898 8492
rect 30944 8489 30972 8520
rect 31754 8508 31760 8560
rect 31812 8548 31818 8560
rect 32554 8551 32612 8557
rect 32554 8548 32566 8551
rect 31812 8520 32566 8548
rect 31812 8508 31818 8520
rect 32554 8517 32566 8520
rect 32600 8517 32612 8551
rect 32554 8511 32612 8517
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8449 30987 8483
rect 32122 8480 32128 8492
rect 30929 8443 30987 8449
rect 31726 8452 32128 8480
rect 31726 8412 31754 8452
rect 32122 8440 32128 8452
rect 32180 8440 32186 8492
rect 32306 8480 32312 8492
rect 32267 8452 32312 8480
rect 32306 8440 32312 8452
rect 32364 8440 32370 8492
rect 30668 8384 31754 8412
rect 17313 8347 17371 8353
rect 17313 8313 17325 8347
rect 17359 8344 17371 8347
rect 19702 8344 19708 8356
rect 17359 8316 19708 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 19702 8304 19708 8316
rect 19760 8304 19766 8356
rect 20993 8347 21051 8353
rect 20993 8313 21005 8347
rect 21039 8344 21051 8347
rect 21174 8344 21180 8356
rect 21039 8316 21180 8344
rect 21039 8313 21051 8316
rect 20993 8307 21051 8313
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 23109 8347 23167 8353
rect 23109 8313 23121 8347
rect 23155 8344 23167 8347
rect 24026 8344 24032 8356
rect 23155 8316 24032 8344
rect 23155 8313 23167 8316
rect 23109 8307 23167 8313
rect 24026 8304 24032 8316
rect 24084 8304 24090 8356
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8276 8171 8279
rect 8202 8276 8208 8288
rect 8159 8248 8208 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 18506 8276 18512 8288
rect 16724 8248 18512 8276
rect 16724 8236 16730 8248
rect 18506 8236 18512 8248
rect 18564 8236 18570 8288
rect 21726 8236 21732 8288
rect 21784 8276 21790 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 21784 8248 22937 8276
rect 21784 8236 21790 8248
rect 22925 8245 22937 8248
rect 22971 8276 22983 8279
rect 28074 8276 28080 8288
rect 22971 8248 28080 8276
rect 22971 8245 22983 8248
rect 22925 8239 22983 8245
rect 28074 8236 28080 8248
rect 28132 8236 28138 8288
rect 1104 8186 34868 8208
rect 1104 8134 5170 8186
rect 5222 8134 5234 8186
rect 5286 8134 5298 8186
rect 5350 8134 5362 8186
rect 5414 8134 5426 8186
rect 5478 8134 13611 8186
rect 13663 8134 13675 8186
rect 13727 8134 13739 8186
rect 13791 8134 13803 8186
rect 13855 8134 13867 8186
rect 13919 8134 22052 8186
rect 22104 8134 22116 8186
rect 22168 8134 22180 8186
rect 22232 8134 22244 8186
rect 22296 8134 22308 8186
rect 22360 8134 30493 8186
rect 30545 8134 30557 8186
rect 30609 8134 30621 8186
rect 30673 8134 30685 8186
rect 30737 8134 30749 8186
rect 30801 8134 34868 8186
rect 1104 8112 34868 8134
rect 18230 8032 18236 8084
rect 18288 8072 18294 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 18288 8044 22937 8072
rect 18288 8032 18294 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 28261 8075 28319 8081
rect 28261 8072 28273 8075
rect 28132 8044 28273 8072
rect 28132 8032 28138 8044
rect 28261 8041 28273 8044
rect 28307 8041 28319 8075
rect 28261 8035 28319 8041
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 32401 8075 32459 8081
rect 32401 8072 32413 8075
rect 32364 8044 32413 8072
rect 32364 8032 32370 8044
rect 32401 8041 32413 8044
rect 32447 8041 32459 8075
rect 32401 8035 32459 8041
rect 7116 7908 8248 7936
rect 7116 7877 7144 7908
rect 8220 7880 8248 7908
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 7331 7840 8156 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 8128 7812 8156 7840
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 8260 7840 9781 7868
rect 8260 7828 8266 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 20714 7868 20720 7880
rect 19475 7840 20720 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 7374 7800 7380 7812
rect 7335 7772 7380 7800
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 9968 7800 9996 7831
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 24026 7828 24032 7880
rect 24084 7868 24090 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24084 7840 24593 7868
rect 24084 7828 24090 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 28537 7871 28595 7877
rect 28537 7837 28549 7871
rect 28583 7868 28595 7871
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 28583 7840 29745 7868
rect 28583 7837 28595 7840
rect 28537 7831 28595 7837
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 33686 7868 33692 7880
rect 33647 7840 33692 7868
rect 29733 7831 29791 7837
rect 33686 7828 33692 7840
rect 33744 7828 33750 7880
rect 8168 7772 9996 7800
rect 10137 7803 10195 7809
rect 8168 7760 8174 7772
rect 10137 7769 10149 7803
rect 10183 7800 10195 7803
rect 10226 7800 10232 7812
rect 10183 7772 10232 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 15930 7760 15936 7812
rect 15988 7800 15994 7812
rect 16301 7803 16359 7809
rect 16301 7800 16313 7803
rect 15988 7772 16313 7800
rect 15988 7760 15994 7772
rect 16301 7769 16313 7772
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 21637 7803 21695 7809
rect 21637 7800 21649 7803
rect 20864 7772 21649 7800
rect 20864 7760 20870 7772
rect 21637 7769 21649 7772
rect 21683 7769 21695 7803
rect 28074 7800 28080 7812
rect 28035 7772 28080 7800
rect 21637 7763 21695 7769
rect 28074 7760 28080 7772
rect 28132 7760 28138 7812
rect 28261 7803 28319 7809
rect 28261 7769 28273 7803
rect 28307 7800 28319 7803
rect 28350 7800 28356 7812
rect 28307 7772 28356 7800
rect 28307 7769 28319 7772
rect 28261 7763 28319 7769
rect 28350 7760 28356 7772
rect 28408 7760 28414 7812
rect 17586 7732 17592 7744
rect 17547 7704 17592 7732
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 20438 7692 20444 7744
rect 20496 7732 20502 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 20496 7704 20729 7732
rect 20496 7692 20502 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 20717 7695 20775 7701
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 25869 7735 25927 7741
rect 25869 7732 25881 7735
rect 23440 7704 25881 7732
rect 23440 7692 23446 7704
rect 25869 7701 25881 7704
rect 25915 7701 25927 7735
rect 25869 7695 25927 7701
rect 30374 7692 30380 7744
rect 30432 7732 30438 7744
rect 31021 7735 31079 7741
rect 31021 7732 31033 7735
rect 30432 7704 31033 7732
rect 30432 7692 30438 7704
rect 31021 7701 31033 7704
rect 31067 7701 31079 7735
rect 31021 7695 31079 7701
rect 1104 7642 35027 7664
rect 1104 7590 9390 7642
rect 9442 7590 9454 7642
rect 9506 7590 9518 7642
rect 9570 7590 9582 7642
rect 9634 7590 9646 7642
rect 9698 7590 17831 7642
rect 17883 7590 17895 7642
rect 17947 7590 17959 7642
rect 18011 7590 18023 7642
rect 18075 7590 18087 7642
rect 18139 7590 26272 7642
rect 26324 7590 26336 7642
rect 26388 7590 26400 7642
rect 26452 7590 26464 7642
rect 26516 7590 26528 7642
rect 26580 7590 34713 7642
rect 34765 7590 34777 7642
rect 34829 7590 34841 7642
rect 34893 7590 34905 7642
rect 34957 7590 34969 7642
rect 35021 7590 35027 7642
rect 1104 7568 35027 7590
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 10560 7500 10701 7528
rect 10560 7488 10566 7500
rect 10689 7497 10701 7500
rect 10735 7528 10747 7531
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 10735 7500 12173 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 15930 7528 15936 7540
rect 15891 7500 15936 7528
rect 12161 7491 12219 7497
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 17402 7488 17408 7540
rect 17460 7528 17466 7540
rect 19518 7528 19524 7540
rect 17460 7500 18920 7528
rect 19479 7500 19524 7528
rect 17460 7488 17466 7500
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 5684 7432 6837 7460
rect 5684 7420 5690 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 7374 7420 7380 7472
rect 7432 7420 7438 7472
rect 10226 7420 10232 7472
rect 10284 7420 10290 7472
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 15565 7463 15623 7469
rect 15565 7460 15577 7463
rect 15252 7432 15577 7460
rect 15252 7420 15258 7432
rect 15565 7429 15577 7432
rect 15611 7429 15623 7463
rect 15565 7423 15623 7429
rect 15749 7463 15807 7469
rect 15749 7429 15761 7463
rect 15795 7460 15807 7463
rect 16666 7460 16672 7472
rect 15795 7432 16672 7460
rect 15795 7429 15807 7432
rect 15749 7423 15807 7429
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 17586 7460 17592 7472
rect 17420 7432 17592 7460
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3786 7392 3792 7404
rect 2731 7364 3792 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8938 7392 8944 7404
rect 8444 7364 8944 7392
rect 8444 7352 8450 7364
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 17420 7392 17448 7432
rect 17586 7420 17592 7432
rect 17644 7460 17650 7472
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 17644 7432 18245 7460
rect 17644 7420 17650 7432
rect 18233 7429 18245 7432
rect 18279 7429 18291 7463
rect 18892 7460 18920 7500
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 20625 7531 20683 7537
rect 20625 7528 20637 7531
rect 20588 7500 20637 7528
rect 20588 7488 20594 7500
rect 20625 7497 20637 7500
rect 20671 7497 20683 7531
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20625 7491 20683 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 22373 7531 22431 7537
rect 22373 7528 22385 7531
rect 21048 7500 22385 7528
rect 21048 7488 21054 7500
rect 22373 7497 22385 7500
rect 22419 7497 22431 7531
rect 25958 7528 25964 7540
rect 25919 7500 25964 7528
rect 22373 7491 22431 7497
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 29086 7528 29092 7540
rect 29047 7500 29092 7528
rect 29086 7488 29092 7500
rect 29144 7488 29150 7540
rect 20438 7460 20444 7472
rect 18892 7432 20444 7460
rect 18233 7423 18291 7429
rect 20438 7420 20444 7432
rect 20496 7420 20502 7472
rect 20898 7420 20904 7472
rect 20956 7460 20962 7472
rect 23382 7460 23388 7472
rect 20956 7432 22508 7460
rect 23343 7432 23388 7460
rect 20956 7420 20962 7432
rect 14783 7364 17448 7392
rect 17497 7395 17555 7401
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 17497 7361 17509 7395
rect 17543 7361 17555 7395
rect 17678 7392 17684 7404
rect 17639 7364 17684 7392
rect 17497 7355 17555 7361
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 8404 7324 8432 7352
rect 6595 7296 8432 7324
rect 9217 7327 9275 7333
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 11054 7324 11060 7336
rect 9263 7296 11060 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 11296 7296 11897 7324
rect 11296 7284 11302 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 11885 7287 11943 7293
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7324 12127 7327
rect 13078 7324 13084 7336
rect 12115 7296 13084 7324
rect 12115 7293 12127 7296
rect 12069 7287 12127 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 17034 7284 17040 7336
rect 17092 7324 17098 7336
rect 17512 7324 17540 7355
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7392 17831 7395
rect 17862 7392 17868 7404
rect 17819 7364 17868 7392
rect 17819 7361 17831 7364
rect 17773 7355 17831 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22370 7392 22376 7404
rect 22235 7364 22376 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 22480 7401 22508 7432
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 25038 7460 25044 7472
rect 24999 7432 25044 7460
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 29362 7460 29368 7472
rect 25792 7432 29368 7460
rect 25792 7401 25820 7432
rect 29362 7420 29368 7432
rect 29420 7420 29426 7472
rect 22465 7395 22523 7401
rect 22465 7361 22477 7395
rect 22511 7361 22523 7395
rect 25777 7395 25835 7401
rect 25777 7392 25789 7395
rect 22465 7355 22523 7361
rect 23952 7364 25789 7392
rect 22388 7324 22416 7352
rect 23750 7324 23756 7336
rect 17092 7296 22094 7324
rect 22388 7296 23756 7324
rect 17092 7284 17098 7296
rect 21726 7256 21732 7268
rect 20640 7228 21732 7256
rect 2590 7188 2596 7200
rect 2551 7160 2596 7188
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 12526 7188 12532 7200
rect 12487 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 15102 7188 15108 7200
rect 13495 7160 15108 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15654 7148 15660 7200
rect 15712 7188 15718 7200
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15712 7160 15761 7188
rect 15712 7148 15718 7160
rect 15749 7157 15761 7160
rect 15795 7188 15807 7191
rect 19426 7188 19432 7200
rect 15795 7160 19432 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 19426 7148 19432 7160
rect 19484 7188 19490 7200
rect 20640 7197 20668 7228
rect 21726 7216 21732 7228
rect 21784 7216 21790 7268
rect 22066 7256 22094 7296
rect 23750 7284 23756 7296
rect 23808 7284 23814 7336
rect 23952 7256 23980 7364
rect 25777 7361 25789 7364
rect 25823 7361 25835 7395
rect 26050 7392 26056 7404
rect 25963 7364 26056 7392
rect 25777 7355 25835 7361
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 30374 7392 30380 7404
rect 30335 7364 30380 7392
rect 30374 7352 30380 7364
rect 30432 7352 30438 7404
rect 24026 7284 24032 7336
rect 24084 7324 24090 7336
rect 24578 7324 24584 7336
rect 24084 7296 24584 7324
rect 24084 7284 24090 7296
rect 24578 7284 24584 7296
rect 24636 7324 24642 7336
rect 26068 7324 26096 7352
rect 24636 7296 26096 7324
rect 24636 7284 24642 7296
rect 22066 7228 23980 7256
rect 20625 7191 20683 7197
rect 20625 7188 20637 7191
rect 19484 7160 20637 7188
rect 19484 7148 19490 7160
rect 20625 7157 20637 7160
rect 20671 7157 20683 7191
rect 20625 7151 20683 7157
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 22005 7191 22063 7197
rect 22005 7188 22017 7191
rect 20772 7160 22017 7188
rect 20772 7148 20778 7160
rect 22005 7157 22017 7160
rect 22051 7157 22063 7191
rect 25590 7188 25596 7200
rect 25551 7160 25596 7188
rect 22005 7151 22063 7157
rect 25590 7148 25596 7160
rect 25648 7148 25654 7200
rect 1104 7098 34868 7120
rect 1104 7046 5170 7098
rect 5222 7046 5234 7098
rect 5286 7046 5298 7098
rect 5350 7046 5362 7098
rect 5414 7046 5426 7098
rect 5478 7046 13611 7098
rect 13663 7046 13675 7098
rect 13727 7046 13739 7098
rect 13791 7046 13803 7098
rect 13855 7046 13867 7098
rect 13919 7046 22052 7098
rect 22104 7046 22116 7098
rect 22168 7046 22180 7098
rect 22232 7046 22244 7098
rect 22296 7046 22308 7098
rect 22360 7046 30493 7098
rect 30545 7046 30557 7098
rect 30609 7046 30621 7098
rect 30673 7046 30685 7098
rect 30737 7046 30749 7098
rect 30801 7046 34868 7098
rect 1104 7024 34868 7046
rect 1844 6987 1902 6993
rect 1844 6953 1856 6987
rect 1890 6984 1902 6987
rect 2590 6984 2596 6996
rect 1890 6956 2596 6984
rect 1890 6953 1902 6956
rect 1844 6947 1902 6953
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 13078 6984 13084 6996
rect 13039 6956 13084 6984
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 20346 6984 20352 6996
rect 19306 6956 20352 6984
rect 17862 6916 17868 6928
rect 17512 6888 17868 6916
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 3142 6848 3148 6860
rect 1627 6820 3148 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 3786 6848 3792 6860
rect 3375 6820 3792 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 5074 6848 5080 6860
rect 4396 6820 5080 6848
rect 4396 6808 4402 6820
rect 5074 6808 5080 6820
rect 5132 6848 5138 6860
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5132 6820 5457 6848
rect 5132 6808 5138 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 5718 6789 5724 6792
rect 5712 6780 5724 6789
rect 5679 6752 5724 6780
rect 5712 6743 5724 6752
rect 5718 6740 5724 6743
rect 5776 6740 5782 6792
rect 2866 6672 2872 6724
rect 2924 6672 2930 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 6840 6684 7757 6712
rect 6840 6653 6868 6684
rect 7745 6681 7757 6684
rect 7791 6681 7803 6715
rect 7944 6712 7972 6811
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 8352 6820 10149 6848
rect 8352 6808 8358 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10686 6848 10692 6860
rect 10647 6820 10692 6848
rect 10137 6811 10195 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15160 6820 15577 6848
rect 15160 6808 15166 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6780 10287 6783
rect 10410 6780 10416 6792
rect 10275 6752 10416 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 10502 6740 10508 6792
rect 10560 6789 10566 6792
rect 10560 6783 10609 6789
rect 10560 6749 10563 6783
rect 10597 6749 10609 6783
rect 11238 6780 11244 6792
rect 10560 6743 10609 6749
rect 10704 6752 11244 6780
rect 10560 6740 10566 6743
rect 10704 6712 10732 6752
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 15654 6780 15660 6792
rect 13771 6752 15660 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 7944 6684 10732 6712
rect 7745 6675 7803 6681
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11946 6715 12004 6721
rect 11946 6712 11958 6715
rect 11112 6684 11958 6712
rect 11112 6672 11118 6684
rect 11946 6681 11958 6684
rect 11992 6681 12004 6715
rect 12802 6712 12808 6724
rect 11946 6675 12004 6681
rect 12406 6684 12808 6712
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 6972 6616 7297 6644
rect 6972 6604 6978 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 8294 6644 8300 6656
rect 7699 6616 8300 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 12406 6644 12434 6684
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 13556 6712 13584 6743
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 17218 6780 17224 6792
rect 15764 6752 17224 6780
rect 15764 6712 15792 6752
rect 17218 6740 17224 6752
rect 17276 6780 17282 6792
rect 17512 6780 17540 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 19306 6848 19334 6956
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 21266 6848 21272 6860
rect 17604 6820 19334 6848
rect 21227 6820 21272 6848
rect 17604 6789 17632 6820
rect 21266 6808 21272 6820
rect 21324 6808 21330 6860
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 22704 6820 23980 6848
rect 22704 6808 22710 6820
rect 17276 6752 17540 6780
rect 17589 6783 17647 6789
rect 17276 6740 17282 6752
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17589 6743 17647 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19518 6780 19524 6792
rect 19475 6752 19524 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19702 6789 19708 6792
rect 19696 6780 19708 6789
rect 19663 6752 19708 6780
rect 19696 6743 19708 6752
rect 19702 6740 19708 6743
rect 19760 6740 19766 6792
rect 21536 6783 21594 6789
rect 21536 6749 21548 6783
rect 21582 6780 21594 6783
rect 21818 6780 21824 6792
rect 21582 6752 21824 6780
rect 21582 6749 21594 6752
rect 21536 6743 21594 6749
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 23750 6780 23756 6792
rect 23711 6752 23756 6780
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 23952 6789 23980 6820
rect 23937 6783 23995 6789
rect 23937 6749 23949 6783
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 24026 6740 24032 6792
rect 24084 6780 24090 6792
rect 24581 6783 24639 6789
rect 24084 6752 24129 6780
rect 24084 6740 24090 6752
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24627 6752 25084 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 25056 6724 25084 6752
rect 28902 6740 28908 6792
rect 28960 6789 28966 6792
rect 28960 6780 28972 6789
rect 28960 6752 29005 6780
rect 28960 6743 28972 6752
rect 28960 6740 28966 6743
rect 29086 6740 29092 6792
rect 29144 6780 29150 6792
rect 29181 6783 29239 6789
rect 29181 6780 29193 6783
rect 29144 6752 29193 6780
rect 29144 6740 29150 6752
rect 29181 6749 29193 6752
rect 29227 6749 29239 6783
rect 29181 6743 29239 6749
rect 29822 6740 29828 6792
rect 29880 6780 29886 6792
rect 30101 6783 30159 6789
rect 30101 6780 30113 6783
rect 29880 6752 30113 6780
rect 29880 6740 29886 6752
rect 30101 6749 30113 6752
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 13556 6684 15792 6712
rect 15832 6715 15890 6721
rect 15832 6681 15844 6715
rect 15878 6712 15890 6715
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 15878 6684 17417 6712
rect 15878 6681 15890 6684
rect 15832 6675 15890 6681
rect 17405 6681 17417 6684
rect 17451 6681 17463 6715
rect 17405 6675 17463 6681
rect 17494 6672 17500 6724
rect 17552 6712 17558 6724
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 17552 6684 17785 6712
rect 17552 6672 17558 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 24848 6715 24906 6721
rect 24848 6681 24860 6715
rect 24894 6712 24906 6715
rect 24946 6712 24952 6724
rect 24894 6684 24952 6712
rect 24894 6681 24906 6684
rect 24848 6675 24906 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 25038 6672 25044 6724
rect 25096 6672 25102 6724
rect 28258 6712 28264 6724
rect 27816 6684 28264 6712
rect 13630 6644 13636 6656
rect 11011 6616 12434 6644
rect 13591 6616 13636 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 16945 6647 17003 6653
rect 16945 6613 16957 6647
rect 16991 6644 17003 6647
rect 17512 6644 17540 6672
rect 16991 6616 17540 6644
rect 16991 6613 17003 6616
rect 16945 6607 17003 6613
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 18380 6616 20821 6644
rect 18380 6604 18386 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 22649 6647 22707 6653
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 22830 6644 22836 6656
rect 22695 6616 22836 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 23566 6644 23572 6656
rect 23527 6616 23572 6644
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 25866 6604 25872 6656
rect 25924 6644 25930 6656
rect 27816 6653 27844 6684
rect 28258 6672 28264 6684
rect 28316 6672 28322 6724
rect 29270 6672 29276 6724
rect 29328 6712 29334 6724
rect 30346 6715 30404 6721
rect 30346 6712 30358 6715
rect 29328 6684 30358 6712
rect 29328 6672 29334 6684
rect 30346 6681 30358 6684
rect 30392 6681 30404 6715
rect 30346 6675 30404 6681
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25924 6616 25973 6644
rect 25924 6604 25930 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 27801 6647 27859 6653
rect 27801 6613 27813 6647
rect 27847 6613 27859 6647
rect 27801 6607 27859 6613
rect 27890 6604 27896 6656
rect 27948 6644 27954 6656
rect 31481 6647 31539 6653
rect 31481 6644 31493 6647
rect 27948 6616 31493 6644
rect 27948 6604 27954 6616
rect 31481 6613 31493 6616
rect 31527 6613 31539 6647
rect 31481 6607 31539 6613
rect 1104 6554 35027 6576
rect 1104 6502 9390 6554
rect 9442 6502 9454 6554
rect 9506 6502 9518 6554
rect 9570 6502 9582 6554
rect 9634 6502 9646 6554
rect 9698 6502 17831 6554
rect 17883 6502 17895 6554
rect 17947 6502 17959 6554
rect 18011 6502 18023 6554
rect 18075 6502 18087 6554
rect 18139 6502 26272 6554
rect 26324 6502 26336 6554
rect 26388 6502 26400 6554
rect 26452 6502 26464 6554
rect 26516 6502 26528 6554
rect 26580 6502 34713 6554
rect 34765 6502 34777 6554
rect 34829 6502 34841 6554
rect 34893 6502 34905 6554
rect 34957 6502 34969 6554
rect 35021 6502 35027 6554
rect 1104 6480 35027 6502
rect 2866 6400 2872 6452
rect 2924 6400 2930 6452
rect 6914 6440 6920 6452
rect 6875 6412 6920 6440
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 12989 6443 13047 6449
rect 12989 6440 13001 6443
rect 12584 6412 13001 6440
rect 12584 6400 12590 6412
rect 12989 6409 13001 6412
rect 13035 6409 13047 6443
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 12989 6403 13047 6409
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 28258 6400 28264 6452
rect 28316 6440 28322 6452
rect 30834 6440 30840 6452
rect 28316 6412 30840 6440
rect 28316 6400 28322 6412
rect 30834 6400 30840 6412
rect 30892 6400 30898 6452
rect 2777 6375 2835 6381
rect 2777 6341 2789 6375
rect 2823 6372 2835 6375
rect 2884 6372 2912 6400
rect 2823 6344 2912 6372
rect 3697 6375 3755 6381
rect 2823 6341 2835 6344
rect 2777 6335 2835 6341
rect 3697 6341 3709 6375
rect 3743 6372 3755 6375
rect 3786 6372 3792 6384
rect 3743 6344 3792 6372
rect 3743 6341 3755 6344
rect 3697 6335 3755 6341
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 7006 6372 7012 6384
rect 6871 6344 7012 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 12897 6375 12955 6381
rect 12897 6341 12909 6375
rect 12943 6372 12955 6375
rect 13630 6372 13636 6384
rect 12943 6344 13636 6372
rect 12943 6341 12955 6344
rect 12897 6335 12955 6341
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 19880 6375 19938 6381
rect 19880 6341 19892 6375
rect 19926 6372 19938 6375
rect 20714 6372 20720 6384
rect 19926 6344 20720 6372
rect 19926 6341 19938 6344
rect 19880 6335 19938 6341
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 24682 6375 24740 6381
rect 24682 6372 24694 6375
rect 23624 6344 24694 6372
rect 23624 6332 23630 6344
rect 24682 6341 24694 6344
rect 24728 6341 24740 6375
rect 24682 6335 24740 6341
rect 29178 6332 29184 6384
rect 29236 6372 29242 6384
rect 29558 6375 29616 6381
rect 29558 6372 29570 6375
rect 29236 6344 29570 6372
rect 29236 6332 29242 6344
rect 29558 6341 29570 6344
rect 29604 6341 29616 6375
rect 29558 6335 29616 6341
rect 2958 6304 2964 6316
rect 2919 6276 2964 6304
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3142 6304 3148 6316
rect 3055 6276 3148 6304
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3160 6236 3188 6264
rect 4062 6236 4068 6248
rect 3160 6208 4068 6236
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6144 6208 6653 6236
rect 6144 6196 6150 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12492 6208 12725 6236
rect 12492 6196 12498 6208
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19576 6208 19625 6236
rect 19576 6196 19582 6208
rect 19613 6205 19625 6208
rect 19659 6205 19671 6239
rect 19613 6199 19671 6205
rect 24949 6239 25007 6245
rect 24949 6205 24961 6239
rect 24995 6205 25007 6239
rect 29822 6236 29828 6248
rect 29783 6208 29828 6236
rect 24949 6199 25007 6205
rect 7285 6171 7343 6177
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 18414 6168 18420 6180
rect 7331 6140 18420 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 18414 6128 18420 6140
rect 18472 6128 18478 6180
rect 22646 6128 22652 6180
rect 22704 6168 22710 6180
rect 23569 6171 23627 6177
rect 23569 6168 23581 6171
rect 22704 6140 23581 6168
rect 22704 6128 22710 6140
rect 23569 6137 23581 6140
rect 23615 6137 23627 6171
rect 23569 6131 23627 6137
rect 3789 6103 3847 6109
rect 3789 6069 3801 6103
rect 3835 6100 3847 6103
rect 3970 6100 3976 6112
rect 3835 6072 3976 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 13357 6103 13415 6109
rect 13357 6069 13369 6103
rect 13403 6100 13415 6103
rect 19978 6100 19984 6112
rect 13403 6072 19984 6100
rect 13403 6069 13415 6072
rect 13357 6063 13415 6069
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 24964 6100 24992 6199
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 28445 6171 28503 6177
rect 28445 6137 28457 6171
rect 28491 6168 28503 6171
rect 28810 6168 28816 6180
rect 28491 6140 28816 6168
rect 28491 6137 28503 6140
rect 28445 6131 28503 6137
rect 28810 6128 28816 6140
rect 28868 6128 28874 6180
rect 24728 6072 24992 6100
rect 24728 6060 24734 6072
rect 1104 6010 34868 6032
rect 1104 5958 5170 6010
rect 5222 5958 5234 6010
rect 5286 5958 5298 6010
rect 5350 5958 5362 6010
rect 5414 5958 5426 6010
rect 5478 5958 13611 6010
rect 13663 5958 13675 6010
rect 13727 5958 13739 6010
rect 13791 5958 13803 6010
rect 13855 5958 13867 6010
rect 13919 5958 22052 6010
rect 22104 5958 22116 6010
rect 22168 5958 22180 6010
rect 22232 5958 22244 6010
rect 22296 5958 22308 6010
rect 22360 5958 30493 6010
rect 30545 5958 30557 6010
rect 30609 5958 30621 6010
rect 30673 5958 30685 6010
rect 30737 5958 30749 6010
rect 30801 5958 34868 6010
rect 1104 5936 34868 5958
rect 25958 5896 25964 5908
rect 25919 5868 25964 5896
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 29181 5899 29239 5905
rect 29181 5865 29193 5899
rect 29227 5896 29239 5899
rect 29270 5896 29276 5908
rect 29227 5868 29276 5896
rect 29227 5865 29239 5868
rect 29181 5859 29239 5865
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 28994 5828 29000 5840
rect 28736 5800 29000 5828
rect 3970 5760 3976 5772
rect 3931 5732 3976 5760
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 5626 5760 5632 5772
rect 4387 5732 5632 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5692 24639 5695
rect 24670 5692 24676 5704
rect 24627 5664 24676 5692
rect 24627 5661 24639 5664
rect 24581 5655 24639 5661
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 24848 5695 24906 5701
rect 24848 5661 24860 5695
rect 24894 5692 24906 5695
rect 25590 5692 25596 5704
rect 24894 5664 25596 5692
rect 24894 5661 24906 5664
rect 24848 5655 24906 5661
rect 25590 5652 25596 5664
rect 25648 5652 25654 5704
rect 28736 5701 28764 5800
rect 28994 5788 29000 5800
rect 29052 5788 29058 5840
rect 28721 5695 28779 5701
rect 28721 5661 28733 5695
rect 28767 5661 28779 5695
rect 28721 5655 28779 5661
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 29362 5692 29368 5704
rect 29043 5664 29368 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 29362 5652 29368 5664
rect 29420 5652 29426 5704
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 8202 5624 8208 5636
rect 5460 5596 8208 5624
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 5460 5556 5488 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 27890 5584 27896 5636
rect 27948 5624 27954 5636
rect 28813 5627 28871 5633
rect 28813 5624 28825 5627
rect 27948 5596 28825 5624
rect 27948 5584 27954 5596
rect 28813 5593 28825 5596
rect 28859 5593 28871 5627
rect 28813 5587 28871 5593
rect 6086 5556 6092 5568
rect 4120 5528 5488 5556
rect 6047 5528 6092 5556
rect 4120 5516 4126 5528
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 1104 5466 35027 5488
rect 1104 5414 9390 5466
rect 9442 5414 9454 5466
rect 9506 5414 9518 5466
rect 9570 5414 9582 5466
rect 9634 5414 9646 5466
rect 9698 5414 17831 5466
rect 17883 5414 17895 5466
rect 17947 5414 17959 5466
rect 18011 5414 18023 5466
rect 18075 5414 18087 5466
rect 18139 5414 26272 5466
rect 26324 5414 26336 5466
rect 26388 5414 26400 5466
rect 26452 5414 26464 5466
rect 26516 5414 26528 5466
rect 26580 5414 34713 5466
rect 34765 5414 34777 5466
rect 34829 5414 34841 5466
rect 34893 5414 34905 5466
rect 34957 5414 34969 5466
rect 35021 5414 35027 5466
rect 1104 5392 35027 5414
rect 5626 5352 5632 5364
rect 5587 5324 5632 5352
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 10502 5352 10508 5364
rect 6144 5324 9628 5352
rect 10463 5324 10508 5352
rect 6144 5312 6150 5324
rect 2958 5244 2964 5296
rect 3016 5284 3022 5296
rect 4341 5287 4399 5293
rect 3016 5256 4292 5284
rect 3016 5244 3022 5256
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4264 5225 4292 5256
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 4706 5284 4712 5296
rect 4387 5256 4712 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 5721 5219 5779 5225
rect 4295 5188 5488 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 5460 5012 5488 5188
rect 5721 5185 5733 5219
rect 5767 5216 5779 5219
rect 6104 5216 6132 5312
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 9493 5287 9551 5293
rect 9493 5284 9505 5287
rect 9364 5256 9505 5284
rect 9364 5244 9370 5256
rect 9493 5253 9505 5256
rect 9539 5253 9551 5287
rect 9600 5284 9628 5324
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 19518 5352 19524 5364
rect 13228 5324 13952 5352
rect 19479 5324 19524 5352
rect 13228 5312 13234 5324
rect 12434 5284 12440 5296
rect 9600 5256 12440 5284
rect 9493 5247 9551 5253
rect 12434 5244 12440 5256
rect 12492 5284 12498 5296
rect 12492 5256 13584 5284
rect 12492 5244 12498 5256
rect 5767 5188 6132 5216
rect 9585 5219 9643 5225
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 6546 5148 6552 5160
rect 5684 5120 6552 5148
rect 5684 5108 5690 5120
rect 6546 5108 6552 5120
rect 6604 5148 6610 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 6604 5120 9321 5148
rect 6604 5108 6610 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9600 5148 9628 5179
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9916 5188 10425 5216
rect 9916 5176 9922 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10870 5216 10876 5228
rect 10643 5188 10876 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 13556 5225 13584 5256
rect 11957 5219 12015 5225
rect 11957 5216 11969 5219
rect 11848 5188 11969 5216
rect 11848 5176 11854 5188
rect 11957 5185 11969 5188
rect 12003 5185 12015 5219
rect 11957 5179 12015 5185
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 10686 5148 10692 5160
rect 9600 5120 10692 5148
rect 9309 5111 9367 5117
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 11698 5148 11704 5160
rect 11611 5120 11704 5148
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 11716 5080 11744 5108
rect 13832 5080 13860 5111
rect 7248 5052 11744 5080
rect 13004 5052 13860 5080
rect 13924 5080 13952 5324
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 18230 5284 18236 5296
rect 18191 5256 18236 5284
rect 18230 5244 18236 5256
rect 18288 5244 18294 5296
rect 23382 5284 23388 5296
rect 23343 5256 23388 5284
rect 23382 5244 23388 5256
rect 23440 5244 23446 5296
rect 15194 5216 15200 5228
rect 15155 5188 15200 5216
rect 15194 5176 15200 5188
rect 15252 5216 15258 5228
rect 17402 5216 17408 5228
rect 15252 5188 17408 5216
rect 15252 5176 15258 5188
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 25774 5216 25780 5228
rect 25735 5188 25780 5216
rect 25774 5176 25780 5188
rect 25832 5176 25838 5228
rect 25961 5219 26019 5225
rect 25961 5185 25973 5219
rect 26007 5185 26019 5219
rect 25961 5179 26019 5185
rect 25976 5148 26004 5179
rect 26602 5148 26608 5160
rect 25056 5120 26608 5148
rect 25056 5092 25084 5120
rect 26602 5108 26608 5120
rect 26660 5108 26666 5160
rect 25038 5080 25044 5092
rect 13924 5052 25044 5080
rect 7248 5040 7254 5052
rect 8110 5012 8116 5024
rect 5460 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 9950 5012 9956 5024
rect 9911 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 11974 5012 11980 5024
rect 11296 4984 11980 5012
rect 11296 4972 11302 4984
rect 11974 4972 11980 4984
rect 12032 5012 12038 5024
rect 13004 5012 13032 5052
rect 25038 5040 25044 5052
rect 25096 5040 25102 5092
rect 12032 4984 13032 5012
rect 13081 5015 13139 5021
rect 12032 4972 12038 4984
rect 13081 4981 13093 5015
rect 13127 5012 13139 5015
rect 13633 5015 13691 5021
rect 13633 5012 13645 5015
rect 13127 4984 13645 5012
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 13633 4981 13645 4984
rect 13679 4981 13691 5015
rect 13633 4975 13691 4981
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 14274 5012 14280 5024
rect 13771 4984 14280 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 14918 4972 14924 5024
rect 14976 5012 14982 5024
rect 15105 5015 15163 5021
rect 15105 5012 15117 5015
rect 14976 4984 15117 5012
rect 14976 4972 14982 4984
rect 15105 4981 15117 4984
rect 15151 4981 15163 5015
rect 15105 4975 15163 4981
rect 25593 5015 25651 5021
rect 25593 4981 25605 5015
rect 25639 5012 25651 5015
rect 25682 5012 25688 5024
rect 25639 4984 25688 5012
rect 25639 4981 25651 4984
rect 25593 4975 25651 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 1104 4922 34868 4944
rect 1104 4870 5170 4922
rect 5222 4870 5234 4922
rect 5286 4870 5298 4922
rect 5350 4870 5362 4922
rect 5414 4870 5426 4922
rect 5478 4870 13611 4922
rect 13663 4870 13675 4922
rect 13727 4870 13739 4922
rect 13791 4870 13803 4922
rect 13855 4870 13867 4922
rect 13919 4870 22052 4922
rect 22104 4870 22116 4922
rect 22168 4870 22180 4922
rect 22232 4870 22244 4922
rect 22296 4870 22308 4922
rect 22360 4870 30493 4922
rect 30545 4870 30557 4922
rect 30609 4870 30621 4922
rect 30673 4870 30685 4922
rect 30737 4870 30749 4922
rect 30801 4870 34868 4922
rect 1104 4848 34868 4870
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11974 4808 11980 4820
rect 11935 4780 11980 4808
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 7190 4672 7196 4684
rect 5132 4644 7196 4672
rect 5132 4632 5138 4644
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 8938 4632 8944 4684
rect 8996 4672 9002 4684
rect 9125 4675 9183 4681
rect 9125 4672 9137 4675
rect 8996 4644 9137 4672
rect 8996 4632 9002 4644
rect 9125 4641 9137 4644
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 9447 4644 10824 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 7466 4613 7472 4616
rect 7460 4604 7472 4613
rect 7427 4576 7472 4604
rect 7460 4567 7472 4576
rect 7466 4564 7472 4567
rect 7524 4564 7530 4616
rect 10502 4564 10508 4616
rect 10560 4564 10566 4616
rect 10796 4536 10824 4644
rect 10888 4604 10916 4768
rect 14553 4743 14611 4749
rect 14553 4709 14565 4743
rect 14599 4740 14611 4743
rect 20714 4740 20720 4752
rect 14599 4712 20720 4740
rect 14599 4709 14611 4712
rect 14553 4703 14611 4709
rect 20714 4700 20720 4712
rect 20772 4700 20778 4752
rect 24670 4740 24676 4752
rect 24631 4712 24676 4740
rect 24670 4700 24676 4712
rect 24728 4700 24734 4752
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 14240 4644 16221 4672
rect 14240 4632 14246 4644
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 10888 4576 11897 4604
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 12434 4604 12440 4616
rect 12299 4576 12440 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14568 4613 14596 4644
rect 16209 4641 16221 4644
rect 16255 4672 16267 4675
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 16255 4644 18705 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 18693 4641 18705 4644
rect 18739 4672 18751 4675
rect 20438 4672 20444 4684
rect 18739 4644 20444 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 25038 4672 25044 4684
rect 24999 4644 25044 4672
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 15838 4564 15844 4616
rect 15896 4604 15902 4616
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 15896 4576 15945 4604
rect 15896 4564 15902 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 15933 4567 15991 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 19978 4564 19984 4616
rect 20036 4604 20042 4616
rect 20165 4607 20223 4613
rect 20165 4604 20177 4607
rect 20036 4576 20177 4604
rect 20036 4564 20042 4576
rect 20165 4573 20177 4576
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 20898 4564 20904 4616
rect 20956 4604 20962 4616
rect 21637 4607 21695 4613
rect 21637 4604 21649 4607
rect 20956 4576 21649 4604
rect 20956 4564 20962 4576
rect 21637 4573 21649 4576
rect 21683 4604 21695 4607
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 21683 4576 22293 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 22281 4573 22293 4576
rect 22327 4604 22339 4607
rect 25866 4604 25872 4616
rect 22327 4576 25872 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 25866 4564 25872 4576
rect 25924 4564 25930 4616
rect 11790 4536 11796 4548
rect 10796 4508 11796 4536
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 26142 4545 26148 4548
rect 26136 4499 26148 4545
rect 26200 4536 26206 4548
rect 26200 4508 26236 4536
rect 26142 4496 26148 4499
rect 26200 4496 26206 4508
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 9766 4468 9772 4480
rect 8619 4440 9772 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 12437 4471 12495 4477
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 14369 4471 14427 4477
rect 14369 4468 14381 4471
rect 12483 4440 14381 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 14369 4437 14381 4440
rect 14415 4437 14427 4471
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 14369 4431 14427 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4468 16083 4471
rect 16298 4468 16304 4480
rect 16071 4440 16304 4468
rect 16071 4437 16083 4440
rect 16025 4431 16083 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 17494 4468 17500 4480
rect 17455 4440 17500 4468
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18230 4468 18236 4480
rect 18095 4440 18236 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4468 18567 4471
rect 19058 4468 19064 4480
rect 18555 4440 19064 4468
rect 18555 4437 18567 4440
rect 18509 4431 18567 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 20806 4468 20812 4480
rect 20303 4440 20812 4468
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 21542 4468 21548 4480
rect 21503 4440 21548 4468
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22189 4471 22247 4477
rect 22189 4468 22201 4471
rect 22152 4440 22201 4468
rect 22152 4428 22158 4440
rect 22189 4437 22201 4440
rect 22235 4437 22247 4471
rect 24578 4468 24584 4480
rect 24539 4440 24584 4468
rect 22189 4431 22247 4437
rect 24578 4428 24584 4440
rect 24636 4428 24642 4480
rect 26786 4428 26792 4480
rect 26844 4468 26850 4480
rect 27249 4471 27307 4477
rect 27249 4468 27261 4471
rect 26844 4440 27261 4468
rect 26844 4428 26850 4440
rect 27249 4437 27261 4440
rect 27295 4437 27307 4471
rect 27249 4431 27307 4437
rect 1104 4378 35027 4400
rect 1104 4326 9390 4378
rect 9442 4326 9454 4378
rect 9506 4326 9518 4378
rect 9570 4326 9582 4378
rect 9634 4326 9646 4378
rect 9698 4326 17831 4378
rect 17883 4326 17895 4378
rect 17947 4326 17959 4378
rect 18011 4326 18023 4378
rect 18075 4326 18087 4378
rect 18139 4326 26272 4378
rect 26324 4326 26336 4378
rect 26388 4326 26400 4378
rect 26452 4326 26464 4378
rect 26516 4326 26528 4378
rect 26580 4326 34713 4378
rect 34765 4326 34777 4378
rect 34829 4326 34841 4378
rect 34893 4326 34905 4378
rect 34957 4326 34969 4378
rect 35021 4326 35027 4378
rect 1104 4304 35027 4326
rect 9306 4264 9312 4276
rect 9267 4236 9312 4264
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9677 4267 9735 4273
rect 9677 4233 9689 4267
rect 9723 4264 9735 4267
rect 9858 4264 9864 4276
rect 9723 4236 9864 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 7377 4199 7435 4205
rect 7377 4165 7389 4199
rect 7423 4196 7435 4199
rect 7466 4196 7472 4208
rect 7423 4168 7472 4196
rect 7423 4165 7435 4168
rect 7377 4159 7435 4165
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 7926 4156 7932 4208
rect 7984 4156 7990 4208
rect 8938 4128 8944 4140
rect 8588 4100 8944 4128
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4060 7159 4063
rect 8588 4060 8616 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 7147 4032 8616 4060
rect 8849 4063 8907 4069
rect 7147 4029 7159 4032
rect 7101 4023 7159 4029
rect 8849 4029 8861 4063
rect 8895 4060 8907 4063
rect 9692 4060 9720 4227
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 22462 4264 22468 4276
rect 10008 4236 22468 4264
rect 10008 4224 10014 4236
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 26142 4264 26148 4276
rect 26103 4236 26148 4264
rect 26142 4224 26148 4236
rect 26200 4224 26206 4276
rect 13354 4196 13360 4208
rect 13315 4168 13360 4196
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 15188 4199 15246 4205
rect 15188 4165 15200 4199
rect 15234 4196 15246 4199
rect 15562 4196 15568 4208
rect 15234 4168 15568 4196
rect 15234 4165 15246 4168
rect 15188 4159 15246 4165
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 25866 4196 25872 4208
rect 17420 4168 18092 4196
rect 17420 4140 17448 4168
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10502 4128 10508 4140
rect 9824 4100 9869 4128
rect 10463 4100 10508 4128
rect 9824 4088 9830 4100
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10594 4088 10600 4140
rect 10652 4128 10658 4140
rect 10870 4128 10876 4140
rect 10652 4100 10697 4128
rect 10831 4100 10876 4128
rect 10652 4088 10658 4100
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 13998 4128 14004 4140
rect 13495 4100 14004 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17402 4128 17408 4140
rect 17083 4100 17408 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17402 4088 17408 4100
rect 17460 4088 17466 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17954 4137 17960 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17552 4100 17693 4128
rect 17552 4088 17558 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17948 4128 17960 4137
rect 17915 4100 17960 4128
rect 17681 4091 17739 4097
rect 17948 4091 17960 4100
rect 17954 4088 17960 4091
rect 18012 4088 18018 4140
rect 18064 4128 18092 4168
rect 24320 4168 25872 4196
rect 19702 4128 19708 4140
rect 18064 4100 19708 4128
rect 19702 4088 19708 4100
rect 19760 4128 19766 4140
rect 20898 4128 20904 4140
rect 19760 4100 20904 4128
rect 19760 4088 19766 4100
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 21174 4128 21180 4140
rect 21232 4137 21238 4140
rect 21144 4100 21180 4128
rect 21174 4088 21180 4100
rect 21232 4091 21244 4137
rect 21453 4131 21511 4137
rect 21453 4097 21465 4131
rect 21499 4128 21511 4131
rect 21542 4128 21548 4140
rect 21499 4100 21548 4128
rect 21499 4097 21511 4100
rect 21453 4091 21511 4097
rect 21232 4088 21238 4091
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22094 4128 22100 4140
rect 22051 4100 22100 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22278 4137 22284 4140
rect 22272 4091 22284 4137
rect 22336 4128 22342 4140
rect 24320 4137 24348 4168
rect 25866 4156 25872 4168
rect 25924 4196 25930 4208
rect 28074 4196 28080 4208
rect 25924 4168 28080 4196
rect 25924 4156 25930 4168
rect 24578 4137 24584 4140
rect 24305 4131 24363 4137
rect 22336 4100 22372 4128
rect 22278 4088 22284 4091
rect 22336 4088 22342 4100
rect 24305 4097 24317 4131
rect 24351 4097 24363 4131
rect 24572 4128 24584 4137
rect 24539 4100 24584 4128
rect 24305 4091 24363 4097
rect 24572 4091 24584 4100
rect 24578 4088 24584 4091
rect 24636 4088 24642 4140
rect 26602 4128 26608 4140
rect 26563 4100 26608 4128
rect 26602 4088 26608 4100
rect 26660 4128 26666 4140
rect 27062 4128 27068 4140
rect 26660 4100 27068 4128
rect 26660 4088 26666 4100
rect 27062 4088 27068 4100
rect 27120 4088 27126 4140
rect 27172 4137 27200 4168
rect 28074 4156 28080 4168
rect 28132 4156 28138 4208
rect 27157 4131 27215 4137
rect 27157 4097 27169 4131
rect 27203 4097 27215 4131
rect 27157 4091 27215 4097
rect 27424 4131 27482 4137
rect 27424 4097 27436 4131
rect 27470 4128 27482 4131
rect 27798 4128 27804 4140
rect 27470 4100 27804 4128
rect 27470 4097 27482 4100
rect 27424 4091 27482 4097
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 8895 4032 9720 4060
rect 9953 4063 10011 4069
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 11238 4060 11244 4072
rect 9999 4032 11244 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 14182 4060 14188 4072
rect 13679 4032 14188 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 26237 3995 26295 4001
rect 26237 3961 26249 3995
rect 26283 3992 26295 3995
rect 26283 3964 26317 3992
rect 26283 3961 26295 3964
rect 26237 3955 26295 3961
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16724 3896 16957 3924
rect 16724 3884 16730 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 19058 3924 19064 3936
rect 19019 3896 19064 3924
rect 16945 3887 17003 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 20073 3927 20131 3933
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 21082 3924 21088 3936
rect 20119 3896 21088 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 23382 3924 23388 3936
rect 23343 3896 23388 3924
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 25685 3927 25743 3933
rect 25685 3893 25697 3927
rect 25731 3924 25743 3927
rect 26252 3924 26280 3955
rect 26602 3924 26608 3936
rect 25731 3896 26608 3924
rect 25731 3893 25743 3896
rect 25685 3887 25743 3893
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 28350 3884 28356 3936
rect 28408 3924 28414 3936
rect 28537 3927 28595 3933
rect 28537 3924 28549 3927
rect 28408 3896 28549 3924
rect 28408 3884 28414 3896
rect 28537 3893 28549 3896
rect 28583 3893 28595 3927
rect 28537 3887 28595 3893
rect 1104 3834 34868 3856
rect 1104 3782 5170 3834
rect 5222 3782 5234 3834
rect 5286 3782 5298 3834
rect 5350 3782 5362 3834
rect 5414 3782 5426 3834
rect 5478 3782 13611 3834
rect 13663 3782 13675 3834
rect 13727 3782 13739 3834
rect 13791 3782 13803 3834
rect 13855 3782 13867 3834
rect 13919 3782 22052 3834
rect 22104 3782 22116 3834
rect 22168 3782 22180 3834
rect 22232 3782 22244 3834
rect 22296 3782 22308 3834
rect 22360 3782 30493 3834
rect 30545 3782 30557 3834
rect 30609 3782 30621 3834
rect 30673 3782 30685 3834
rect 30737 3782 30749 3834
rect 30801 3782 34868 3834
rect 1104 3760 34868 3782
rect 7926 3720 7932 3732
rect 7887 3692 7932 3720
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 13998 3720 14004 3732
rect 13771 3692 14004 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 16850 3680 16856 3732
rect 16908 3720 16914 3732
rect 20806 3720 20812 3732
rect 16908 3692 20392 3720
rect 20767 3692 20812 3720
rect 16908 3680 16914 3692
rect 20364 3652 20392 3692
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22370 3720 22376 3732
rect 22143 3692 22376 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 24578 3720 24584 3732
rect 24539 3692 24584 3720
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 27065 3723 27123 3729
rect 27065 3720 27077 3723
rect 24688 3692 27077 3720
rect 24688 3652 24716 3692
rect 27065 3689 27077 3692
rect 27111 3689 27123 3723
rect 27798 3720 27804 3732
rect 27759 3692 27804 3720
rect 27065 3683 27123 3689
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 26786 3652 26792 3664
rect 20364 3624 24716 3652
rect 26747 3624 26792 3652
rect 26786 3612 26792 3624
rect 26844 3612 26850 3664
rect 26881 3655 26939 3661
rect 26881 3621 26893 3655
rect 26927 3652 26939 3655
rect 26927 3624 27108 3652
rect 26927 3621 26939 3624
rect 26881 3615 26939 3621
rect 8202 3584 8208 3596
rect 7944 3556 8208 3584
rect 7944 3525 7972 3556
rect 8202 3544 8208 3556
rect 8260 3584 8266 3596
rect 10870 3584 10876 3596
rect 8260 3556 10876 3584
rect 8260 3544 8266 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 16666 3584 16672 3596
rect 16627 3556 16672 3584
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 22738 3584 22744 3596
rect 22699 3556 22744 3584
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 26142 3544 26148 3596
rect 26200 3584 26206 3596
rect 26973 3587 27031 3593
rect 26973 3584 26985 3587
rect 26200 3556 26985 3584
rect 26200 3544 26206 3556
rect 26973 3553 26985 3556
rect 27019 3553 27031 3587
rect 26973 3547 27031 3553
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 10594 3516 10600 3528
rect 8168 3488 10600 3516
rect 8168 3476 8174 3488
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 12342 3516 12348 3528
rect 12303 3488 12348 3516
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 12612 3519 12670 3525
rect 12612 3485 12624 3519
rect 12658 3516 12670 3519
rect 12986 3516 12992 3528
rect 12658 3488 12992 3516
rect 12658 3485 12670 3488
rect 12612 3479 12670 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 15654 3516 15660 3528
rect 15615 3488 15660 3516
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 19426 3516 19432 3528
rect 19387 3488 19432 3516
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 22462 3516 22468 3528
rect 22423 3488 22468 3516
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3516 22615 3519
rect 23382 3516 23388 3528
rect 22603 3488 23388 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 25682 3476 25688 3528
rect 25740 3525 25746 3528
rect 25740 3516 25752 3525
rect 25740 3488 25785 3516
rect 25740 3479 25752 3488
rect 25740 3476 25746 3479
rect 25866 3476 25872 3528
rect 25924 3516 25930 3528
rect 25961 3519 26019 3525
rect 25961 3516 25973 3519
rect 25924 3488 25973 3516
rect 25924 3476 25930 3488
rect 25961 3485 25973 3488
rect 26007 3485 26019 3519
rect 25961 3479 26019 3485
rect 26421 3519 26479 3525
rect 26421 3485 26433 3519
rect 26467 3516 26479 3519
rect 26602 3516 26608 3528
rect 26467 3488 26608 3516
rect 26467 3485 26479 3488
rect 26421 3479 26479 3485
rect 26602 3476 26608 3488
rect 26660 3476 26666 3528
rect 27080 3516 27108 3624
rect 27614 3612 27620 3664
rect 27672 3652 27678 3664
rect 27893 3655 27951 3661
rect 27893 3652 27905 3655
rect 27672 3624 27905 3652
rect 27672 3612 27678 3624
rect 27893 3621 27905 3624
rect 27939 3621 27951 3655
rect 27893 3615 27951 3621
rect 27154 3544 27160 3596
rect 27212 3584 27218 3596
rect 28261 3587 28319 3593
rect 28261 3584 28273 3587
rect 27212 3556 28273 3584
rect 27212 3544 27218 3556
rect 28261 3553 28273 3556
rect 28307 3553 28319 3587
rect 28261 3547 28319 3553
rect 28350 3516 28356 3528
rect 27080 3488 28356 3516
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 16942 3457 16948 3460
rect 15390 3451 15448 3457
rect 15390 3448 15402 3451
rect 14792 3420 15402 3448
rect 14792 3408 14798 3420
rect 15390 3417 15402 3420
rect 15436 3417 15448 3451
rect 15390 3411 15448 3417
rect 16936 3411 16948 3457
rect 17000 3448 17006 3460
rect 19696 3451 19754 3457
rect 17000 3420 17036 3448
rect 16942 3408 16948 3411
rect 17000 3408 17006 3420
rect 19696 3417 19708 3451
rect 19742 3448 19754 3451
rect 19794 3448 19800 3460
rect 19742 3420 19800 3448
rect 19742 3417 19754 3420
rect 19696 3411 19754 3417
rect 19794 3408 19800 3420
rect 19852 3408 19858 3460
rect 25774 3408 25780 3460
rect 25832 3448 25838 3460
rect 27080 3448 27108 3488
rect 28350 3476 28356 3488
rect 28408 3476 28414 3528
rect 25832 3420 27108 3448
rect 25832 3408 25838 3420
rect 14274 3380 14280 3392
rect 14235 3352 14280 3380
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 18230 3380 18236 3392
rect 18095 3352 18236 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 18230 3340 18236 3352
rect 18288 3340 18294 3392
rect 1104 3290 35027 3312
rect 1104 3238 9390 3290
rect 9442 3238 9454 3290
rect 9506 3238 9518 3290
rect 9570 3238 9582 3290
rect 9634 3238 9646 3290
rect 9698 3238 17831 3290
rect 17883 3238 17895 3290
rect 17947 3238 17959 3290
rect 18011 3238 18023 3290
rect 18075 3238 18087 3290
rect 18139 3238 26272 3290
rect 26324 3238 26336 3290
rect 26388 3238 26400 3290
rect 26452 3238 26464 3290
rect 26516 3238 26528 3290
rect 26580 3238 34713 3290
rect 34765 3238 34777 3290
rect 34829 3238 34841 3290
rect 34893 3238 34905 3290
rect 34957 3238 34969 3290
rect 35021 3238 35027 3290
rect 1104 3216 35027 3238
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12529 3179 12587 3185
rect 12529 3176 12541 3179
rect 12400 3148 12541 3176
rect 12400 3136 12406 3148
rect 12529 3145 12541 3148
rect 12575 3145 12587 3179
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 12529 3139 12587 3145
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14734 3176 14740 3188
rect 14695 3148 14740 3176
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15654 3176 15660 3188
rect 15335 3148 15660 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16942 3176 16948 3188
rect 16903 3148 16948 3176
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17184 3148 17325 3176
rect 17184 3136 17190 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 18230 3176 18236 3188
rect 17451 3148 18236 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19484 3148 19625 3176
rect 19484 3136 19490 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 19613 3139 19671 3145
rect 20717 3179 20775 3185
rect 20717 3145 20729 3179
rect 20763 3176 20775 3179
rect 21174 3176 21180 3188
rect 20763 3148 21180 3176
rect 20763 3145 20775 3148
rect 20717 3139 20775 3145
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 29089 3179 29147 3185
rect 29089 3145 29101 3179
rect 29135 3176 29147 3179
rect 29822 3176 29828 3188
rect 29135 3148 29828 3176
rect 29135 3145 29147 3148
rect 29089 3139 29147 3145
rect 29822 3136 29828 3148
rect 29880 3136 29886 3188
rect 21082 3108 21088 3120
rect 12636 3080 15240 3108
rect 21043 3080 21088 3108
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 12636 3049 12664 3080
rect 15212 3049 15240 3080
rect 21082 3068 21088 3080
rect 21140 3068 21146 3120
rect 30374 3108 30380 3120
rect 30335 3080 30380 3108
rect 30374 3068 30380 3080
rect 30432 3068 30438 3120
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 10928 3012 12633 3040
rect 10928 3000 10934 3012
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 15197 3043 15255 3049
rect 15197 3009 15209 3043
rect 15243 3009 15255 3043
rect 19702 3040 19708 3052
rect 19663 3012 19708 3040
rect 15197 3003 15255 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 20772 3012 20913 3040
rect 20772 3000 20778 3012
rect 20901 3009 20913 3012
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21177 3043 21235 3049
rect 21177 3009 21189 3043
rect 21223 3040 21235 3043
rect 22738 3040 22744 3052
rect 21223 3012 22744 3040
rect 21223 3009 21235 3012
rect 21177 3003 21235 3009
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 15470 2972 15476 2984
rect 14332 2944 15476 2972
rect 14332 2932 14338 2944
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 17589 2975 17647 2981
rect 17589 2941 17601 2975
rect 17635 2972 17647 2975
rect 20438 2972 20444 2984
rect 17635 2944 20444 2972
rect 17635 2941 17647 2944
rect 17589 2935 17647 2941
rect 20438 2932 20444 2944
rect 20496 2972 20502 2984
rect 21192 2972 21220 3003
rect 22738 3000 22744 3012
rect 22796 3040 22802 3052
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 22796 3012 25145 3040
rect 22796 3000 22802 3012
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3040 26111 3043
rect 26786 3040 26792 3052
rect 26099 3012 26792 3040
rect 26099 3009 26111 3012
rect 26053 3003 26111 3009
rect 26786 3000 26792 3012
rect 26844 3040 26850 3052
rect 27614 3040 27620 3052
rect 26844 3012 27620 3040
rect 26844 3000 26850 3012
rect 27614 3000 27620 3012
rect 27672 3000 27678 3052
rect 20496 2944 21220 2972
rect 20496 2932 20502 2944
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 25501 2975 25559 2981
rect 25501 2972 25513 2975
rect 25096 2944 25513 2972
rect 25096 2932 25102 2944
rect 25501 2941 25513 2944
rect 25547 2972 25559 2975
rect 26142 2972 26148 2984
rect 25547 2944 26148 2972
rect 25547 2941 25559 2944
rect 25501 2935 25559 2941
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 25593 2907 25651 2913
rect 25593 2873 25605 2907
rect 25639 2904 25651 2907
rect 25639 2876 26004 2904
rect 25639 2873 25651 2876
rect 25593 2867 25651 2873
rect 25685 2839 25743 2845
rect 25685 2805 25697 2839
rect 25731 2836 25743 2839
rect 25774 2836 25780 2848
rect 25731 2808 25780 2836
rect 25731 2805 25743 2808
rect 25685 2799 25743 2805
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 25976 2836 26004 2876
rect 26234 2836 26240 2848
rect 25976 2808 26240 2836
rect 26234 2796 26240 2808
rect 26292 2836 26298 2848
rect 26602 2836 26608 2848
rect 26292 2808 26608 2836
rect 26292 2796 26298 2808
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 1104 2746 34868 2768
rect 1104 2694 5170 2746
rect 5222 2694 5234 2746
rect 5286 2694 5298 2746
rect 5350 2694 5362 2746
rect 5414 2694 5426 2746
rect 5478 2694 13611 2746
rect 13663 2694 13675 2746
rect 13727 2694 13739 2746
rect 13791 2694 13803 2746
rect 13855 2694 13867 2746
rect 13919 2694 22052 2746
rect 22104 2694 22116 2746
rect 22168 2694 22180 2746
rect 22232 2694 22244 2746
rect 22296 2694 22308 2746
rect 22360 2694 30493 2746
rect 30545 2694 30557 2746
rect 30609 2694 30621 2746
rect 30673 2694 30685 2746
rect 30737 2694 30749 2746
rect 30801 2694 34868 2746
rect 1104 2672 34868 2694
rect 15930 2632 15936 2644
rect 4448 2604 15936 2632
rect 2056 2468 4384 2496
rect 2056 2437 2084 2468
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 1268 2332 1777 2360
rect 1268 2320 1274 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 2777 2363 2835 2369
rect 2777 2360 2789 2363
rect 2556 2332 2789 2360
rect 2556 2320 2562 2332
rect 2777 2329 2789 2332
rect 2823 2329 2835 2363
rect 2777 2323 2835 2329
rect 3068 2292 3096 2391
rect 3786 2320 3792 2372
rect 3844 2360 3850 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3844 2332 4169 2360
rect 3844 2320 3850 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4356 2360 4384 2468
rect 4448 2437 4476 2604
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 10134 2564 10140 2576
rect 5644 2536 10140 2564
rect 5644 2437 5672 2536
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 14366 2496 14372 2508
rect 7668 2468 14372 2496
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2397 4491 2431
rect 5629 2431 5687 2437
rect 4433 2391 4491 2397
rect 5000 2400 5488 2428
rect 5000 2360 5028 2400
rect 4356 2332 5028 2360
rect 4157 2323 4215 2329
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5132 2332 5365 2360
rect 5132 2320 5138 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5460 2360 5488 2400
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6420 2400 6561 2428
rect 6420 2388 6426 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7558 2360 7564 2372
rect 5460 2332 7564 2360
rect 5353 2323 5411 2329
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 7668 2292 7696 2468
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 18230 2456 18236 2508
rect 18288 2456 18294 2508
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7800 2400 7845 2428
rect 7800 2388 7806 2400
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8996 2400 9137 2428
rect 8996 2388 9002 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10284 2400 10333 2428
rect 10284 2388 10290 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11572 2400 11713 2428
rect 11572 2388 11578 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12860 2400 12909 2428
rect 12860 2388 12866 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 15470 2428 15476 2440
rect 15431 2400 15476 2428
rect 14277 2391 14335 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 18248 2428 18276 2456
rect 18095 2400 18276 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 19058 2388 19064 2440
rect 19116 2428 19122 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19116 2400 19441 2428
rect 19116 2388 19122 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 20806 2428 20812 2440
rect 20671 2400 20812 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21140 2400 22017 2428
rect 21140 2388 21146 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 23382 2428 23388 2440
rect 23247 2400 23388 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 23382 2388 23388 2400
rect 23440 2388 23446 2440
rect 25038 2428 25044 2440
rect 24999 2400 25044 2428
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 27614 2428 27620 2440
rect 26292 2400 26337 2428
rect 27575 2400 27620 2428
rect 26292 2388 26298 2400
rect 27614 2388 27620 2400
rect 27672 2388 27678 2440
rect 28350 2428 28356 2440
rect 28311 2400 28356 2428
rect 28350 2388 28356 2400
rect 28408 2388 28414 2440
rect 29546 2388 29552 2440
rect 29604 2428 29610 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29604 2400 29745 2428
rect 29604 2388 29610 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30892 2400 30941 2428
rect 30892 2388 30898 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 32122 2388 32128 2440
rect 32180 2428 32186 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32180 2400 32321 2428
rect 32180 2388 32186 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33505 2431 33563 2437
rect 33505 2428 33517 2431
rect 33468 2400 33517 2428
rect 33468 2388 33474 2400
rect 33505 2397 33517 2400
rect 33551 2397 33563 2431
rect 33505 2391 33563 2397
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14148 2332 14565 2360
rect 14148 2320 14154 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 15378 2320 15384 2372
rect 15436 2360 15442 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15436 2332 15761 2360
rect 15436 2320 15442 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15749 2323 15807 2329
rect 16666 2320 16672 2372
rect 16724 2360 16730 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 16724 2332 17141 2360
rect 16724 2320 16730 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 17129 2323 17187 2329
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 18288 2332 18337 2360
rect 18288 2320 18294 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 18325 2323 18383 2329
rect 19242 2320 19248 2372
rect 19300 2360 19306 2372
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 19300 2332 19717 2360
rect 19300 2320 19306 2332
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 20530 2320 20536 2372
rect 20588 2360 20594 2372
rect 20901 2363 20959 2369
rect 20901 2360 20913 2363
rect 20588 2332 20913 2360
rect 20588 2320 20594 2332
rect 20901 2329 20913 2332
rect 20947 2329 20959 2363
rect 20901 2323 20959 2329
rect 21818 2320 21824 2372
rect 21876 2360 21882 2372
rect 22281 2363 22339 2369
rect 22281 2360 22293 2363
rect 21876 2332 22293 2360
rect 21876 2320 21882 2332
rect 22281 2329 22293 2332
rect 22327 2329 22339 2363
rect 22281 2323 22339 2329
rect 23106 2320 23112 2372
rect 23164 2360 23170 2372
rect 23477 2363 23535 2369
rect 23477 2360 23489 2363
rect 23164 2332 23489 2360
rect 23164 2320 23170 2332
rect 23477 2329 23489 2332
rect 23523 2329 23535 2363
rect 23477 2323 23535 2329
rect 24394 2320 24400 2372
rect 24452 2360 24458 2372
rect 24765 2363 24823 2369
rect 24765 2360 24777 2363
rect 24452 2332 24777 2360
rect 24452 2320 24458 2332
rect 24765 2329 24777 2332
rect 24811 2329 24823 2363
rect 24765 2323 24823 2329
rect 25682 2320 25688 2372
rect 25740 2360 25746 2372
rect 25961 2363 26019 2369
rect 25961 2360 25973 2363
rect 25740 2332 25973 2360
rect 25740 2320 25746 2332
rect 25961 2329 25973 2332
rect 26007 2329 26019 2363
rect 25961 2323 26019 2329
rect 26970 2320 26976 2372
rect 27028 2360 27034 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 27028 2332 27353 2360
rect 27028 2320 27034 2332
rect 27341 2329 27353 2332
rect 27387 2329 27399 2363
rect 27341 2323 27399 2329
rect 28258 2320 28264 2372
rect 28316 2360 28322 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28316 2332 28641 2360
rect 28316 2320 28322 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 3068 2264 7696 2292
rect 34333 2295 34391 2301
rect 34333 2261 34345 2295
rect 34379 2292 34391 2295
rect 34606 2292 34612 2304
rect 34379 2264 34612 2292
rect 34379 2261 34391 2264
rect 34333 2255 34391 2261
rect 34606 2252 34612 2264
rect 34664 2252 34670 2304
rect 1104 2202 35027 2224
rect 1104 2150 9390 2202
rect 9442 2150 9454 2202
rect 9506 2150 9518 2202
rect 9570 2150 9582 2202
rect 9634 2150 9646 2202
rect 9698 2150 17831 2202
rect 17883 2150 17895 2202
rect 17947 2150 17959 2202
rect 18011 2150 18023 2202
rect 18075 2150 18087 2202
rect 18139 2150 26272 2202
rect 26324 2150 26336 2202
rect 26388 2150 26400 2202
rect 26452 2150 26464 2202
rect 26516 2150 26528 2202
rect 26580 2150 34713 2202
rect 34765 2150 34777 2202
rect 34829 2150 34841 2202
rect 34893 2150 34905 2202
rect 34957 2150 34969 2202
rect 35021 2150 35027 2202
rect 1104 2128 35027 2150
<< via1 >>
rect 9390 33702 9442 33754
rect 9454 33702 9506 33754
rect 9518 33702 9570 33754
rect 9582 33702 9634 33754
rect 9646 33702 9698 33754
rect 17831 33702 17883 33754
rect 17895 33702 17947 33754
rect 17959 33702 18011 33754
rect 18023 33702 18075 33754
rect 18087 33702 18139 33754
rect 26272 33702 26324 33754
rect 26336 33702 26388 33754
rect 26400 33702 26452 33754
rect 26464 33702 26516 33754
rect 26528 33702 26580 33754
rect 34713 33702 34765 33754
rect 34777 33702 34829 33754
rect 34841 33702 34893 33754
rect 34905 33702 34957 33754
rect 34969 33702 35021 33754
rect 4896 33575 4948 33584
rect 4896 33541 4905 33575
rect 4905 33541 4939 33575
rect 4939 33541 4948 33575
rect 4896 33532 4948 33541
rect 7840 33575 7892 33584
rect 7840 33541 7849 33575
rect 7849 33541 7883 33575
rect 7883 33541 7892 33575
rect 7840 33532 7892 33541
rect 10600 33532 10652 33584
rect 13820 33532 13872 33584
rect 16580 33532 16632 33584
rect 19432 33532 19484 33584
rect 22652 33575 22704 33584
rect 22652 33541 22661 33575
rect 22661 33541 22695 33575
rect 22695 33541 22704 33575
rect 22652 33532 22704 33541
rect 25596 33575 25648 33584
rect 25596 33541 25605 33575
rect 25605 33541 25639 33575
rect 25639 33541 25648 33575
rect 25596 33532 25648 33541
rect 28540 33575 28592 33584
rect 28540 33541 28549 33575
rect 28549 33541 28583 33575
rect 28583 33541 28592 33575
rect 28540 33532 28592 33541
rect 31484 33575 31536 33584
rect 31484 33541 31493 33575
rect 31493 33541 31527 33575
rect 31527 33541 31536 33575
rect 31484 33532 31536 33541
rect 34244 33575 34296 33584
rect 34244 33541 34253 33575
rect 34253 33541 34287 33575
rect 34287 33541 34296 33575
rect 34244 33532 34296 33541
rect 8024 33371 8076 33380
rect 8024 33337 8033 33371
rect 8033 33337 8067 33371
rect 8067 33337 8076 33371
rect 8024 33328 8076 33337
rect 12256 33328 12308 33380
rect 14280 33371 14332 33380
rect 14280 33337 14289 33371
rect 14289 33337 14323 33371
rect 14323 33337 14332 33371
rect 14280 33328 14332 33337
rect 16856 33371 16908 33380
rect 16856 33337 16865 33371
rect 16865 33337 16899 33371
rect 16899 33337 16908 33371
rect 16856 33328 16908 33337
rect 19524 33371 19576 33380
rect 19524 33337 19533 33371
rect 19533 33337 19567 33371
rect 19567 33337 19576 33371
rect 19524 33328 19576 33337
rect 20260 33328 20312 33380
rect 25412 33371 25464 33380
rect 25412 33337 25421 33371
rect 25421 33337 25455 33371
rect 25455 33337 25464 33371
rect 25412 33328 25464 33337
rect 31300 33371 31352 33380
rect 31300 33337 31309 33371
rect 31309 33337 31343 33371
rect 31343 33337 31352 33371
rect 31300 33328 31352 33337
rect 33324 33328 33376 33380
rect 4988 33303 5040 33312
rect 4988 33269 4997 33303
rect 4997 33269 5031 33303
rect 5031 33269 5040 33303
rect 4988 33260 5040 33269
rect 20444 33260 20496 33312
rect 5170 33158 5222 33210
rect 5234 33158 5286 33210
rect 5298 33158 5350 33210
rect 5362 33158 5414 33210
rect 5426 33158 5478 33210
rect 13611 33158 13663 33210
rect 13675 33158 13727 33210
rect 13739 33158 13791 33210
rect 13803 33158 13855 33210
rect 13867 33158 13919 33210
rect 22052 33158 22104 33210
rect 22116 33158 22168 33210
rect 22180 33158 22232 33210
rect 22244 33158 22296 33210
rect 22308 33158 22360 33210
rect 30493 33158 30545 33210
rect 30557 33158 30609 33210
rect 30621 33158 30673 33210
rect 30685 33158 30737 33210
rect 30749 33158 30801 33210
rect 12072 33056 12124 33108
rect 20260 32988 20312 33040
rect 20444 32920 20496 32972
rect 20628 32963 20680 32972
rect 20628 32929 20637 32963
rect 20637 32929 20671 32963
rect 20671 32929 20680 32963
rect 20628 32920 20680 32929
rect 10508 32852 10560 32904
rect 16212 32784 16264 32836
rect 16856 32852 16908 32904
rect 19340 32852 19392 32904
rect 24584 32920 24636 32972
rect 22836 32852 22888 32904
rect 16764 32784 16816 32836
rect 10140 32759 10192 32768
rect 10140 32725 10149 32759
rect 10149 32725 10183 32759
rect 10183 32725 10192 32759
rect 10140 32716 10192 32725
rect 13268 32716 13320 32768
rect 25412 32784 25464 32836
rect 21272 32716 21324 32768
rect 22008 32716 22060 32768
rect 9390 32614 9442 32666
rect 9454 32614 9506 32666
rect 9518 32614 9570 32666
rect 9582 32614 9634 32666
rect 9646 32614 9698 32666
rect 17831 32614 17883 32666
rect 17895 32614 17947 32666
rect 17959 32614 18011 32666
rect 18023 32614 18075 32666
rect 18087 32614 18139 32666
rect 26272 32614 26324 32666
rect 26336 32614 26388 32666
rect 26400 32614 26452 32666
rect 26464 32614 26516 32666
rect 26528 32614 26580 32666
rect 34713 32614 34765 32666
rect 34777 32614 34829 32666
rect 34841 32614 34893 32666
rect 34905 32614 34957 32666
rect 34969 32614 35021 32666
rect 12256 32555 12308 32564
rect 12256 32521 12265 32555
rect 12265 32521 12299 32555
rect 12299 32521 12308 32555
rect 12256 32512 12308 32521
rect 14280 32512 14332 32564
rect 12072 32487 12124 32496
rect 12072 32453 12081 32487
rect 12081 32453 12115 32487
rect 12115 32453 12124 32487
rect 12072 32444 12124 32453
rect 13268 32487 13320 32496
rect 13268 32453 13277 32487
rect 13277 32453 13311 32487
rect 13311 32453 13320 32487
rect 13268 32444 13320 32453
rect 10324 32376 10376 32428
rect 10508 32419 10560 32428
rect 10508 32385 10517 32419
rect 10517 32385 10551 32419
rect 10551 32385 10560 32419
rect 10508 32376 10560 32385
rect 11428 32376 11480 32428
rect 19524 32444 19576 32496
rect 17868 32376 17920 32428
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 22468 32376 22520 32428
rect 23204 32419 23256 32428
rect 12348 32351 12400 32360
rect 8576 32240 8628 32292
rect 12348 32317 12357 32351
rect 12357 32317 12391 32351
rect 12391 32317 12400 32351
rect 12348 32308 12400 32317
rect 16764 32308 16816 32360
rect 17408 32351 17460 32360
rect 17408 32317 17417 32351
rect 17417 32317 17451 32351
rect 17451 32317 17460 32351
rect 17408 32308 17460 32317
rect 21272 32351 21324 32360
rect 21272 32317 21281 32351
rect 21281 32317 21315 32351
rect 21315 32317 21324 32351
rect 21272 32308 21324 32317
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 24492 32419 24544 32428
rect 24492 32385 24501 32419
rect 24501 32385 24535 32419
rect 24535 32385 24544 32419
rect 24492 32376 24544 32385
rect 24584 32376 24636 32428
rect 27712 32419 27764 32428
rect 27712 32385 27721 32419
rect 27721 32385 27755 32419
rect 27755 32385 27764 32419
rect 27712 32376 27764 32385
rect 28080 32419 28132 32428
rect 28080 32385 28089 32419
rect 28089 32385 28123 32419
rect 28123 32385 28132 32419
rect 28080 32376 28132 32385
rect 31300 32376 31352 32428
rect 33324 32419 33376 32428
rect 33324 32385 33333 32419
rect 33333 32385 33367 32419
rect 33367 32385 33376 32419
rect 33324 32376 33376 32385
rect 23388 32308 23440 32360
rect 21088 32240 21140 32292
rect 10048 32172 10100 32224
rect 10600 32215 10652 32224
rect 10600 32181 10609 32215
rect 10609 32181 10643 32215
rect 10643 32181 10652 32215
rect 10600 32172 10652 32181
rect 11888 32172 11940 32224
rect 13176 32172 13228 32224
rect 22836 32172 22888 32224
rect 25044 32172 25096 32224
rect 30196 32172 30248 32224
rect 33140 32215 33192 32224
rect 33140 32181 33149 32215
rect 33149 32181 33183 32215
rect 33183 32181 33192 32215
rect 33140 32172 33192 32181
rect 5170 32070 5222 32122
rect 5234 32070 5286 32122
rect 5298 32070 5350 32122
rect 5362 32070 5414 32122
rect 5426 32070 5478 32122
rect 13611 32070 13663 32122
rect 13675 32070 13727 32122
rect 13739 32070 13791 32122
rect 13803 32070 13855 32122
rect 13867 32070 13919 32122
rect 22052 32070 22104 32122
rect 22116 32070 22168 32122
rect 22180 32070 22232 32122
rect 22244 32070 22296 32122
rect 22308 32070 22360 32122
rect 30493 32070 30545 32122
rect 30557 32070 30609 32122
rect 30621 32070 30673 32122
rect 30685 32070 30737 32122
rect 30749 32070 30801 32122
rect 16120 31968 16172 32020
rect 18236 31968 18288 32020
rect 20628 31968 20680 32020
rect 23204 31968 23256 32020
rect 8760 31900 8812 31952
rect 11704 31900 11756 31952
rect 16856 31900 16908 31952
rect 9864 31875 9916 31884
rect 9864 31841 9873 31875
rect 9873 31841 9907 31875
rect 9907 31841 9916 31875
rect 9864 31832 9916 31841
rect 10508 31832 10560 31884
rect 17132 31875 17184 31884
rect 17132 31841 17141 31875
rect 17141 31841 17175 31875
rect 17175 31841 17184 31875
rect 17132 31832 17184 31841
rect 20536 31900 20588 31952
rect 8576 31807 8628 31816
rect 8576 31773 8585 31807
rect 8585 31773 8619 31807
rect 8619 31773 8628 31807
rect 8576 31764 8628 31773
rect 10140 31764 10192 31816
rect 11428 31807 11480 31816
rect 11428 31773 11437 31807
rect 11437 31773 11471 31807
rect 11471 31773 11480 31807
rect 11428 31764 11480 31773
rect 12348 31764 12400 31816
rect 14004 31764 14056 31816
rect 14280 31807 14332 31816
rect 14280 31773 14289 31807
rect 14289 31773 14323 31807
rect 14323 31773 14332 31807
rect 14280 31764 14332 31773
rect 14648 31764 14700 31816
rect 16120 31764 16172 31816
rect 10048 31696 10100 31748
rect 15568 31739 15620 31748
rect 15568 31705 15577 31739
rect 15577 31705 15611 31739
rect 15611 31705 15620 31739
rect 15568 31696 15620 31705
rect 17316 31807 17368 31816
rect 17316 31773 17325 31807
rect 17325 31773 17359 31807
rect 17359 31773 17368 31807
rect 17316 31764 17368 31773
rect 17868 31764 17920 31816
rect 21088 31832 21140 31884
rect 22468 31900 22520 31952
rect 8024 31628 8076 31680
rect 15752 31671 15804 31680
rect 15752 31637 15777 31671
rect 15777 31637 15804 31671
rect 20812 31764 20864 31816
rect 21180 31764 21232 31816
rect 21364 31764 21416 31816
rect 25044 31875 25096 31884
rect 25044 31841 25053 31875
rect 25053 31841 25087 31875
rect 25087 31841 25096 31875
rect 25044 31832 25096 31841
rect 25136 31875 25188 31884
rect 25136 31841 25145 31875
rect 25145 31841 25179 31875
rect 25179 31841 25188 31875
rect 25136 31832 25188 31841
rect 22836 31807 22888 31816
rect 21088 31739 21140 31748
rect 21088 31705 21097 31739
rect 21097 31705 21131 31739
rect 21131 31705 21140 31739
rect 21088 31696 21140 31705
rect 22836 31773 22845 31807
rect 22845 31773 22879 31807
rect 22879 31773 22888 31807
rect 22836 31764 22888 31773
rect 23664 31807 23716 31816
rect 23664 31773 23673 31807
rect 23673 31773 23707 31807
rect 23707 31773 23716 31807
rect 23664 31764 23716 31773
rect 26608 31807 26660 31816
rect 23388 31696 23440 31748
rect 26608 31773 26617 31807
rect 26617 31773 26651 31807
rect 26651 31773 26660 31807
rect 26608 31764 26660 31773
rect 26700 31696 26752 31748
rect 27712 31696 27764 31748
rect 15752 31628 15804 31637
rect 22744 31628 22796 31680
rect 23480 31671 23532 31680
rect 23480 31637 23489 31671
rect 23489 31637 23523 31671
rect 23523 31637 23532 31671
rect 23480 31628 23532 31637
rect 24768 31628 24820 31680
rect 9390 31526 9442 31578
rect 9454 31526 9506 31578
rect 9518 31526 9570 31578
rect 9582 31526 9634 31578
rect 9646 31526 9698 31578
rect 17831 31526 17883 31578
rect 17895 31526 17947 31578
rect 17959 31526 18011 31578
rect 18023 31526 18075 31578
rect 18087 31526 18139 31578
rect 26272 31526 26324 31578
rect 26336 31526 26388 31578
rect 26400 31526 26452 31578
rect 26464 31526 26516 31578
rect 26528 31526 26580 31578
rect 34713 31526 34765 31578
rect 34777 31526 34829 31578
rect 34841 31526 34893 31578
rect 34905 31526 34957 31578
rect 34969 31526 35021 31578
rect 9864 31424 9916 31476
rect 14280 31424 14332 31476
rect 16120 31467 16172 31476
rect 16120 31433 16129 31467
rect 16129 31433 16163 31467
rect 16163 31433 16172 31467
rect 16120 31424 16172 31433
rect 17316 31424 17368 31476
rect 20812 31467 20864 31476
rect 20812 31433 20846 31467
rect 20846 31433 20864 31467
rect 20812 31424 20864 31433
rect 25136 31424 25188 31476
rect 25228 31424 25280 31476
rect 25780 31424 25832 31476
rect 26608 31424 26660 31476
rect 9772 31356 9824 31408
rect 10048 31356 10100 31408
rect 10600 31356 10652 31408
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 9404 31220 9456 31272
rect 10048 31220 10100 31272
rect 12624 31288 12676 31340
rect 15568 31356 15620 31408
rect 19340 31356 19392 31408
rect 14096 31331 14148 31340
rect 14096 31297 14105 31331
rect 14105 31297 14139 31331
rect 14139 31297 14148 31331
rect 14096 31288 14148 31297
rect 14832 31331 14884 31340
rect 14832 31297 14841 31331
rect 14841 31297 14875 31331
rect 14875 31297 14884 31331
rect 14832 31288 14884 31297
rect 10600 31220 10652 31272
rect 13268 31263 13320 31272
rect 13268 31229 13277 31263
rect 13277 31229 13311 31263
rect 13311 31229 13320 31263
rect 13268 31220 13320 31229
rect 10692 31152 10744 31204
rect 10324 31084 10376 31136
rect 14280 31127 14332 31136
rect 14280 31093 14289 31127
rect 14289 31093 14323 31127
rect 14323 31093 14332 31127
rect 14280 31084 14332 31093
rect 14648 31220 14700 31272
rect 15476 31288 15528 31340
rect 16304 31331 16356 31340
rect 16304 31297 16313 31331
rect 16313 31297 16347 31331
rect 16347 31297 16356 31331
rect 16304 31288 16356 31297
rect 17132 31331 17184 31340
rect 17132 31297 17141 31331
rect 17141 31297 17175 31331
rect 17175 31297 17184 31331
rect 17132 31288 17184 31297
rect 15752 31220 15804 31272
rect 17684 31288 17736 31340
rect 20352 31288 20404 31340
rect 20996 31288 21048 31340
rect 22652 31331 22704 31340
rect 22652 31297 22661 31331
rect 22661 31297 22695 31331
rect 22695 31297 22704 31331
rect 22652 31288 22704 31297
rect 22744 31331 22796 31340
rect 22744 31297 22753 31331
rect 22753 31297 22787 31331
rect 22787 31297 22796 31331
rect 23020 31331 23072 31340
rect 22744 31288 22796 31297
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 23480 31331 23532 31340
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 21364 31220 21416 31272
rect 21456 31220 21508 31272
rect 23480 31297 23489 31331
rect 23489 31297 23523 31331
rect 23523 31297 23532 31331
rect 23480 31288 23532 31297
rect 24492 31288 24544 31340
rect 25228 31331 25280 31340
rect 23664 31220 23716 31272
rect 25228 31297 25237 31331
rect 25237 31297 25271 31331
rect 25271 31297 25280 31331
rect 25228 31288 25280 31297
rect 25320 31288 25372 31340
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 25044 31220 25096 31272
rect 26700 31288 26752 31340
rect 25780 31220 25832 31272
rect 29092 31263 29144 31272
rect 29092 31229 29101 31263
rect 29101 31229 29135 31263
rect 29135 31229 29144 31263
rect 29092 31220 29144 31229
rect 17040 31084 17092 31136
rect 21916 31084 21968 31136
rect 26056 31084 26108 31136
rect 28540 31084 28592 31136
rect 5170 30982 5222 31034
rect 5234 30982 5286 31034
rect 5298 30982 5350 31034
rect 5362 30982 5414 31034
rect 5426 30982 5478 31034
rect 13611 30982 13663 31034
rect 13675 30982 13727 31034
rect 13739 30982 13791 31034
rect 13803 30982 13855 31034
rect 13867 30982 13919 31034
rect 22052 30982 22104 31034
rect 22116 30982 22168 31034
rect 22180 30982 22232 31034
rect 22244 30982 22296 31034
rect 22308 30982 22360 31034
rect 30493 30982 30545 31034
rect 30557 30982 30609 31034
rect 30621 30982 30673 31034
rect 30685 30982 30737 31034
rect 30749 30982 30801 31034
rect 9404 30923 9456 30932
rect 9404 30889 9413 30923
rect 9413 30889 9447 30923
rect 9447 30889 9456 30923
rect 9404 30880 9456 30889
rect 10048 30923 10100 30932
rect 10048 30889 10057 30923
rect 10057 30889 10091 30923
rect 10091 30889 10100 30923
rect 10048 30880 10100 30889
rect 10232 30880 10284 30932
rect 13268 30880 13320 30932
rect 17408 30880 17460 30932
rect 20996 30923 21048 30932
rect 20996 30889 21005 30923
rect 21005 30889 21039 30923
rect 21039 30889 21048 30923
rect 20996 30880 21048 30889
rect 23020 30880 23072 30932
rect 14832 30812 14884 30864
rect 10508 30744 10560 30796
rect 9956 30719 10008 30728
rect 9956 30685 9965 30719
rect 9965 30685 9999 30719
rect 9999 30685 10008 30719
rect 9956 30676 10008 30685
rect 10140 30719 10192 30728
rect 10140 30685 10149 30719
rect 10149 30685 10183 30719
rect 10183 30685 10192 30719
rect 10140 30676 10192 30685
rect 10324 30676 10376 30728
rect 15752 30787 15804 30796
rect 15752 30753 15761 30787
rect 15761 30753 15795 30787
rect 15795 30753 15804 30787
rect 15752 30744 15804 30753
rect 14096 30676 14148 30728
rect 14556 30719 14608 30728
rect 14556 30685 14565 30719
rect 14565 30685 14599 30719
rect 14599 30685 14608 30719
rect 14556 30676 14608 30685
rect 14924 30719 14976 30728
rect 14924 30685 14933 30719
rect 14933 30685 14967 30719
rect 14967 30685 14976 30719
rect 14924 30676 14976 30685
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 23388 30812 23440 30864
rect 16856 30719 16908 30728
rect 16856 30685 16865 30719
rect 16865 30685 16899 30719
rect 16899 30685 16908 30719
rect 16856 30676 16908 30685
rect 17040 30719 17092 30728
rect 17040 30685 17049 30719
rect 17049 30685 17083 30719
rect 17083 30685 17092 30719
rect 17040 30676 17092 30685
rect 10600 30540 10652 30592
rect 14004 30540 14056 30592
rect 16304 30608 16356 30660
rect 18788 30608 18840 30660
rect 21456 30676 21508 30728
rect 23664 30744 23716 30796
rect 25228 30744 25280 30796
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 25044 30719 25096 30728
rect 25044 30685 25053 30719
rect 25053 30685 25087 30719
rect 25087 30685 25096 30719
rect 25044 30676 25096 30685
rect 25596 30719 25648 30728
rect 25596 30685 25605 30719
rect 25605 30685 25639 30719
rect 25639 30685 25648 30719
rect 25596 30676 25648 30685
rect 26056 30719 26108 30728
rect 26056 30685 26065 30719
rect 26065 30685 26099 30719
rect 26099 30685 26108 30719
rect 26056 30676 26108 30685
rect 29092 30744 29144 30796
rect 28908 30719 28960 30728
rect 26976 30608 27028 30660
rect 27620 30608 27672 30660
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 28724 30608 28776 30660
rect 9390 30438 9442 30490
rect 9454 30438 9506 30490
rect 9518 30438 9570 30490
rect 9582 30438 9634 30490
rect 9646 30438 9698 30490
rect 17831 30438 17883 30490
rect 17895 30438 17947 30490
rect 17959 30438 18011 30490
rect 18023 30438 18075 30490
rect 18087 30438 18139 30490
rect 26272 30438 26324 30490
rect 26336 30438 26388 30490
rect 26400 30438 26452 30490
rect 26464 30438 26516 30490
rect 26528 30438 26580 30490
rect 34713 30438 34765 30490
rect 34777 30438 34829 30490
rect 34841 30438 34893 30490
rect 34905 30438 34957 30490
rect 34969 30438 35021 30490
rect 18788 30268 18840 30320
rect 14280 30243 14332 30252
rect 14280 30209 14289 30243
rect 14289 30209 14323 30243
rect 14323 30209 14332 30243
rect 14280 30200 14332 30209
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 20168 30200 20220 30252
rect 20812 30200 20864 30252
rect 20904 30200 20956 30252
rect 24676 30243 24728 30252
rect 24676 30209 24685 30243
rect 24685 30209 24719 30243
rect 24719 30209 24728 30243
rect 24676 30200 24728 30209
rect 25136 30243 25188 30252
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 25228 30200 25280 30252
rect 26056 30336 26108 30388
rect 25688 30200 25740 30252
rect 25044 30132 25096 30184
rect 26976 30200 27028 30252
rect 27528 30200 27580 30252
rect 29092 30336 29144 30388
rect 28080 30311 28132 30320
rect 28080 30277 28089 30311
rect 28089 30277 28123 30311
rect 28123 30277 28132 30311
rect 28080 30268 28132 30277
rect 28540 30311 28592 30320
rect 28540 30277 28549 30311
rect 28549 30277 28583 30311
rect 28583 30277 28592 30311
rect 28540 30268 28592 30277
rect 28724 30243 28776 30252
rect 28724 30209 28733 30243
rect 28733 30209 28767 30243
rect 28767 30209 28776 30243
rect 28724 30200 28776 30209
rect 29000 30243 29052 30252
rect 29000 30209 29009 30243
rect 29009 30209 29043 30243
rect 29043 30209 29052 30243
rect 29000 30200 29052 30209
rect 29184 30243 29236 30252
rect 29184 30209 29193 30243
rect 29193 30209 29227 30243
rect 29227 30209 29236 30243
rect 29184 30200 29236 30209
rect 28632 30132 28684 30184
rect 28080 30064 28132 30116
rect 12900 29996 12952 30048
rect 20628 29996 20680 30048
rect 27436 29996 27488 30048
rect 28632 29996 28684 30048
rect 5170 29894 5222 29946
rect 5234 29894 5286 29946
rect 5298 29894 5350 29946
rect 5362 29894 5414 29946
rect 5426 29894 5478 29946
rect 13611 29894 13663 29946
rect 13675 29894 13727 29946
rect 13739 29894 13791 29946
rect 13803 29894 13855 29946
rect 13867 29894 13919 29946
rect 22052 29894 22104 29946
rect 22116 29894 22168 29946
rect 22180 29894 22232 29946
rect 22244 29894 22296 29946
rect 22308 29894 22360 29946
rect 30493 29894 30545 29946
rect 30557 29894 30609 29946
rect 30621 29894 30673 29946
rect 30685 29894 30737 29946
rect 30749 29894 30801 29946
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 25044 29835 25096 29844
rect 25044 29801 25053 29835
rect 25053 29801 25087 29835
rect 25087 29801 25096 29835
rect 25044 29792 25096 29801
rect 25136 29792 25188 29844
rect 9036 29724 9088 29776
rect 10692 29656 10744 29708
rect 10416 29631 10468 29640
rect 10416 29597 10425 29631
rect 10425 29597 10459 29631
rect 10459 29597 10468 29631
rect 10416 29588 10468 29597
rect 10140 29520 10192 29572
rect 12900 29588 12952 29640
rect 10692 29563 10744 29572
rect 10692 29529 10701 29563
rect 10701 29529 10735 29563
rect 10735 29529 10744 29563
rect 10692 29520 10744 29529
rect 15016 29588 15068 29640
rect 19248 29588 19300 29640
rect 20536 29656 20588 29708
rect 20812 29656 20864 29708
rect 23204 29724 23256 29776
rect 27160 29656 27212 29708
rect 20352 29588 20404 29640
rect 20720 29588 20772 29640
rect 24768 29631 24820 29640
rect 14280 29520 14332 29572
rect 15108 29563 15160 29572
rect 15108 29529 15117 29563
rect 15117 29529 15151 29563
rect 15151 29529 15160 29563
rect 15108 29520 15160 29529
rect 20904 29520 20956 29572
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 21640 29520 21692 29572
rect 24584 29520 24636 29572
rect 26976 29588 27028 29640
rect 27528 29631 27580 29640
rect 27528 29597 27537 29631
rect 27537 29597 27571 29631
rect 27571 29597 27580 29631
rect 27528 29588 27580 29597
rect 27620 29631 27672 29640
rect 27620 29597 27629 29631
rect 27629 29597 27663 29631
rect 27663 29597 27672 29631
rect 27620 29588 27672 29597
rect 28356 29631 28408 29640
rect 27712 29520 27764 29572
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 28908 29724 28960 29776
rect 29000 29656 29052 29708
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 29184 29588 29236 29640
rect 9312 29452 9364 29504
rect 9956 29452 10008 29504
rect 10416 29452 10468 29504
rect 12624 29452 12676 29504
rect 12808 29495 12860 29504
rect 12808 29461 12817 29495
rect 12817 29461 12851 29495
rect 12851 29461 12860 29495
rect 12808 29452 12860 29461
rect 19524 29495 19576 29504
rect 19524 29461 19533 29495
rect 19533 29461 19567 29495
rect 19567 29461 19576 29495
rect 19524 29452 19576 29461
rect 21456 29452 21508 29504
rect 9390 29350 9442 29402
rect 9454 29350 9506 29402
rect 9518 29350 9570 29402
rect 9582 29350 9634 29402
rect 9646 29350 9698 29402
rect 17831 29350 17883 29402
rect 17895 29350 17947 29402
rect 17959 29350 18011 29402
rect 18023 29350 18075 29402
rect 18087 29350 18139 29402
rect 26272 29350 26324 29402
rect 26336 29350 26388 29402
rect 26400 29350 26452 29402
rect 26464 29350 26516 29402
rect 26528 29350 26580 29402
rect 34713 29350 34765 29402
rect 34777 29350 34829 29402
rect 34841 29350 34893 29402
rect 34905 29350 34957 29402
rect 34969 29350 35021 29402
rect 12900 29248 12952 29300
rect 14556 29291 14608 29300
rect 14556 29257 14565 29291
rect 14565 29257 14599 29291
rect 14599 29257 14608 29291
rect 14556 29248 14608 29257
rect 14924 29248 14976 29300
rect 20168 29291 20220 29300
rect 9036 29155 9088 29164
rect 9036 29121 9045 29155
rect 9045 29121 9079 29155
rect 9079 29121 9088 29155
rect 9036 29112 9088 29121
rect 9312 29155 9364 29164
rect 9312 29121 9321 29155
rect 9321 29121 9355 29155
rect 9355 29121 9364 29155
rect 9312 29112 9364 29121
rect 9496 29155 9548 29164
rect 9496 29121 9505 29155
rect 9505 29121 9539 29155
rect 9539 29121 9548 29155
rect 9496 29112 9548 29121
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 15108 29180 15160 29232
rect 20168 29257 20177 29291
rect 20177 29257 20211 29291
rect 20211 29257 20220 29291
rect 20168 29248 20220 29257
rect 21364 29248 21416 29300
rect 27620 29248 27672 29300
rect 28356 29248 28408 29300
rect 29184 29248 29236 29300
rect 12624 29155 12676 29164
rect 12624 29121 12633 29155
rect 12633 29121 12667 29155
rect 12667 29121 12676 29155
rect 12624 29112 12676 29121
rect 12808 29112 12860 29164
rect 13452 29112 13504 29164
rect 15568 29155 15620 29164
rect 15568 29121 15577 29155
rect 15577 29121 15611 29155
rect 15611 29121 15620 29155
rect 15568 29112 15620 29121
rect 15752 29155 15804 29164
rect 15752 29121 15761 29155
rect 15761 29121 15795 29155
rect 15795 29121 15804 29155
rect 15752 29112 15804 29121
rect 19340 29112 19392 29164
rect 19524 29155 19576 29164
rect 19524 29121 19533 29155
rect 19533 29121 19567 29155
rect 19567 29121 19576 29155
rect 19524 29112 19576 29121
rect 20536 29180 20588 29232
rect 20444 29155 20496 29164
rect 20444 29121 20453 29155
rect 20453 29121 20487 29155
rect 20487 29121 20496 29155
rect 20628 29155 20680 29164
rect 20444 29112 20496 29121
rect 20628 29121 20637 29155
rect 20637 29121 20671 29155
rect 20671 29121 20680 29155
rect 20628 29112 20680 29121
rect 20720 29155 20772 29164
rect 20720 29121 20729 29155
rect 20729 29121 20763 29155
rect 20763 29121 20772 29155
rect 21640 29180 21692 29232
rect 25228 29223 25280 29232
rect 20720 29112 20772 29121
rect 15016 29044 15068 29096
rect 22376 29112 22428 29164
rect 25228 29189 25237 29223
rect 25237 29189 25271 29223
rect 25271 29189 25280 29223
rect 25228 29180 25280 29189
rect 22744 29155 22796 29164
rect 22744 29121 22753 29155
rect 22753 29121 22787 29155
rect 22787 29121 22796 29155
rect 22744 29112 22796 29121
rect 22836 29112 22888 29164
rect 23388 29112 23440 29164
rect 25780 29112 25832 29164
rect 27160 29155 27212 29164
rect 27160 29121 27169 29155
rect 27169 29121 27203 29155
rect 27203 29121 27212 29155
rect 27160 29112 27212 29121
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 28080 29155 28132 29164
rect 28080 29121 28089 29155
rect 28089 29121 28123 29155
rect 28123 29121 28132 29155
rect 28080 29112 28132 29121
rect 28172 29044 28224 29096
rect 28632 29044 28684 29096
rect 21272 29019 21324 29028
rect 21272 28985 21281 29019
rect 21281 28985 21315 29019
rect 21315 28985 21324 29019
rect 21272 28976 21324 28985
rect 8944 28908 8996 28960
rect 10600 28908 10652 28960
rect 20720 28908 20772 28960
rect 22468 29019 22520 29028
rect 22468 28985 22477 29019
rect 22477 28985 22511 29019
rect 22511 28985 22520 29019
rect 22468 28976 22520 28985
rect 27528 28976 27580 29028
rect 28908 28951 28960 28960
rect 28908 28917 28917 28951
rect 28917 28917 28951 28951
rect 28951 28917 28960 28951
rect 28908 28908 28960 28917
rect 5170 28806 5222 28858
rect 5234 28806 5286 28858
rect 5298 28806 5350 28858
rect 5362 28806 5414 28858
rect 5426 28806 5478 28858
rect 13611 28806 13663 28858
rect 13675 28806 13727 28858
rect 13739 28806 13791 28858
rect 13803 28806 13855 28858
rect 13867 28806 13919 28858
rect 22052 28806 22104 28858
rect 22116 28806 22168 28858
rect 22180 28806 22232 28858
rect 22244 28806 22296 28858
rect 22308 28806 22360 28858
rect 30493 28806 30545 28858
rect 30557 28806 30609 28858
rect 30621 28806 30673 28858
rect 30685 28806 30737 28858
rect 30749 28806 30801 28858
rect 21180 28747 21232 28756
rect 21180 28713 21189 28747
rect 21189 28713 21223 28747
rect 21223 28713 21232 28747
rect 21180 28704 21232 28713
rect 28908 28704 28960 28756
rect 13452 28636 13504 28688
rect 9496 28568 9548 28620
rect 11796 28568 11848 28620
rect 12532 28568 12584 28620
rect 15016 28568 15068 28620
rect 20720 28636 20772 28688
rect 20812 28568 20864 28620
rect 9036 28432 9088 28484
rect 10692 28500 10744 28552
rect 11336 28543 11388 28552
rect 11336 28509 11345 28543
rect 11345 28509 11379 28543
rect 11379 28509 11388 28543
rect 11336 28500 11388 28509
rect 12808 28500 12860 28552
rect 13084 28543 13136 28552
rect 13084 28509 13093 28543
rect 13093 28509 13127 28543
rect 13127 28509 13136 28543
rect 13084 28500 13136 28509
rect 13268 28543 13320 28552
rect 13268 28509 13277 28543
rect 13277 28509 13311 28543
rect 13311 28509 13320 28543
rect 14556 28543 14608 28552
rect 13268 28500 13320 28509
rect 14556 28509 14565 28543
rect 14565 28509 14599 28543
rect 14599 28509 14608 28543
rect 14556 28500 14608 28509
rect 15108 28500 15160 28552
rect 15384 28543 15436 28552
rect 15384 28509 15393 28543
rect 15393 28509 15427 28543
rect 15427 28509 15436 28543
rect 15384 28500 15436 28509
rect 15476 28500 15528 28552
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 19984 28543 20036 28552
rect 19984 28509 19993 28543
rect 19993 28509 20027 28543
rect 20027 28509 20036 28543
rect 19984 28500 20036 28509
rect 13452 28432 13504 28484
rect 15752 28432 15804 28484
rect 19248 28432 19300 28484
rect 20720 28543 20772 28552
rect 20720 28509 20751 28543
rect 20751 28509 20772 28543
rect 20720 28500 20772 28509
rect 20904 28543 20956 28552
rect 20904 28509 20913 28543
rect 20913 28509 20947 28543
rect 20947 28509 20956 28543
rect 20904 28500 20956 28509
rect 26700 28568 26752 28620
rect 27620 28568 27672 28620
rect 22836 28543 22888 28552
rect 22836 28509 22845 28543
rect 22845 28509 22879 28543
rect 22879 28509 22888 28543
rect 22836 28500 22888 28509
rect 23572 28500 23624 28552
rect 24676 28500 24728 28552
rect 27896 28500 27948 28552
rect 28724 28543 28776 28552
rect 28724 28509 28733 28543
rect 28733 28509 28767 28543
rect 28767 28509 28776 28543
rect 28724 28500 28776 28509
rect 9128 28407 9180 28416
rect 9128 28373 9137 28407
rect 9137 28373 9171 28407
rect 9171 28373 9180 28407
rect 9128 28364 9180 28373
rect 9312 28364 9364 28416
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 13084 28364 13136 28416
rect 15936 28364 15988 28416
rect 20536 28364 20588 28416
rect 22744 28364 22796 28416
rect 27252 28407 27304 28416
rect 27252 28373 27261 28407
rect 27261 28373 27295 28407
rect 27295 28373 27304 28407
rect 27252 28364 27304 28373
rect 9390 28262 9442 28314
rect 9454 28262 9506 28314
rect 9518 28262 9570 28314
rect 9582 28262 9634 28314
rect 9646 28262 9698 28314
rect 17831 28262 17883 28314
rect 17895 28262 17947 28314
rect 17959 28262 18011 28314
rect 18023 28262 18075 28314
rect 18087 28262 18139 28314
rect 26272 28262 26324 28314
rect 26336 28262 26388 28314
rect 26400 28262 26452 28314
rect 26464 28262 26516 28314
rect 26528 28262 26580 28314
rect 34713 28262 34765 28314
rect 34777 28262 34829 28314
rect 34841 28262 34893 28314
rect 34905 28262 34957 28314
rect 34969 28262 35021 28314
rect 8944 28160 8996 28212
rect 11336 28160 11388 28212
rect 9128 28024 9180 28076
rect 13084 28160 13136 28212
rect 15384 28203 15436 28212
rect 15384 28169 15393 28203
rect 15393 28169 15427 28203
rect 15427 28169 15436 28203
rect 15384 28160 15436 28169
rect 19800 28160 19852 28212
rect 12532 28067 12584 28076
rect 8760 27999 8812 28008
rect 8760 27965 8769 27999
rect 8769 27965 8803 27999
rect 8803 27965 8812 27999
rect 8760 27956 8812 27965
rect 8944 27999 8996 28008
rect 8944 27965 8953 27999
rect 8953 27965 8987 27999
rect 8987 27965 8996 27999
rect 12532 28033 12541 28067
rect 12541 28033 12575 28067
rect 12575 28033 12584 28067
rect 12532 28024 12584 28033
rect 13452 28092 13504 28144
rect 15016 28092 15068 28144
rect 15568 28092 15620 28144
rect 16028 28092 16080 28144
rect 19340 28092 19392 28144
rect 13268 28024 13320 28076
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 14280 28024 14332 28076
rect 15476 28024 15528 28076
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 20904 28092 20956 28144
rect 22376 28160 22428 28212
rect 22468 28160 22520 28212
rect 8944 27956 8996 27965
rect 9772 27956 9824 28008
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 14556 27956 14608 28008
rect 19984 27956 20036 28008
rect 22284 28024 22336 28076
rect 9128 27820 9180 27872
rect 9312 27820 9364 27872
rect 9588 27820 9640 27872
rect 9772 27863 9824 27872
rect 9772 27829 9781 27863
rect 9781 27829 9815 27863
rect 9815 27829 9824 27863
rect 9772 27820 9824 27829
rect 23572 28092 23624 28144
rect 22836 27956 22888 28008
rect 27344 28092 27396 28144
rect 31116 28092 31168 28144
rect 24860 28024 24912 28076
rect 25688 28067 25740 28076
rect 25688 28033 25697 28067
rect 25697 28033 25731 28067
rect 25731 28033 25740 28067
rect 25688 28024 25740 28033
rect 27068 28024 27120 28076
rect 27712 28024 27764 28076
rect 29000 28024 29052 28076
rect 32680 28024 32732 28076
rect 25136 27956 25188 28008
rect 25780 27999 25832 28008
rect 25780 27965 25789 27999
rect 25789 27965 25823 27999
rect 25823 27965 25832 27999
rect 25780 27956 25832 27965
rect 26240 27956 26292 28008
rect 25872 27888 25924 27940
rect 26608 27820 26660 27872
rect 30012 27820 30064 27872
rect 5170 27718 5222 27770
rect 5234 27718 5286 27770
rect 5298 27718 5350 27770
rect 5362 27718 5414 27770
rect 5426 27718 5478 27770
rect 13611 27718 13663 27770
rect 13675 27718 13727 27770
rect 13739 27718 13791 27770
rect 13803 27718 13855 27770
rect 13867 27718 13919 27770
rect 22052 27718 22104 27770
rect 22116 27718 22168 27770
rect 22180 27718 22232 27770
rect 22244 27718 22296 27770
rect 22308 27718 22360 27770
rect 30493 27718 30545 27770
rect 30557 27718 30609 27770
rect 30621 27718 30673 27770
rect 30685 27718 30737 27770
rect 30749 27718 30801 27770
rect 22376 27616 22428 27668
rect 24676 27616 24728 27668
rect 16028 27548 16080 27600
rect 24584 27548 24636 27600
rect 27896 27591 27948 27600
rect 27896 27557 27905 27591
rect 27905 27557 27939 27591
rect 27939 27557 27948 27591
rect 27896 27548 27948 27557
rect 9036 27480 9088 27532
rect 12532 27480 12584 27532
rect 9128 27412 9180 27464
rect 9588 27412 9640 27464
rect 14004 27480 14056 27532
rect 19892 27480 19944 27532
rect 13820 27412 13872 27464
rect 8208 27344 8260 27396
rect 12348 27344 12400 27396
rect 12624 27344 12676 27396
rect 13728 27344 13780 27396
rect 16028 27455 16080 27464
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 18236 27455 18288 27464
rect 16304 27344 16356 27396
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 21180 27412 21232 27464
rect 25872 27480 25924 27532
rect 25688 27455 25740 27464
rect 19524 27344 19576 27396
rect 20996 27344 21048 27396
rect 19800 27276 19852 27328
rect 21916 27276 21968 27328
rect 22376 27276 22428 27328
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 25596 27344 25648 27396
rect 26148 27412 26200 27464
rect 27712 27455 27764 27464
rect 26240 27344 26292 27396
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 28172 27412 28224 27464
rect 25780 27276 25832 27328
rect 26700 27276 26752 27328
rect 27068 27276 27120 27328
rect 29920 27412 29972 27464
rect 32220 27344 32272 27396
rect 28724 27276 28776 27328
rect 31208 27319 31260 27328
rect 31208 27285 31217 27319
rect 31217 27285 31251 27319
rect 31251 27285 31260 27319
rect 31208 27276 31260 27285
rect 9390 27174 9442 27226
rect 9454 27174 9506 27226
rect 9518 27174 9570 27226
rect 9582 27174 9634 27226
rect 9646 27174 9698 27226
rect 17831 27174 17883 27226
rect 17895 27174 17947 27226
rect 17959 27174 18011 27226
rect 18023 27174 18075 27226
rect 18087 27174 18139 27226
rect 26272 27174 26324 27226
rect 26336 27174 26388 27226
rect 26400 27174 26452 27226
rect 26464 27174 26516 27226
rect 26528 27174 26580 27226
rect 34713 27174 34765 27226
rect 34777 27174 34829 27226
rect 34841 27174 34893 27226
rect 34905 27174 34957 27226
rect 34969 27174 35021 27226
rect 12900 27072 12952 27124
rect 18236 27072 18288 27124
rect 9128 27004 9180 27056
rect 10324 27004 10376 27056
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 9772 26936 9824 26988
rect 12624 27004 12676 27056
rect 13820 27004 13872 27056
rect 14280 27004 14332 27056
rect 19800 27004 19852 27056
rect 25228 27072 25280 27124
rect 25504 27072 25556 27124
rect 31116 27115 31168 27124
rect 31116 27081 31125 27115
rect 31125 27081 31159 27115
rect 31159 27081 31168 27115
rect 31116 27072 31168 27081
rect 12440 26936 12492 26988
rect 13452 26936 13504 26988
rect 13728 26979 13780 26988
rect 13728 26945 13737 26979
rect 13737 26945 13771 26979
rect 13771 26945 13780 26979
rect 13728 26936 13780 26945
rect 9128 26911 9180 26920
rect 9128 26877 9137 26911
rect 9137 26877 9171 26911
rect 9171 26877 9180 26911
rect 9128 26868 9180 26877
rect 15752 26979 15804 26988
rect 15752 26945 15761 26979
rect 15761 26945 15795 26979
rect 15795 26945 15804 26979
rect 15752 26936 15804 26945
rect 16396 26936 16448 26988
rect 18328 26936 18380 26988
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 21180 26936 21232 26988
rect 24768 26936 24820 26988
rect 25136 26979 25188 26988
rect 25136 26945 25145 26979
rect 25145 26945 25179 26979
rect 25179 26945 25188 26979
rect 25136 26936 25188 26945
rect 25596 26979 25648 26988
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 26148 27004 26200 27056
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 27436 26979 27488 26988
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 30012 26979 30064 26988
rect 30012 26945 30021 26979
rect 30021 26945 30055 26979
rect 30055 26945 30064 26979
rect 30012 26936 30064 26945
rect 16672 26868 16724 26920
rect 26148 26868 26200 26920
rect 27620 26868 27672 26920
rect 29920 26868 29972 26920
rect 8760 26732 8812 26784
rect 9220 26732 9272 26784
rect 11152 26732 11204 26784
rect 12624 26732 12676 26784
rect 20536 26732 20588 26784
rect 20904 26732 20956 26784
rect 5170 26630 5222 26682
rect 5234 26630 5286 26682
rect 5298 26630 5350 26682
rect 5362 26630 5414 26682
rect 5426 26630 5478 26682
rect 13611 26630 13663 26682
rect 13675 26630 13727 26682
rect 13739 26630 13791 26682
rect 13803 26630 13855 26682
rect 13867 26630 13919 26682
rect 22052 26630 22104 26682
rect 22116 26630 22168 26682
rect 22180 26630 22232 26682
rect 22244 26630 22296 26682
rect 22308 26630 22360 26682
rect 30493 26630 30545 26682
rect 30557 26630 30609 26682
rect 30621 26630 30673 26682
rect 30685 26630 30737 26682
rect 30749 26630 30801 26682
rect 12440 26528 12492 26580
rect 12900 26528 12952 26580
rect 13360 26528 13412 26580
rect 16672 26571 16724 26580
rect 16672 26537 16681 26571
rect 16681 26537 16715 26571
rect 16715 26537 16724 26571
rect 16672 26528 16724 26537
rect 25136 26528 25188 26580
rect 27068 26571 27120 26580
rect 27068 26537 27077 26571
rect 27077 26537 27111 26571
rect 27111 26537 27120 26571
rect 27068 26528 27120 26537
rect 32220 26571 32272 26580
rect 32220 26537 32229 26571
rect 32229 26537 32263 26571
rect 32263 26537 32272 26571
rect 32220 26528 32272 26537
rect 9312 26460 9364 26512
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 11152 26392 11204 26401
rect 18972 26460 19024 26512
rect 12808 26392 12860 26444
rect 13452 26392 13504 26444
rect 12624 26367 12676 26376
rect 12624 26333 12633 26367
rect 12633 26333 12667 26367
rect 12667 26333 12676 26367
rect 12624 26324 12676 26333
rect 9036 26256 9088 26308
rect 12532 26256 12584 26308
rect 13452 26299 13504 26308
rect 13452 26265 13463 26299
rect 13463 26265 13504 26299
rect 18236 26392 18288 26444
rect 19340 26392 19392 26444
rect 21180 26460 21232 26512
rect 22744 26460 22796 26512
rect 25504 26435 25556 26444
rect 25504 26401 25513 26435
rect 25513 26401 25547 26435
rect 25547 26401 25556 26435
rect 25504 26392 25556 26401
rect 13452 26256 13504 26265
rect 16856 26256 16908 26308
rect 18236 26256 18288 26308
rect 24860 26324 24912 26376
rect 25320 26324 25372 26376
rect 25596 26367 25648 26376
rect 25596 26333 25605 26367
rect 25605 26333 25639 26367
rect 25639 26333 25648 26367
rect 25596 26324 25648 26333
rect 26516 26460 26568 26512
rect 26792 26460 26844 26512
rect 28632 26460 28684 26512
rect 22560 26299 22612 26308
rect 22560 26265 22569 26299
rect 22569 26265 22603 26299
rect 22603 26265 22612 26299
rect 22560 26256 22612 26265
rect 24584 26256 24636 26308
rect 26516 26367 26568 26376
rect 9312 26188 9364 26240
rect 19892 26188 19944 26240
rect 21180 26188 21232 26240
rect 26516 26333 26525 26367
rect 26525 26333 26559 26367
rect 26559 26333 26568 26367
rect 26516 26324 26568 26333
rect 26608 26367 26660 26376
rect 26608 26333 26617 26367
rect 26617 26333 26651 26367
rect 26651 26333 26660 26367
rect 26608 26324 26660 26333
rect 27160 26324 27212 26376
rect 32404 26367 32456 26376
rect 32404 26333 32413 26367
rect 32413 26333 32447 26367
rect 32447 26333 32456 26367
rect 32404 26324 32456 26333
rect 32680 26367 32732 26376
rect 32680 26333 32689 26367
rect 32689 26333 32723 26367
rect 32723 26333 32732 26367
rect 32680 26324 32732 26333
rect 26608 26188 26660 26240
rect 29092 26256 29144 26308
rect 31208 26256 31260 26308
rect 27528 26188 27580 26240
rect 9390 26086 9442 26138
rect 9454 26086 9506 26138
rect 9518 26086 9570 26138
rect 9582 26086 9634 26138
rect 9646 26086 9698 26138
rect 17831 26086 17883 26138
rect 17895 26086 17947 26138
rect 17959 26086 18011 26138
rect 18023 26086 18075 26138
rect 18087 26086 18139 26138
rect 26272 26086 26324 26138
rect 26336 26086 26388 26138
rect 26400 26086 26452 26138
rect 26464 26086 26516 26138
rect 26528 26086 26580 26138
rect 34713 26086 34765 26138
rect 34777 26086 34829 26138
rect 34841 26086 34893 26138
rect 34905 26086 34957 26138
rect 34969 26086 35021 26138
rect 12532 25984 12584 26036
rect 9312 25848 9364 25900
rect 12348 25959 12400 25968
rect 12348 25925 12357 25959
rect 12357 25925 12391 25959
rect 12391 25925 12400 25959
rect 12348 25916 12400 25925
rect 12440 25959 12492 25968
rect 12440 25925 12449 25959
rect 12449 25925 12483 25959
rect 12483 25925 12492 25959
rect 12440 25916 12492 25925
rect 9220 25780 9272 25832
rect 9588 25823 9640 25832
rect 9588 25789 9597 25823
rect 9597 25789 9631 25823
rect 9631 25789 9640 25823
rect 9588 25780 9640 25789
rect 12256 25848 12308 25900
rect 14740 25984 14792 26036
rect 16856 26027 16908 26036
rect 16856 25993 16865 26027
rect 16865 25993 16899 26027
rect 16899 25993 16908 26027
rect 16856 25984 16908 25993
rect 13360 25959 13412 25968
rect 13360 25925 13369 25959
rect 13369 25925 13403 25959
rect 13403 25925 13412 25959
rect 13360 25916 13412 25925
rect 16672 25916 16724 25968
rect 21916 25916 21968 25968
rect 9864 25780 9916 25832
rect 13452 25891 13504 25900
rect 13452 25857 13466 25891
rect 13466 25857 13500 25891
rect 13500 25857 13504 25891
rect 17040 25891 17092 25900
rect 13452 25848 13504 25857
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 19616 25891 19668 25900
rect 16304 25780 16356 25832
rect 16488 25780 16540 25832
rect 19616 25857 19625 25891
rect 19625 25857 19659 25891
rect 19659 25857 19668 25891
rect 19616 25848 19668 25857
rect 14464 25712 14516 25764
rect 21180 25848 21232 25900
rect 22376 25848 22428 25900
rect 25044 25984 25096 26036
rect 25688 25984 25740 26036
rect 27252 25984 27304 26036
rect 29920 26027 29972 26036
rect 29920 25993 29929 26027
rect 29929 25993 29963 26027
rect 29963 25993 29972 26027
rect 29920 25984 29972 25993
rect 25504 25916 25556 25968
rect 28632 25959 28684 25968
rect 28632 25925 28641 25959
rect 28641 25925 28675 25959
rect 28675 25925 28684 25959
rect 28632 25916 28684 25925
rect 31484 25916 31536 25968
rect 24676 25891 24728 25900
rect 24676 25857 24685 25891
rect 24685 25857 24719 25891
rect 24719 25857 24728 25891
rect 24676 25848 24728 25857
rect 26516 25891 26568 25900
rect 26516 25857 26525 25891
rect 26525 25857 26559 25891
rect 26559 25857 26568 25891
rect 26516 25848 26568 25857
rect 27620 25891 27672 25900
rect 27620 25857 27629 25891
rect 27629 25857 27663 25891
rect 27663 25857 27672 25891
rect 27620 25848 27672 25857
rect 31944 25848 31996 25900
rect 32772 25891 32824 25900
rect 32772 25857 32781 25891
rect 32781 25857 32815 25891
rect 32815 25857 32824 25891
rect 32772 25848 32824 25857
rect 23388 25780 23440 25832
rect 26700 25780 26752 25832
rect 27068 25780 27120 25832
rect 25044 25712 25096 25764
rect 27160 25712 27212 25764
rect 27528 25823 27580 25832
rect 27528 25789 27537 25823
rect 27537 25789 27571 25823
rect 27571 25789 27580 25823
rect 27528 25780 27580 25789
rect 12716 25644 12768 25696
rect 13084 25687 13136 25696
rect 13084 25653 13093 25687
rect 13093 25653 13127 25687
rect 13127 25653 13136 25687
rect 13084 25644 13136 25653
rect 18328 25687 18380 25696
rect 18328 25653 18337 25687
rect 18337 25653 18371 25687
rect 18371 25653 18380 25687
rect 18328 25644 18380 25653
rect 32312 25687 32364 25696
rect 32312 25653 32321 25687
rect 32321 25653 32355 25687
rect 32355 25653 32364 25687
rect 32312 25644 32364 25653
rect 5170 25542 5222 25594
rect 5234 25542 5286 25594
rect 5298 25542 5350 25594
rect 5362 25542 5414 25594
rect 5426 25542 5478 25594
rect 13611 25542 13663 25594
rect 13675 25542 13727 25594
rect 13739 25542 13791 25594
rect 13803 25542 13855 25594
rect 13867 25542 13919 25594
rect 22052 25542 22104 25594
rect 22116 25542 22168 25594
rect 22180 25542 22232 25594
rect 22244 25542 22296 25594
rect 22308 25542 22360 25594
rect 30493 25542 30545 25594
rect 30557 25542 30609 25594
rect 30621 25542 30673 25594
rect 30685 25542 30737 25594
rect 30749 25542 30801 25594
rect 16304 25415 16356 25424
rect 16304 25381 16313 25415
rect 16313 25381 16347 25415
rect 16347 25381 16356 25415
rect 16304 25372 16356 25381
rect 3332 25236 3384 25288
rect 4068 25279 4120 25288
rect 4068 25245 4077 25279
rect 4077 25245 4111 25279
rect 4111 25245 4120 25279
rect 4068 25236 4120 25245
rect 4252 25279 4304 25288
rect 4252 25245 4261 25279
rect 4261 25245 4295 25279
rect 4295 25245 4304 25279
rect 4252 25236 4304 25245
rect 6828 25236 6880 25288
rect 7840 25236 7892 25288
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 13084 25304 13136 25356
rect 12716 25279 12768 25288
rect 12716 25245 12725 25279
rect 12725 25245 12759 25279
rect 12759 25245 12768 25279
rect 12716 25236 12768 25245
rect 4160 25168 4212 25220
rect 15660 25236 15712 25288
rect 15936 25236 15988 25288
rect 16672 25440 16724 25492
rect 19800 25483 19852 25492
rect 19800 25449 19809 25483
rect 19809 25449 19843 25483
rect 19843 25449 19852 25483
rect 19800 25440 19852 25449
rect 25596 25440 25648 25492
rect 26792 25440 26844 25492
rect 27620 25440 27672 25492
rect 21180 25347 21232 25356
rect 21180 25313 21189 25347
rect 21189 25313 21223 25347
rect 21223 25313 21232 25347
rect 21180 25304 21232 25313
rect 26608 25347 26660 25356
rect 26608 25313 26617 25347
rect 26617 25313 26651 25347
rect 26651 25313 26660 25347
rect 26608 25304 26660 25313
rect 20904 25279 20956 25288
rect 20904 25245 20922 25279
rect 20922 25245 20956 25279
rect 20904 25236 20956 25245
rect 23480 25236 23532 25288
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 24676 25236 24728 25288
rect 27344 25279 27396 25288
rect 27344 25245 27352 25279
rect 27352 25245 27386 25279
rect 27386 25245 27396 25279
rect 27344 25236 27396 25245
rect 30104 25279 30156 25288
rect 15476 25168 15528 25220
rect 2872 25100 2924 25152
rect 5540 25100 5592 25152
rect 13452 25100 13504 25152
rect 15200 25143 15252 25152
rect 15200 25109 15209 25143
rect 15209 25109 15243 25143
rect 15243 25109 15252 25143
rect 15200 25100 15252 25109
rect 21088 25168 21140 25220
rect 25136 25168 25188 25220
rect 26516 25168 26568 25220
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 31484 25236 31536 25288
rect 16120 25143 16172 25152
rect 16120 25109 16129 25143
rect 16129 25109 16163 25143
rect 16163 25109 16172 25143
rect 16120 25100 16172 25109
rect 22560 25100 22612 25152
rect 27068 25143 27120 25152
rect 27068 25109 27077 25143
rect 27077 25109 27111 25143
rect 27111 25109 27120 25143
rect 27068 25100 27120 25109
rect 30380 25211 30432 25220
rect 30380 25177 30414 25211
rect 30414 25177 30432 25211
rect 30380 25168 30432 25177
rect 31392 25100 31444 25152
rect 9390 24998 9442 25050
rect 9454 24998 9506 25050
rect 9518 24998 9570 25050
rect 9582 24998 9634 25050
rect 9646 24998 9698 25050
rect 17831 24998 17883 25050
rect 17895 24998 17947 25050
rect 17959 24998 18011 25050
rect 18023 24998 18075 25050
rect 18087 24998 18139 25050
rect 26272 24998 26324 25050
rect 26336 24998 26388 25050
rect 26400 24998 26452 25050
rect 26464 24998 26516 25050
rect 26528 24998 26580 25050
rect 34713 24998 34765 25050
rect 34777 24998 34829 25050
rect 34841 24998 34893 25050
rect 34905 24998 34957 25050
rect 34969 24998 35021 25050
rect 12256 24896 12308 24948
rect 15292 24896 15344 24948
rect 17040 24896 17092 24948
rect 23572 24896 23624 24948
rect 25136 24896 25188 24948
rect 31484 24939 31536 24948
rect 31484 24905 31493 24939
rect 31493 24905 31527 24939
rect 31527 24905 31536 24939
rect 31484 24896 31536 24905
rect 5080 24828 5132 24880
rect 3884 24760 3936 24812
rect 4160 24760 4212 24812
rect 6828 24760 6880 24812
rect 7840 24760 7892 24812
rect 12808 24760 12860 24812
rect 2780 24692 2832 24744
rect 4712 24735 4764 24744
rect 4712 24701 4721 24735
rect 4721 24701 4755 24735
rect 4755 24701 4764 24735
rect 4712 24692 4764 24701
rect 8484 24692 8536 24744
rect 4068 24624 4120 24676
rect 4988 24624 5040 24676
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 20628 24828 20680 24880
rect 22100 24828 22152 24880
rect 23664 24871 23716 24880
rect 23664 24837 23673 24871
rect 23673 24837 23707 24871
rect 23707 24837 23716 24871
rect 23664 24828 23716 24837
rect 15384 24760 15436 24769
rect 16304 24760 16356 24812
rect 18236 24760 18288 24812
rect 20996 24803 21048 24812
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 17316 24692 17368 24744
rect 19340 24735 19392 24744
rect 19340 24701 19349 24735
rect 19349 24701 19383 24735
rect 19383 24701 19392 24735
rect 19340 24692 19392 24701
rect 15476 24624 15528 24676
rect 21548 24760 21600 24812
rect 23756 24760 23808 24812
rect 25228 24803 25280 24812
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 25320 24803 25372 24812
rect 25320 24769 25329 24803
rect 25329 24769 25363 24803
rect 25363 24769 25372 24803
rect 27068 24828 27120 24880
rect 27160 24828 27212 24880
rect 25320 24760 25372 24769
rect 28724 24760 28776 24812
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 32312 24760 32364 24812
rect 22192 24692 22244 24744
rect 28172 24692 28224 24744
rect 30104 24735 30156 24744
rect 30104 24701 30113 24735
rect 30113 24701 30147 24735
rect 30147 24701 30156 24735
rect 30104 24692 30156 24701
rect 15016 24556 15068 24608
rect 18052 24556 18104 24608
rect 21272 24624 21324 24676
rect 20444 24556 20496 24608
rect 25044 24624 25096 24676
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 26608 24556 26660 24608
rect 5170 24454 5222 24506
rect 5234 24454 5286 24506
rect 5298 24454 5350 24506
rect 5362 24454 5414 24506
rect 5426 24454 5478 24506
rect 13611 24454 13663 24506
rect 13675 24454 13727 24506
rect 13739 24454 13791 24506
rect 13803 24454 13855 24506
rect 13867 24454 13919 24506
rect 22052 24454 22104 24506
rect 22116 24454 22168 24506
rect 22180 24454 22232 24506
rect 22244 24454 22296 24506
rect 22308 24454 22360 24506
rect 30493 24454 30545 24506
rect 30557 24454 30609 24506
rect 30621 24454 30673 24506
rect 30685 24454 30737 24506
rect 30749 24454 30801 24506
rect 2780 24395 2832 24404
rect 2780 24361 2789 24395
rect 2789 24361 2823 24395
rect 2823 24361 2832 24395
rect 2780 24352 2832 24361
rect 4344 24352 4396 24404
rect 6828 24395 6880 24404
rect 2688 24284 2740 24336
rect 2964 24284 3016 24336
rect 6828 24361 6837 24395
rect 6837 24361 6871 24395
rect 6871 24361 6880 24395
rect 6828 24352 6880 24361
rect 16488 24352 16540 24404
rect 2780 24216 2832 24268
rect 2964 24191 3016 24200
rect 2964 24157 2973 24191
rect 2973 24157 3007 24191
rect 3007 24157 3016 24191
rect 2964 24148 3016 24157
rect 5080 24216 5132 24268
rect 6920 24216 6972 24268
rect 5540 24191 5592 24200
rect 2320 24123 2372 24132
rect 2320 24089 2329 24123
rect 2329 24089 2363 24123
rect 2363 24089 2372 24123
rect 2320 24080 2372 24089
rect 2688 24080 2740 24132
rect 3424 24123 3476 24132
rect 3424 24089 3433 24123
rect 3433 24089 3467 24123
rect 3467 24089 3476 24123
rect 3424 24080 3476 24089
rect 4344 24012 4396 24064
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 15108 24284 15160 24336
rect 20996 24352 21048 24404
rect 13452 24216 13504 24268
rect 7748 24080 7800 24132
rect 9312 24148 9364 24200
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12440 24148 12492 24200
rect 13268 24148 13320 24200
rect 8576 24080 8628 24132
rect 5816 24012 5868 24064
rect 12256 24080 12308 24132
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 15568 24080 15620 24132
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 16396 24148 16448 24200
rect 17960 24148 18012 24200
rect 20904 24216 20956 24268
rect 21088 24216 21140 24268
rect 25228 24352 25280 24404
rect 27528 24352 27580 24404
rect 30380 24352 30432 24404
rect 23480 24284 23532 24336
rect 23756 24284 23808 24336
rect 29000 24284 29052 24336
rect 18696 24080 18748 24132
rect 19708 24080 19760 24132
rect 21272 24148 21324 24200
rect 23572 24080 23624 24132
rect 32404 24216 32456 24268
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 26700 24148 26752 24200
rect 30932 24148 30984 24200
rect 25136 24080 25188 24132
rect 32772 24148 32824 24200
rect 12624 24012 12676 24064
rect 12900 24012 12952 24064
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 17132 24055 17184 24064
rect 17132 24021 17141 24055
rect 17141 24021 17175 24055
rect 17175 24021 17184 24055
rect 17132 24012 17184 24021
rect 17592 24012 17644 24064
rect 24676 24012 24728 24064
rect 25320 24055 25372 24064
rect 25320 24021 25329 24055
rect 25329 24021 25363 24055
rect 25363 24021 25372 24055
rect 25320 24012 25372 24021
rect 31392 24012 31444 24064
rect 9390 23910 9442 23962
rect 9454 23910 9506 23962
rect 9518 23910 9570 23962
rect 9582 23910 9634 23962
rect 9646 23910 9698 23962
rect 17831 23910 17883 23962
rect 17895 23910 17947 23962
rect 17959 23910 18011 23962
rect 18023 23910 18075 23962
rect 18087 23910 18139 23962
rect 26272 23910 26324 23962
rect 26336 23910 26388 23962
rect 26400 23910 26452 23962
rect 26464 23910 26516 23962
rect 26528 23910 26580 23962
rect 34713 23910 34765 23962
rect 34777 23910 34829 23962
rect 34841 23910 34893 23962
rect 34905 23910 34957 23962
rect 34969 23910 35021 23962
rect 2320 23808 2372 23860
rect 7748 23808 7800 23860
rect 3332 23740 3384 23792
rect 3700 23715 3752 23724
rect 3700 23681 3709 23715
rect 3709 23681 3743 23715
rect 3743 23681 3752 23715
rect 3700 23672 3752 23681
rect 5816 23740 5868 23792
rect 8484 23740 8536 23792
rect 15016 23808 15068 23860
rect 15384 23808 15436 23860
rect 16120 23808 16172 23860
rect 19340 23808 19392 23860
rect 20628 23808 20680 23860
rect 30104 23851 30156 23860
rect 4712 23604 4764 23656
rect 5080 23672 5132 23724
rect 7196 23672 7248 23724
rect 20720 23740 20772 23792
rect 21916 23740 21968 23792
rect 30104 23817 30113 23851
rect 30113 23817 30147 23851
rect 30147 23817 30156 23851
rect 30104 23808 30156 23817
rect 25228 23740 25280 23792
rect 28632 23783 28684 23792
rect 28632 23749 28641 23783
rect 28641 23749 28675 23783
rect 28675 23749 28684 23783
rect 28632 23740 28684 23749
rect 6736 23604 6788 23656
rect 7104 23647 7156 23656
rect 7104 23613 7113 23647
rect 7113 23613 7147 23647
rect 7147 23613 7156 23647
rect 7104 23604 7156 23613
rect 3884 23468 3936 23520
rect 4252 23468 4304 23520
rect 4620 23468 4672 23520
rect 12900 23715 12952 23724
rect 7932 23604 7984 23656
rect 9496 23604 9548 23656
rect 8300 23536 8352 23588
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 15476 23672 15528 23724
rect 15844 23672 15896 23724
rect 17132 23672 17184 23724
rect 20444 23715 20496 23724
rect 20444 23681 20453 23715
rect 20453 23681 20487 23715
rect 20487 23681 20496 23715
rect 20444 23672 20496 23681
rect 20904 23672 20956 23724
rect 12256 23647 12308 23656
rect 12256 23613 12265 23647
rect 12265 23613 12299 23647
rect 12299 23613 12308 23647
rect 12256 23604 12308 23613
rect 13176 23647 13228 23656
rect 13176 23613 13185 23647
rect 13185 23613 13219 23647
rect 13219 23613 13228 23647
rect 13176 23604 13228 23613
rect 14740 23604 14792 23656
rect 15200 23647 15252 23656
rect 15200 23613 15209 23647
rect 15209 23613 15243 23647
rect 15243 23613 15252 23647
rect 15200 23604 15252 23613
rect 15292 23647 15344 23656
rect 15292 23613 15301 23647
rect 15301 23613 15335 23647
rect 15335 23613 15344 23647
rect 15292 23604 15344 23613
rect 18420 23604 18472 23656
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 23664 23672 23716 23724
rect 24676 23672 24728 23724
rect 27160 23604 27212 23656
rect 14188 23536 14240 23588
rect 19708 23536 19760 23588
rect 8024 23468 8076 23520
rect 9496 23468 9548 23520
rect 15476 23511 15528 23520
rect 15476 23477 15485 23511
rect 15485 23477 15519 23511
rect 15519 23477 15528 23511
rect 15476 23468 15528 23477
rect 24952 23468 25004 23520
rect 5170 23366 5222 23418
rect 5234 23366 5286 23418
rect 5298 23366 5350 23418
rect 5362 23366 5414 23418
rect 5426 23366 5478 23418
rect 13611 23366 13663 23418
rect 13675 23366 13727 23418
rect 13739 23366 13791 23418
rect 13803 23366 13855 23418
rect 13867 23366 13919 23418
rect 22052 23366 22104 23418
rect 22116 23366 22168 23418
rect 22180 23366 22232 23418
rect 22244 23366 22296 23418
rect 22308 23366 22360 23418
rect 30493 23366 30545 23418
rect 30557 23366 30609 23418
rect 30621 23366 30673 23418
rect 30685 23366 30737 23418
rect 30749 23366 30801 23418
rect 2872 23264 2924 23316
rect 3424 23264 3476 23316
rect 4252 23264 4304 23316
rect 7104 23264 7156 23316
rect 10232 23264 10284 23316
rect 18696 23307 18748 23316
rect 7380 23196 7432 23248
rect 9864 23196 9916 23248
rect 4160 23128 4212 23180
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 7380 23103 7432 23112
rect 7380 23069 7415 23103
rect 7415 23069 7432 23103
rect 7564 23103 7616 23112
rect 7380 23060 7432 23069
rect 7564 23069 7573 23103
rect 7573 23069 7607 23103
rect 7607 23069 7616 23103
rect 7564 23060 7616 23069
rect 8024 23128 8076 23180
rect 5080 22992 5132 23044
rect 7196 23035 7248 23044
rect 7196 23001 7205 23035
rect 7205 23001 7239 23035
rect 7239 23001 7248 23035
rect 7196 22992 7248 23001
rect 7748 22992 7800 23044
rect 3976 22967 4028 22976
rect 3976 22933 3985 22967
rect 3985 22933 4019 22967
rect 4019 22933 4028 22967
rect 3976 22924 4028 22933
rect 4712 22924 4764 22976
rect 6736 22924 6788 22976
rect 8392 23103 8444 23112
rect 8392 23069 8401 23103
rect 8401 23069 8435 23103
rect 8435 23069 8444 23103
rect 8392 23060 8444 23069
rect 9496 23128 9548 23180
rect 10048 23128 10100 23180
rect 8668 23060 8720 23112
rect 9404 23103 9456 23112
rect 9404 23069 9413 23103
rect 9413 23069 9447 23103
rect 9447 23069 9456 23103
rect 9404 23060 9456 23069
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 9772 22992 9824 23044
rect 11888 22992 11940 23044
rect 18696 23273 18705 23307
rect 18705 23273 18739 23307
rect 18739 23273 18748 23307
rect 18696 23264 18748 23273
rect 21916 23307 21968 23316
rect 21916 23273 21925 23307
rect 21925 23273 21959 23307
rect 21959 23273 21968 23307
rect 21916 23264 21968 23273
rect 31852 23264 31904 23316
rect 33140 23264 33192 23316
rect 15200 23171 15252 23180
rect 15200 23137 15209 23171
rect 15209 23137 15243 23171
rect 15243 23137 15252 23171
rect 15200 23128 15252 23137
rect 15384 23196 15436 23248
rect 19616 23196 19668 23248
rect 19984 23196 20036 23248
rect 28724 23196 28776 23248
rect 15476 23128 15528 23180
rect 17316 23171 17368 23180
rect 17316 23137 17325 23171
rect 17325 23137 17359 23171
rect 17359 23137 17368 23171
rect 17316 23128 17368 23137
rect 24952 23171 25004 23180
rect 24952 23137 24961 23171
rect 24961 23137 24995 23171
rect 24995 23137 25004 23171
rect 24952 23128 25004 23137
rect 25320 23171 25372 23180
rect 25320 23137 25329 23171
rect 25329 23137 25363 23171
rect 25363 23137 25372 23171
rect 25320 23128 25372 23137
rect 31024 23128 31076 23180
rect 32680 23171 32732 23180
rect 32680 23137 32689 23171
rect 32689 23137 32723 23171
rect 32723 23137 32732 23171
rect 32680 23128 32732 23137
rect 33140 23171 33192 23180
rect 33140 23137 33149 23171
rect 33149 23137 33183 23171
rect 33183 23137 33192 23171
rect 33140 23128 33192 23137
rect 14004 23060 14056 23112
rect 15016 23060 15068 23112
rect 17592 23103 17644 23112
rect 17592 23069 17626 23103
rect 17626 23069 17644 23103
rect 10324 22967 10376 22976
rect 10324 22933 10333 22967
rect 10333 22933 10367 22967
rect 10367 22933 10376 22967
rect 10324 22924 10376 22933
rect 10416 22924 10468 22976
rect 14740 22992 14792 23044
rect 17592 23060 17644 23069
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 20812 23060 20864 23112
rect 22744 23060 22796 23112
rect 27528 23103 27580 23112
rect 27528 23069 27537 23103
rect 27537 23069 27571 23103
rect 27571 23069 27580 23103
rect 27528 23060 27580 23069
rect 27988 23103 28040 23112
rect 27988 23069 27997 23103
rect 27997 23069 28031 23103
rect 28031 23069 28040 23103
rect 27988 23060 28040 23069
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 31760 23103 31812 23112
rect 31760 23069 31769 23103
rect 31769 23069 31803 23103
rect 31803 23069 31812 23103
rect 31760 23060 31812 23069
rect 32036 23103 32088 23112
rect 32036 23069 32045 23103
rect 32045 23069 32079 23103
rect 32079 23069 32088 23103
rect 32036 23060 32088 23069
rect 32404 23060 32456 23112
rect 33324 23060 33376 23112
rect 27620 22992 27672 23044
rect 28540 22992 28592 23044
rect 14648 22924 14700 22976
rect 24860 22924 24912 22976
rect 24952 22924 25004 22976
rect 25228 22967 25280 22976
rect 25228 22933 25237 22967
rect 25237 22933 25271 22967
rect 25271 22933 25280 22967
rect 25228 22924 25280 22933
rect 29736 22924 29788 22976
rect 33508 22924 33560 22976
rect 9390 22822 9442 22874
rect 9454 22822 9506 22874
rect 9518 22822 9570 22874
rect 9582 22822 9634 22874
rect 9646 22822 9698 22874
rect 17831 22822 17883 22874
rect 17895 22822 17947 22874
rect 17959 22822 18011 22874
rect 18023 22822 18075 22874
rect 18087 22822 18139 22874
rect 26272 22822 26324 22874
rect 26336 22822 26388 22874
rect 26400 22822 26452 22874
rect 26464 22822 26516 22874
rect 26528 22822 26580 22874
rect 34713 22822 34765 22874
rect 34777 22822 34829 22874
rect 34841 22822 34893 22874
rect 34905 22822 34957 22874
rect 34969 22822 35021 22874
rect 7564 22720 7616 22772
rect 9312 22720 9364 22772
rect 7104 22652 7156 22704
rect 8300 22695 8352 22704
rect 8300 22661 8309 22695
rect 8309 22661 8343 22695
rect 8343 22661 8352 22695
rect 8300 22652 8352 22661
rect 8484 22695 8536 22704
rect 8484 22661 8493 22695
rect 8493 22661 8527 22695
rect 8527 22661 8536 22695
rect 8484 22652 8536 22661
rect 9772 22652 9824 22704
rect 10324 22720 10376 22772
rect 10784 22720 10836 22772
rect 4344 22584 4396 22636
rect 7472 22584 7524 22636
rect 3700 22516 3752 22568
rect 8392 22516 8444 22568
rect 8668 22448 8720 22500
rect 10416 22584 10468 22636
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 12440 22584 12492 22636
rect 12624 22584 12676 22636
rect 11796 22516 11848 22568
rect 5080 22380 5132 22432
rect 9220 22380 9272 22432
rect 11980 22448 12032 22500
rect 12900 22448 12952 22500
rect 13452 22584 13504 22636
rect 31852 22720 31904 22772
rect 32036 22720 32088 22772
rect 14740 22652 14792 22704
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 15476 22627 15528 22636
rect 14188 22516 14240 22568
rect 15476 22593 15485 22627
rect 15485 22593 15519 22627
rect 15519 22593 15528 22627
rect 15476 22584 15528 22593
rect 15568 22627 15620 22636
rect 15568 22593 15577 22627
rect 15577 22593 15611 22627
rect 15611 22593 15620 22627
rect 15568 22584 15620 22593
rect 16396 22584 16448 22636
rect 17132 22584 17184 22636
rect 18696 22584 18748 22636
rect 19984 22627 20036 22636
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 18052 22448 18104 22500
rect 19340 22516 19392 22568
rect 20536 22584 20588 22636
rect 20996 22584 21048 22636
rect 21824 22584 21876 22636
rect 25228 22695 25280 22704
rect 25228 22661 25237 22695
rect 25237 22661 25271 22695
rect 25271 22661 25280 22695
rect 25228 22652 25280 22661
rect 28264 22652 28316 22704
rect 10324 22380 10376 22432
rect 12992 22380 13044 22432
rect 17960 22423 18012 22432
rect 17960 22389 17969 22423
rect 17969 22389 18003 22423
rect 18003 22389 18012 22423
rect 17960 22380 18012 22389
rect 19800 22423 19852 22432
rect 19800 22389 19809 22423
rect 19809 22389 19843 22423
rect 19843 22389 19852 22423
rect 19800 22380 19852 22389
rect 27160 22584 27212 22636
rect 27988 22627 28040 22636
rect 27988 22593 27997 22627
rect 27997 22593 28031 22627
rect 28031 22593 28040 22627
rect 27988 22584 28040 22593
rect 28540 22584 28592 22636
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 26148 22516 26200 22568
rect 26976 22516 27028 22568
rect 29736 22559 29788 22568
rect 29736 22525 29745 22559
rect 29745 22525 29779 22559
rect 29779 22525 29788 22559
rect 29736 22516 29788 22525
rect 33140 22652 33192 22704
rect 33508 22695 33560 22704
rect 33508 22661 33517 22695
rect 33517 22661 33551 22695
rect 33551 22661 33560 22695
rect 33508 22652 33560 22661
rect 31024 22627 31076 22636
rect 31024 22593 31033 22627
rect 31033 22593 31067 22627
rect 31067 22593 31076 22627
rect 31024 22584 31076 22593
rect 31392 22584 31444 22636
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 33692 22627 33744 22636
rect 33692 22593 33701 22627
rect 33701 22593 33735 22627
rect 33735 22593 33744 22627
rect 33692 22584 33744 22593
rect 31116 22559 31168 22568
rect 27988 22448 28040 22500
rect 30104 22491 30156 22500
rect 30104 22457 30113 22491
rect 30113 22457 30147 22491
rect 30147 22457 30156 22491
rect 30104 22448 30156 22457
rect 23020 22380 23072 22432
rect 24584 22423 24636 22432
rect 24584 22389 24593 22423
rect 24593 22389 24627 22423
rect 24627 22389 24636 22423
rect 24584 22380 24636 22389
rect 26976 22380 27028 22432
rect 30380 22380 30432 22432
rect 31116 22525 31125 22559
rect 31125 22525 31159 22559
rect 31159 22525 31168 22559
rect 31116 22516 31168 22525
rect 31300 22559 31352 22568
rect 31300 22525 31310 22559
rect 31310 22525 31344 22559
rect 31344 22525 31352 22559
rect 31300 22516 31352 22525
rect 32404 22516 32456 22568
rect 33324 22516 33376 22568
rect 5170 22278 5222 22330
rect 5234 22278 5286 22330
rect 5298 22278 5350 22330
rect 5362 22278 5414 22330
rect 5426 22278 5478 22330
rect 13611 22278 13663 22330
rect 13675 22278 13727 22330
rect 13739 22278 13791 22330
rect 13803 22278 13855 22330
rect 13867 22278 13919 22330
rect 22052 22278 22104 22330
rect 22116 22278 22168 22330
rect 22180 22278 22232 22330
rect 22244 22278 22296 22330
rect 22308 22278 22360 22330
rect 30493 22278 30545 22330
rect 30557 22278 30609 22330
rect 30621 22278 30673 22330
rect 30685 22278 30737 22330
rect 30749 22278 30801 22330
rect 4896 22176 4948 22228
rect 9864 22176 9916 22228
rect 10232 22219 10284 22228
rect 10232 22185 10241 22219
rect 10241 22185 10275 22219
rect 10275 22185 10284 22219
rect 10232 22176 10284 22185
rect 10968 22176 11020 22228
rect 11704 22219 11756 22228
rect 11704 22185 11725 22219
rect 11725 22185 11756 22219
rect 11704 22176 11756 22185
rect 16396 22176 16448 22228
rect 19984 22176 20036 22228
rect 23020 22219 23072 22228
rect 23020 22185 23029 22219
rect 23029 22185 23063 22219
rect 23063 22185 23072 22219
rect 23020 22176 23072 22185
rect 13360 22108 13412 22160
rect 17960 22108 18012 22160
rect 22652 22108 22704 22160
rect 23848 22176 23900 22228
rect 24768 22176 24820 22228
rect 28448 22176 28500 22228
rect 33692 22176 33744 22228
rect 11612 22040 11664 22092
rect 12072 22040 12124 22092
rect 20076 22040 20128 22092
rect 24952 22108 25004 22160
rect 25228 22040 25280 22092
rect 26148 22040 26200 22092
rect 26976 22083 27028 22092
rect 7196 22015 7248 22024
rect 7196 21981 7205 22015
rect 7205 21981 7239 22015
rect 7239 21981 7248 22015
rect 7196 21972 7248 21981
rect 7472 21972 7524 22024
rect 9312 21972 9364 22024
rect 12716 22015 12768 22024
rect 12716 21981 12725 22015
rect 12725 21981 12759 22015
rect 12759 21981 12768 22015
rect 12716 21972 12768 21981
rect 12900 22015 12952 22024
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 18052 21972 18104 22024
rect 18420 21972 18472 22024
rect 19432 21972 19484 22024
rect 19524 21972 19576 22024
rect 20720 21972 20772 22024
rect 22928 21972 22980 22024
rect 24584 21972 24636 22024
rect 25964 21972 26016 22024
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 30380 22108 30432 22160
rect 33140 22083 33192 22092
rect 33140 22049 33149 22083
rect 33149 22049 33183 22083
rect 33183 22049 33192 22083
rect 33140 22040 33192 22049
rect 26332 21972 26384 22024
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 31024 22015 31076 22024
rect 11704 21904 11756 21956
rect 19340 21904 19392 21956
rect 19892 21904 19944 21956
rect 6920 21836 6972 21888
rect 7196 21879 7248 21888
rect 7196 21845 7205 21879
rect 7205 21845 7239 21879
rect 7239 21845 7248 21879
rect 7196 21836 7248 21845
rect 8392 21836 8444 21888
rect 9036 21836 9088 21888
rect 10692 21836 10744 21888
rect 19616 21836 19668 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 23112 21904 23164 21956
rect 24952 21836 25004 21888
rect 25044 21836 25096 21888
rect 27528 21904 27580 21956
rect 28448 21947 28500 21956
rect 28448 21913 28457 21947
rect 28457 21913 28491 21947
rect 28491 21913 28500 21947
rect 28448 21904 28500 21913
rect 31024 21981 31033 22015
rect 31033 21981 31067 22015
rect 31067 21981 31076 22015
rect 31392 22015 31444 22024
rect 31024 21972 31076 21981
rect 30288 21904 30340 21956
rect 31392 21981 31401 22015
rect 31401 21981 31435 22015
rect 31435 21981 31444 22015
rect 31392 21972 31444 21981
rect 31576 22015 31628 22024
rect 31576 21981 31585 22015
rect 31585 21981 31619 22015
rect 31619 21981 31628 22015
rect 31576 21972 31628 21981
rect 32404 22015 32456 22024
rect 32404 21981 32413 22015
rect 32413 21981 32447 22015
rect 32447 21981 32456 22015
rect 32404 21972 32456 21981
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 29736 21879 29788 21888
rect 29736 21845 29745 21879
rect 29745 21845 29779 21879
rect 29779 21845 29788 21879
rect 29736 21836 29788 21845
rect 9390 21734 9442 21786
rect 9454 21734 9506 21786
rect 9518 21734 9570 21786
rect 9582 21734 9634 21786
rect 9646 21734 9698 21786
rect 17831 21734 17883 21786
rect 17895 21734 17947 21786
rect 17959 21734 18011 21786
rect 18023 21734 18075 21786
rect 18087 21734 18139 21786
rect 26272 21734 26324 21786
rect 26336 21734 26388 21786
rect 26400 21734 26452 21786
rect 26464 21734 26516 21786
rect 26528 21734 26580 21786
rect 34713 21734 34765 21786
rect 34777 21734 34829 21786
rect 34841 21734 34893 21786
rect 34905 21734 34957 21786
rect 34969 21734 35021 21786
rect 12716 21632 12768 21684
rect 27160 21675 27212 21684
rect 11704 21607 11756 21616
rect 11704 21573 11713 21607
rect 11713 21573 11747 21607
rect 11747 21573 11756 21607
rect 11704 21564 11756 21573
rect 20444 21564 20496 21616
rect 3976 21496 4028 21548
rect 4160 21496 4212 21548
rect 11796 21539 11848 21548
rect 11796 21505 11805 21539
rect 11805 21505 11839 21539
rect 11839 21505 11848 21539
rect 11796 21496 11848 21505
rect 11980 21496 12032 21548
rect 12348 21496 12400 21548
rect 14004 21496 14056 21548
rect 16028 21496 16080 21548
rect 16488 21496 16540 21548
rect 19432 21539 19484 21548
rect 19432 21505 19441 21539
rect 19441 21505 19475 21539
rect 19475 21505 19484 21539
rect 19432 21496 19484 21505
rect 19800 21539 19852 21548
rect 19800 21505 19809 21539
rect 19809 21505 19843 21539
rect 19843 21505 19852 21539
rect 19800 21496 19852 21505
rect 23112 21564 23164 21616
rect 22284 21539 22336 21548
rect 2964 21471 3016 21480
rect 2964 21437 2973 21471
rect 2973 21437 3007 21471
rect 3007 21437 3016 21471
rect 2964 21428 3016 21437
rect 10968 21428 11020 21480
rect 19616 21428 19668 21480
rect 4068 21360 4120 21412
rect 3056 21335 3108 21344
rect 3056 21301 3065 21335
rect 3065 21301 3099 21335
rect 3099 21301 3108 21335
rect 3056 21292 3108 21301
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 16856 21292 16908 21344
rect 19892 21292 19944 21344
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 30104 21632 30156 21684
rect 30288 21675 30340 21684
rect 30288 21641 30297 21675
rect 30297 21641 30331 21675
rect 30331 21641 30340 21675
rect 30288 21632 30340 21641
rect 31760 21632 31812 21684
rect 27988 21496 28040 21548
rect 28448 21564 28500 21616
rect 31024 21564 31076 21616
rect 31392 21564 31444 21616
rect 29736 21496 29788 21548
rect 30380 21496 30432 21548
rect 31116 21496 31168 21548
rect 32588 21496 32640 21548
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 23572 21428 23624 21480
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 23848 21292 23900 21344
rect 23940 21292 23992 21344
rect 30104 21360 30156 21412
rect 32220 21360 32272 21412
rect 27896 21292 27948 21344
rect 28448 21292 28500 21344
rect 5170 21190 5222 21242
rect 5234 21190 5286 21242
rect 5298 21190 5350 21242
rect 5362 21190 5414 21242
rect 5426 21190 5478 21242
rect 13611 21190 13663 21242
rect 13675 21190 13727 21242
rect 13739 21190 13791 21242
rect 13803 21190 13855 21242
rect 13867 21190 13919 21242
rect 22052 21190 22104 21242
rect 22116 21190 22168 21242
rect 22180 21190 22232 21242
rect 22244 21190 22296 21242
rect 22308 21190 22360 21242
rect 30493 21190 30545 21242
rect 30557 21190 30609 21242
rect 30621 21190 30673 21242
rect 30685 21190 30737 21242
rect 30749 21190 30801 21242
rect 12900 21088 12952 21140
rect 7472 20952 7524 21004
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 3700 20884 3752 20936
rect 7288 20884 7340 20936
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 10324 20884 10376 20936
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 13452 20884 13504 20936
rect 14464 20884 14516 20936
rect 17316 21088 17368 21140
rect 21272 21131 21324 21140
rect 21272 21097 21281 21131
rect 21281 21097 21315 21131
rect 21315 21097 21324 21131
rect 21272 21088 21324 21097
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 24952 21088 25004 21140
rect 30932 21088 30984 21140
rect 31944 21088 31996 21140
rect 32404 21131 32456 21140
rect 32404 21097 32413 21131
rect 32413 21097 32447 21131
rect 32447 21097 32456 21131
rect 32404 21088 32456 21097
rect 19892 20952 19944 21004
rect 19984 20952 20036 21004
rect 21180 20952 21232 21004
rect 18328 20884 18380 20936
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 3148 20748 3200 20800
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 10232 20791 10284 20800
rect 10232 20757 10241 20791
rect 10241 20757 10275 20791
rect 10275 20757 10284 20791
rect 10232 20748 10284 20757
rect 10968 20748 11020 20800
rect 14372 20791 14424 20800
rect 14372 20757 14381 20791
rect 14381 20757 14415 20791
rect 14415 20757 14424 20791
rect 14372 20748 14424 20757
rect 19708 20816 19760 20868
rect 23940 20927 23992 20936
rect 23940 20893 23949 20927
rect 23949 20893 23983 20927
rect 23983 20893 23992 20927
rect 23940 20884 23992 20893
rect 24952 20952 25004 21004
rect 31116 20952 31168 21004
rect 23388 20816 23440 20868
rect 25136 20884 25188 20936
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 32496 20927 32548 20936
rect 32496 20893 32505 20927
rect 32505 20893 32539 20927
rect 32539 20893 32548 20927
rect 32496 20884 32548 20893
rect 32956 20927 33008 20936
rect 32956 20893 32965 20927
rect 32965 20893 32999 20927
rect 32999 20893 33008 20927
rect 32956 20884 33008 20893
rect 33048 20884 33100 20936
rect 32772 20816 32824 20868
rect 22560 20748 22612 20800
rect 25228 20748 25280 20800
rect 9390 20646 9442 20698
rect 9454 20646 9506 20698
rect 9518 20646 9570 20698
rect 9582 20646 9634 20698
rect 9646 20646 9698 20698
rect 17831 20646 17883 20698
rect 17895 20646 17947 20698
rect 17959 20646 18011 20698
rect 18023 20646 18075 20698
rect 18087 20646 18139 20698
rect 26272 20646 26324 20698
rect 26336 20646 26388 20698
rect 26400 20646 26452 20698
rect 26464 20646 26516 20698
rect 26528 20646 26580 20698
rect 34713 20646 34765 20698
rect 34777 20646 34829 20698
rect 34841 20646 34893 20698
rect 34905 20646 34957 20698
rect 34969 20646 35021 20698
rect 8300 20544 8352 20596
rect 3608 20519 3660 20528
rect 3608 20485 3617 20519
rect 3617 20485 3651 20519
rect 3651 20485 3660 20519
rect 3608 20476 3660 20485
rect 7748 20476 7800 20528
rect 3148 20451 3200 20460
rect 3148 20417 3157 20451
rect 3157 20417 3191 20451
rect 3191 20417 3200 20451
rect 3148 20408 3200 20417
rect 3976 20408 4028 20460
rect 4528 20408 4580 20460
rect 7288 20408 7340 20460
rect 8024 20408 8076 20460
rect 8484 20451 8536 20460
rect 3056 20340 3108 20392
rect 3424 20340 3476 20392
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 10232 20408 10284 20460
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 14188 20544 14240 20596
rect 14372 20476 14424 20528
rect 2412 20272 2464 20324
rect 8944 20340 8996 20392
rect 10324 20383 10376 20392
rect 10324 20349 10333 20383
rect 10333 20349 10367 20383
rect 10367 20349 10376 20383
rect 10324 20340 10376 20349
rect 7840 20272 7892 20324
rect 13360 20340 13412 20392
rect 16212 20476 16264 20528
rect 15660 20451 15712 20460
rect 12900 20272 12952 20324
rect 14188 20340 14240 20392
rect 14648 20383 14700 20392
rect 14648 20349 14657 20383
rect 14657 20349 14691 20383
rect 14691 20349 14700 20383
rect 14648 20340 14700 20349
rect 14740 20340 14792 20392
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 16028 20408 16080 20460
rect 19064 20544 19116 20596
rect 19616 20544 19668 20596
rect 19800 20544 19852 20596
rect 18788 20476 18840 20528
rect 22744 20544 22796 20596
rect 31576 20587 31628 20596
rect 31576 20553 31585 20587
rect 31585 20553 31619 20587
rect 31619 20553 31628 20587
rect 31576 20544 31628 20553
rect 32588 20587 32640 20596
rect 32588 20553 32597 20587
rect 32597 20553 32631 20587
rect 32631 20553 32640 20587
rect 32588 20544 32640 20553
rect 22376 20476 22428 20528
rect 18972 20408 19024 20460
rect 19156 20408 19208 20460
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 19708 20408 19760 20460
rect 20444 20408 20496 20460
rect 20628 20408 20680 20460
rect 21088 20408 21140 20460
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 27988 20408 28040 20417
rect 19800 20340 19852 20392
rect 22560 20340 22612 20392
rect 25872 20340 25924 20392
rect 27896 20383 27948 20392
rect 27896 20349 27905 20383
rect 27905 20349 27939 20383
rect 27939 20349 27948 20383
rect 27896 20340 27948 20349
rect 32404 20408 32456 20460
rect 32772 20451 32824 20460
rect 32772 20417 32781 20451
rect 32781 20417 32815 20451
rect 32815 20417 32824 20451
rect 32772 20408 32824 20417
rect 33048 20451 33100 20460
rect 33048 20417 33057 20451
rect 33057 20417 33091 20451
rect 33091 20417 33100 20451
rect 33048 20408 33100 20417
rect 31944 20340 31996 20392
rect 16672 20272 16724 20324
rect 20260 20272 20312 20324
rect 21364 20272 21416 20324
rect 32312 20272 32364 20324
rect 32956 20315 33008 20324
rect 32956 20281 32965 20315
rect 32965 20281 32999 20315
rect 32999 20281 33008 20315
rect 32956 20272 33008 20281
rect 2964 20247 3016 20256
rect 2964 20213 2973 20247
rect 2973 20213 3007 20247
rect 3007 20213 3016 20247
rect 2964 20204 3016 20213
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 19064 20204 19116 20256
rect 19708 20204 19760 20256
rect 21732 20204 21784 20256
rect 28080 20204 28132 20256
rect 5170 20102 5222 20154
rect 5234 20102 5286 20154
rect 5298 20102 5350 20154
rect 5362 20102 5414 20154
rect 5426 20102 5478 20154
rect 13611 20102 13663 20154
rect 13675 20102 13727 20154
rect 13739 20102 13791 20154
rect 13803 20102 13855 20154
rect 13867 20102 13919 20154
rect 22052 20102 22104 20154
rect 22116 20102 22168 20154
rect 22180 20102 22232 20154
rect 22244 20102 22296 20154
rect 22308 20102 22360 20154
rect 30493 20102 30545 20154
rect 30557 20102 30609 20154
rect 30621 20102 30673 20154
rect 30685 20102 30737 20154
rect 30749 20102 30801 20154
rect 3976 20043 4028 20052
rect 3976 20009 3985 20043
rect 3985 20009 4019 20043
rect 4019 20009 4028 20043
rect 3976 20000 4028 20009
rect 4160 20000 4212 20052
rect 2412 19907 2464 19916
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2412 19864 2464 19873
rect 3240 19907 3292 19916
rect 3240 19873 3249 19907
rect 3249 19873 3283 19907
rect 3283 19873 3292 19907
rect 7472 20000 7524 20052
rect 7104 19975 7156 19984
rect 7104 19941 7113 19975
rect 7113 19941 7147 19975
rect 7147 19941 7156 19975
rect 7104 19932 7156 19941
rect 3240 19864 3292 19873
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 3700 19796 3752 19848
rect 4160 19839 4212 19848
rect 4160 19805 4169 19839
rect 4169 19805 4203 19839
rect 4203 19805 4212 19839
rect 4160 19796 4212 19805
rect 7656 20000 7708 20052
rect 15660 20000 15712 20052
rect 19248 20000 19300 20052
rect 19340 20000 19392 20052
rect 19524 20000 19576 20052
rect 20076 20043 20128 20052
rect 20076 20009 20085 20043
rect 20085 20009 20119 20043
rect 20119 20009 20128 20043
rect 20076 20000 20128 20009
rect 7748 19975 7800 19984
rect 7748 19941 7757 19975
rect 7757 19941 7791 19975
rect 7791 19941 7800 19975
rect 7748 19932 7800 19941
rect 14740 19932 14792 19984
rect 14832 19932 14884 19984
rect 21364 19932 21416 19984
rect 32312 19975 32364 19984
rect 32312 19941 32321 19975
rect 32321 19941 32355 19975
rect 32355 19941 32364 19975
rect 32312 19932 32364 19941
rect 5356 19839 5408 19848
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 3332 19728 3384 19780
rect 4252 19771 4304 19780
rect 4252 19737 4261 19771
rect 4261 19737 4295 19771
rect 4295 19737 4304 19771
rect 4252 19728 4304 19737
rect 5080 19771 5132 19780
rect 5080 19737 5089 19771
rect 5089 19737 5123 19771
rect 5123 19737 5132 19771
rect 5080 19728 5132 19737
rect 5264 19771 5316 19780
rect 5264 19737 5273 19771
rect 5273 19737 5307 19771
rect 5307 19737 5316 19771
rect 5264 19728 5316 19737
rect 6552 19660 6604 19712
rect 7380 19796 7432 19848
rect 8024 19839 8076 19848
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 8484 19796 8536 19848
rect 9956 19796 10008 19848
rect 10324 19796 10376 19848
rect 10968 19864 11020 19916
rect 7288 19728 7340 19780
rect 8944 19728 8996 19780
rect 9772 19728 9824 19780
rect 10232 19728 10284 19780
rect 10692 19728 10744 19780
rect 12716 19796 12768 19848
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13452 19796 13504 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 14556 19796 14608 19848
rect 19340 19864 19392 19916
rect 15844 19796 15896 19848
rect 15660 19771 15712 19780
rect 15660 19737 15669 19771
rect 15669 19737 15703 19771
rect 15703 19737 15712 19771
rect 15660 19728 15712 19737
rect 17132 19728 17184 19780
rect 7840 19660 7892 19712
rect 11520 19703 11572 19712
rect 11520 19669 11529 19703
rect 11529 19669 11563 19703
rect 11563 19669 11572 19703
rect 11520 19660 11572 19669
rect 19524 19839 19576 19848
rect 19524 19805 19534 19839
rect 19534 19805 19568 19839
rect 19568 19805 19576 19839
rect 20628 19864 20680 19916
rect 23204 19864 23256 19916
rect 19524 19796 19576 19805
rect 19616 19728 19668 19780
rect 20168 19796 20220 19848
rect 20076 19728 20128 19780
rect 21088 19796 21140 19848
rect 31944 19839 31996 19848
rect 31944 19805 31953 19839
rect 31953 19805 31987 19839
rect 31987 19805 31996 19839
rect 31944 19796 31996 19805
rect 32496 19864 32548 19916
rect 32220 19796 32272 19848
rect 20812 19771 20864 19780
rect 20812 19737 20821 19771
rect 20821 19737 20855 19771
rect 20855 19737 20864 19771
rect 20812 19728 20864 19737
rect 21732 19728 21784 19780
rect 19892 19660 19944 19712
rect 32404 19660 32456 19712
rect 9390 19558 9442 19610
rect 9454 19558 9506 19610
rect 9518 19558 9570 19610
rect 9582 19558 9634 19610
rect 9646 19558 9698 19610
rect 17831 19558 17883 19610
rect 17895 19558 17947 19610
rect 17959 19558 18011 19610
rect 18023 19558 18075 19610
rect 18087 19558 18139 19610
rect 26272 19558 26324 19610
rect 26336 19558 26388 19610
rect 26400 19558 26452 19610
rect 26464 19558 26516 19610
rect 26528 19558 26580 19610
rect 34713 19558 34765 19610
rect 34777 19558 34829 19610
rect 34841 19558 34893 19610
rect 34905 19558 34957 19610
rect 34969 19558 35021 19610
rect 1860 19456 1912 19508
rect 4528 19456 4580 19508
rect 5080 19456 5132 19508
rect 19524 19456 19576 19508
rect 19800 19456 19852 19508
rect 29184 19456 29236 19508
rect 32220 19456 32272 19508
rect 32588 19456 32640 19508
rect 33048 19456 33100 19508
rect 2964 19388 3016 19440
rect 3516 19320 3568 19372
rect 3884 19320 3936 19372
rect 4620 19363 4672 19372
rect 4620 19329 4629 19363
rect 4629 19329 4663 19363
rect 4663 19329 4672 19363
rect 4620 19320 4672 19329
rect 6644 19320 6696 19372
rect 16028 19388 16080 19440
rect 7656 19320 7708 19372
rect 8944 19320 8996 19372
rect 9772 19320 9824 19372
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 13360 19320 13412 19372
rect 17132 19320 17184 19372
rect 19432 19388 19484 19440
rect 25228 19388 25280 19440
rect 28172 19388 28224 19440
rect 19064 19320 19116 19372
rect 23204 19320 23256 19372
rect 27252 19363 27304 19372
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 27896 19320 27948 19372
rect 29000 19363 29052 19372
rect 29000 19329 29009 19363
rect 29009 19329 29043 19363
rect 29043 19329 29052 19363
rect 29000 19320 29052 19329
rect 29368 19363 29420 19372
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 31944 19388 31996 19440
rect 31392 19363 31444 19372
rect 31392 19329 31401 19363
rect 31401 19329 31435 19363
rect 31435 19329 31444 19363
rect 31392 19320 31444 19329
rect 32404 19320 32456 19372
rect 4252 19116 4304 19168
rect 11060 19252 11112 19304
rect 11520 19252 11572 19304
rect 14740 19252 14792 19304
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 28540 19252 28592 19304
rect 29276 19295 29328 19304
rect 29276 19261 29285 19295
rect 29285 19261 29319 19295
rect 29319 19261 29328 19295
rect 29276 19252 29328 19261
rect 10140 19184 10192 19236
rect 32680 19184 32732 19236
rect 8116 19116 8168 19168
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 10232 19159 10284 19168
rect 10232 19125 10241 19159
rect 10241 19125 10275 19159
rect 10275 19125 10284 19159
rect 10232 19116 10284 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 19156 19116 19208 19168
rect 20996 19116 21048 19168
rect 27344 19159 27396 19168
rect 27344 19125 27353 19159
rect 27353 19125 27387 19159
rect 27387 19125 27396 19159
rect 27344 19116 27396 19125
rect 5170 19014 5222 19066
rect 5234 19014 5286 19066
rect 5298 19014 5350 19066
rect 5362 19014 5414 19066
rect 5426 19014 5478 19066
rect 13611 19014 13663 19066
rect 13675 19014 13727 19066
rect 13739 19014 13791 19066
rect 13803 19014 13855 19066
rect 13867 19014 13919 19066
rect 22052 19014 22104 19066
rect 22116 19014 22168 19066
rect 22180 19014 22232 19066
rect 22244 19014 22296 19066
rect 22308 19014 22360 19066
rect 30493 19014 30545 19066
rect 30557 19014 30609 19066
rect 30621 19014 30673 19066
rect 30685 19014 30737 19066
rect 30749 19014 30801 19066
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 14648 18912 14700 18964
rect 16672 18955 16724 18964
rect 2964 18844 3016 18896
rect 7104 18776 7156 18828
rect 8484 18844 8536 18896
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 19340 18912 19392 18964
rect 19616 18912 19668 18964
rect 25872 18955 25924 18964
rect 25872 18921 25881 18955
rect 25881 18921 25915 18955
rect 25915 18921 25924 18955
rect 25872 18912 25924 18921
rect 33324 18912 33376 18964
rect 9128 18776 9180 18828
rect 27712 18844 27764 18896
rect 32772 18844 32824 18896
rect 27344 18776 27396 18828
rect 32404 18776 32456 18828
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 10232 18708 10284 18760
rect 3240 18640 3292 18692
rect 7196 18640 7248 18692
rect 8116 18640 8168 18692
rect 10692 18708 10744 18760
rect 12440 18708 12492 18760
rect 14740 18708 14792 18760
rect 15384 18708 15436 18760
rect 19432 18751 19484 18760
rect 19432 18717 19441 18751
rect 19441 18717 19475 18751
rect 19475 18717 19484 18751
rect 19432 18708 19484 18717
rect 12348 18640 12400 18692
rect 15200 18572 15252 18624
rect 15752 18640 15804 18692
rect 19340 18640 19392 18692
rect 20904 18708 20956 18760
rect 23480 18708 23532 18760
rect 23848 18708 23900 18760
rect 24768 18751 24820 18760
rect 19708 18683 19760 18692
rect 19708 18649 19742 18683
rect 19742 18649 19760 18683
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 25136 18708 25188 18760
rect 25964 18708 26016 18760
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 19708 18640 19760 18649
rect 25688 18640 25740 18692
rect 27252 18708 27304 18760
rect 27896 18751 27948 18760
rect 27896 18717 27905 18751
rect 27905 18717 27939 18751
rect 27939 18717 27948 18751
rect 27896 18708 27948 18717
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 28632 18708 28684 18760
rect 29276 18708 29328 18760
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 30104 18751 30156 18760
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 32036 18751 32088 18760
rect 32036 18717 32045 18751
rect 32045 18717 32079 18751
rect 32079 18717 32088 18751
rect 32036 18708 32088 18717
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 16948 18572 17000 18624
rect 18512 18615 18564 18624
rect 18512 18581 18521 18615
rect 18521 18581 18555 18615
rect 18555 18581 18564 18615
rect 18512 18572 18564 18581
rect 19616 18572 19668 18624
rect 20076 18572 20128 18624
rect 23572 18615 23624 18624
rect 23572 18581 23581 18615
rect 23581 18581 23615 18615
rect 23615 18581 23624 18615
rect 23572 18572 23624 18581
rect 24400 18572 24452 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 26240 18572 26292 18624
rect 27068 18572 27120 18624
rect 29368 18640 29420 18692
rect 28356 18615 28408 18624
rect 28356 18581 28365 18615
rect 28365 18581 28399 18615
rect 28399 18581 28408 18615
rect 28356 18572 28408 18581
rect 9390 18470 9442 18522
rect 9454 18470 9506 18522
rect 9518 18470 9570 18522
rect 9582 18470 9634 18522
rect 9646 18470 9698 18522
rect 17831 18470 17883 18522
rect 17895 18470 17947 18522
rect 17959 18470 18011 18522
rect 18023 18470 18075 18522
rect 18087 18470 18139 18522
rect 26272 18470 26324 18522
rect 26336 18470 26388 18522
rect 26400 18470 26452 18522
rect 26464 18470 26516 18522
rect 26528 18470 26580 18522
rect 34713 18470 34765 18522
rect 34777 18470 34829 18522
rect 34841 18470 34893 18522
rect 34905 18470 34957 18522
rect 34969 18470 35021 18522
rect 8944 18368 8996 18420
rect 12440 18368 12492 18420
rect 15752 18411 15804 18420
rect 7104 18300 7156 18352
rect 12072 18300 12124 18352
rect 12348 18300 12400 18352
rect 14740 18343 14792 18352
rect 6644 18232 6696 18284
rect 8116 18232 8168 18284
rect 11060 18232 11112 18284
rect 11796 18232 11848 18284
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 15752 18377 15761 18411
rect 15761 18377 15795 18411
rect 15795 18377 15804 18411
rect 15752 18368 15804 18377
rect 16672 18368 16724 18420
rect 24952 18368 25004 18420
rect 25688 18411 25740 18420
rect 25688 18377 25697 18411
rect 25697 18377 25731 18411
rect 25731 18377 25740 18411
rect 25688 18368 25740 18377
rect 16028 18300 16080 18352
rect 12992 18275 13044 18284
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 7288 18139 7340 18148
rect 7288 18105 7297 18139
rect 7297 18105 7331 18139
rect 7331 18105 7340 18139
rect 7288 18096 7340 18105
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 15660 18232 15712 18284
rect 18512 18300 18564 18352
rect 29092 18368 29144 18420
rect 24584 18232 24636 18284
rect 24860 18232 24912 18284
rect 25504 18275 25556 18284
rect 25504 18241 25513 18275
rect 25513 18241 25547 18275
rect 25547 18241 25556 18275
rect 25504 18232 25556 18241
rect 28356 18232 28408 18284
rect 31392 18300 31444 18352
rect 20352 18164 20404 18216
rect 23112 18164 23164 18216
rect 23848 18164 23900 18216
rect 12440 18096 12492 18148
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 18236 18028 18288 18080
rect 25320 18071 25372 18080
rect 25320 18037 25329 18071
rect 25329 18037 25363 18071
rect 25363 18037 25372 18071
rect 25320 18028 25372 18037
rect 27252 18164 27304 18216
rect 29000 18164 29052 18216
rect 29184 18232 29236 18284
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 30104 18164 30156 18216
rect 28540 18096 28592 18148
rect 32496 18368 32548 18420
rect 32680 18368 32732 18420
rect 32404 18232 32456 18284
rect 32312 18207 32364 18216
rect 32312 18173 32321 18207
rect 32321 18173 32355 18207
rect 32355 18173 32364 18207
rect 32312 18164 32364 18173
rect 32864 18207 32916 18216
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 34336 18207 34388 18216
rect 34336 18173 34345 18207
rect 34345 18173 34379 18207
rect 34379 18173 34388 18207
rect 34336 18164 34388 18173
rect 5170 17926 5222 17978
rect 5234 17926 5286 17978
rect 5298 17926 5350 17978
rect 5362 17926 5414 17978
rect 5426 17926 5478 17978
rect 13611 17926 13663 17978
rect 13675 17926 13727 17978
rect 13739 17926 13791 17978
rect 13803 17926 13855 17978
rect 13867 17926 13919 17978
rect 22052 17926 22104 17978
rect 22116 17926 22168 17978
rect 22180 17926 22232 17978
rect 22244 17926 22296 17978
rect 22308 17926 22360 17978
rect 30493 17926 30545 17978
rect 30557 17926 30609 17978
rect 30621 17926 30673 17978
rect 30685 17926 30737 17978
rect 30749 17926 30801 17978
rect 6736 17824 6788 17876
rect 15384 17824 15436 17876
rect 27988 17867 28040 17876
rect 3516 17756 3568 17808
rect 11520 17688 11572 17740
rect 3240 17663 3292 17672
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 15200 17663 15252 17672
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 17500 17620 17552 17672
rect 2688 17552 2740 17604
rect 12164 17552 12216 17604
rect 12900 17552 12952 17604
rect 17316 17552 17368 17604
rect 19248 17620 19300 17672
rect 27988 17833 27997 17867
rect 27997 17833 28031 17867
rect 28031 17833 28040 17867
rect 27988 17824 28040 17833
rect 29000 17824 29052 17876
rect 21548 17799 21600 17808
rect 21548 17765 21557 17799
rect 21557 17765 21591 17799
rect 21591 17765 21600 17799
rect 21548 17756 21600 17765
rect 24768 17756 24820 17808
rect 27896 17688 27948 17740
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 21548 17552 21600 17604
rect 25688 17620 25740 17672
rect 27712 17663 27764 17672
rect 27712 17629 27721 17663
rect 27721 17629 27755 17663
rect 27755 17629 27764 17663
rect 27712 17620 27764 17629
rect 27804 17663 27856 17672
rect 27804 17629 27813 17663
rect 27813 17629 27847 17663
rect 27847 17629 27856 17663
rect 27804 17620 27856 17629
rect 28540 17620 28592 17672
rect 28908 17663 28960 17672
rect 28908 17629 28917 17663
rect 28917 17629 28951 17663
rect 28951 17629 28960 17663
rect 28908 17620 28960 17629
rect 30932 17663 30984 17672
rect 30932 17629 30941 17663
rect 30941 17629 30975 17663
rect 30975 17629 30984 17663
rect 32312 17688 32364 17740
rect 30932 17620 30984 17629
rect 26608 17552 26660 17604
rect 31116 17595 31168 17604
rect 31116 17561 31125 17595
rect 31125 17561 31159 17595
rect 31159 17561 31168 17595
rect 31116 17552 31168 17561
rect 32772 17620 32824 17672
rect 3056 17527 3108 17536
rect 3056 17493 3065 17527
rect 3065 17493 3099 17527
rect 3099 17493 3108 17527
rect 3056 17484 3108 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 7104 17484 7156 17536
rect 9956 17484 10008 17536
rect 10968 17484 11020 17536
rect 12992 17484 13044 17536
rect 16580 17484 16632 17536
rect 17592 17484 17644 17536
rect 20904 17484 20956 17536
rect 24860 17484 24912 17536
rect 25780 17484 25832 17536
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 28816 17484 28868 17493
rect 33232 17484 33284 17536
rect 9390 17382 9442 17434
rect 9454 17382 9506 17434
rect 9518 17382 9570 17434
rect 9582 17382 9634 17434
rect 9646 17382 9698 17434
rect 17831 17382 17883 17434
rect 17895 17382 17947 17434
rect 17959 17382 18011 17434
rect 18023 17382 18075 17434
rect 18087 17382 18139 17434
rect 26272 17382 26324 17434
rect 26336 17382 26388 17434
rect 26400 17382 26452 17434
rect 26464 17382 26516 17434
rect 26528 17382 26580 17434
rect 34713 17382 34765 17434
rect 34777 17382 34829 17434
rect 34841 17382 34893 17434
rect 34905 17382 34957 17434
rect 34969 17382 35021 17434
rect 6920 17280 6972 17332
rect 2964 17255 3016 17264
rect 2964 17221 2973 17255
rect 2973 17221 3007 17255
rect 3007 17221 3016 17255
rect 2964 17212 3016 17221
rect 4252 17144 4304 17196
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 6828 17144 6880 17196
rect 7472 17144 7524 17196
rect 7748 17144 7800 17196
rect 9220 17212 9272 17264
rect 10324 17280 10376 17332
rect 14372 17280 14424 17332
rect 19432 17280 19484 17332
rect 12256 17212 12308 17264
rect 13176 17212 13228 17264
rect 16856 17255 16908 17264
rect 16856 17221 16865 17255
rect 16865 17221 16899 17255
rect 16899 17221 16908 17255
rect 16856 17212 16908 17221
rect 18236 17255 18288 17264
rect 18236 17221 18245 17255
rect 18245 17221 18279 17255
rect 18279 17221 18288 17255
rect 18236 17212 18288 17221
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 10048 17144 10100 17196
rect 15384 17144 15436 17196
rect 17224 17144 17276 17196
rect 21180 17212 21232 17264
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 6644 17119 6696 17128
rect 6644 17085 6653 17119
rect 6653 17085 6687 17119
rect 6687 17085 6696 17119
rect 6644 17076 6696 17085
rect 10140 17076 10192 17128
rect 11520 17076 11572 17128
rect 15936 17119 15988 17128
rect 15936 17085 15945 17119
rect 15945 17085 15979 17119
rect 15979 17085 15988 17119
rect 15936 17076 15988 17085
rect 17500 17076 17552 17128
rect 20996 17144 21048 17196
rect 23204 17280 23256 17332
rect 25688 17323 25740 17332
rect 23572 17212 23624 17264
rect 23848 17144 23900 17196
rect 25044 17187 25096 17196
rect 25044 17153 25053 17187
rect 25053 17153 25087 17187
rect 25087 17153 25096 17187
rect 25044 17144 25096 17153
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 27804 17280 27856 17332
rect 28816 17280 28868 17332
rect 29092 17280 29144 17332
rect 30932 17323 30984 17332
rect 30932 17289 30941 17323
rect 30941 17289 30975 17323
rect 30975 17289 30984 17323
rect 30932 17280 30984 17289
rect 25780 17212 25832 17264
rect 32220 17280 32272 17332
rect 32864 17280 32916 17332
rect 33232 17323 33284 17332
rect 33232 17289 33241 17323
rect 33241 17289 33275 17323
rect 33275 17289 33284 17323
rect 33232 17280 33284 17289
rect 22560 17076 22612 17128
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 8116 17008 8168 17060
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 11152 16940 11204 16992
rect 19248 17008 19300 17060
rect 19524 17008 19576 17060
rect 25596 17144 25648 17196
rect 26056 17144 26108 17196
rect 28540 17187 28592 17196
rect 28540 17153 28549 17187
rect 28549 17153 28583 17187
rect 28583 17153 28592 17187
rect 28540 17144 28592 17153
rect 28908 17144 28960 17196
rect 26608 17076 26660 17128
rect 30288 17076 30340 17128
rect 31392 17144 31444 17196
rect 31576 17144 31628 17196
rect 32404 17144 32456 17196
rect 32772 17144 32824 17196
rect 12624 16940 12676 16992
rect 20444 16983 20496 16992
rect 20444 16949 20453 16983
rect 20453 16949 20487 16983
rect 20487 16949 20496 16983
rect 20444 16940 20496 16949
rect 23388 16940 23440 16992
rect 24400 16940 24452 16992
rect 24768 16940 24820 16992
rect 31300 16940 31352 16992
rect 32772 16940 32824 16992
rect 5170 16838 5222 16890
rect 5234 16838 5286 16890
rect 5298 16838 5350 16890
rect 5362 16838 5414 16890
rect 5426 16838 5478 16890
rect 13611 16838 13663 16890
rect 13675 16838 13727 16890
rect 13739 16838 13791 16890
rect 13803 16838 13855 16890
rect 13867 16838 13919 16890
rect 22052 16838 22104 16890
rect 22116 16838 22168 16890
rect 22180 16838 22232 16890
rect 22244 16838 22296 16890
rect 22308 16838 22360 16890
rect 30493 16838 30545 16890
rect 30557 16838 30609 16890
rect 30621 16838 30673 16890
rect 30685 16838 30737 16890
rect 30749 16838 30801 16890
rect 2688 16736 2740 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 6552 16736 6604 16788
rect 6644 16668 6696 16720
rect 11060 16736 11112 16788
rect 12256 16779 12308 16788
rect 12256 16745 12265 16779
rect 12265 16745 12299 16779
rect 12299 16745 12308 16779
rect 12256 16736 12308 16745
rect 15476 16736 15528 16788
rect 15936 16736 15988 16788
rect 19432 16736 19484 16788
rect 7196 16711 7248 16720
rect 7196 16677 7205 16711
rect 7205 16677 7239 16711
rect 7239 16677 7248 16711
rect 7196 16668 7248 16677
rect 8208 16668 8260 16720
rect 7288 16643 7340 16652
rect 4252 16575 4304 16584
rect 3056 16464 3108 16516
rect 4252 16541 4261 16575
rect 4261 16541 4295 16575
rect 4295 16541 4304 16575
rect 4252 16532 4304 16541
rect 6460 16532 6512 16584
rect 7288 16609 7334 16643
rect 7334 16609 7340 16643
rect 10968 16668 11020 16720
rect 15200 16668 15252 16720
rect 20996 16736 21048 16788
rect 26148 16736 26200 16788
rect 31116 16736 31168 16788
rect 31300 16736 31352 16788
rect 32220 16779 32272 16788
rect 7288 16600 7340 16609
rect 12440 16600 12492 16652
rect 14740 16600 14792 16652
rect 17500 16643 17552 16652
rect 17500 16609 17509 16643
rect 17509 16609 17543 16643
rect 17543 16609 17552 16643
rect 17500 16600 17552 16609
rect 26056 16600 26108 16652
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 11060 16532 11112 16584
rect 12072 16532 12124 16584
rect 5080 16464 5132 16516
rect 6368 16396 6420 16448
rect 6552 16396 6604 16448
rect 11152 16464 11204 16516
rect 14280 16464 14332 16516
rect 15384 16532 15436 16584
rect 16580 16532 16632 16584
rect 17224 16575 17276 16584
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 19524 16532 19576 16584
rect 20444 16532 20496 16584
rect 24584 16575 24636 16584
rect 17316 16464 17368 16516
rect 19248 16464 19300 16516
rect 24584 16541 24593 16575
rect 24593 16541 24627 16575
rect 24627 16541 24636 16575
rect 24584 16532 24636 16541
rect 22468 16464 22520 16516
rect 29000 16600 29052 16652
rect 29736 16643 29788 16652
rect 29736 16609 29745 16643
rect 29745 16609 29779 16643
rect 29779 16609 29788 16643
rect 29736 16600 29788 16609
rect 26056 16464 26108 16516
rect 26700 16507 26752 16516
rect 26700 16473 26709 16507
rect 26709 16473 26743 16507
rect 26743 16473 26752 16507
rect 26700 16464 26752 16473
rect 29092 16464 29144 16516
rect 31392 16600 31444 16652
rect 31576 16668 31628 16720
rect 32220 16745 32229 16779
rect 32229 16745 32263 16779
rect 32263 16745 32272 16779
rect 32220 16736 32272 16745
rect 33692 16668 33744 16720
rect 32588 16643 32640 16652
rect 32588 16609 32597 16643
rect 32597 16609 32631 16643
rect 32631 16609 32640 16643
rect 32588 16600 32640 16609
rect 32036 16532 32088 16584
rect 10416 16396 10468 16448
rect 14464 16439 14516 16448
rect 14464 16405 14473 16439
rect 14473 16405 14507 16439
rect 14507 16405 14516 16439
rect 14464 16396 14516 16405
rect 17592 16396 17644 16448
rect 21180 16396 21232 16448
rect 25964 16439 26016 16448
rect 25964 16405 25973 16439
rect 25973 16405 26007 16439
rect 26007 16405 26016 16439
rect 25964 16396 26016 16405
rect 30104 16439 30156 16448
rect 30104 16405 30113 16439
rect 30113 16405 30147 16439
rect 30147 16405 30156 16439
rect 30288 16439 30340 16448
rect 30104 16396 30156 16405
rect 30288 16405 30297 16439
rect 30297 16405 30331 16439
rect 30331 16405 30340 16439
rect 30288 16396 30340 16405
rect 9390 16294 9442 16346
rect 9454 16294 9506 16346
rect 9518 16294 9570 16346
rect 9582 16294 9634 16346
rect 9646 16294 9698 16346
rect 17831 16294 17883 16346
rect 17895 16294 17947 16346
rect 17959 16294 18011 16346
rect 18023 16294 18075 16346
rect 18087 16294 18139 16346
rect 26272 16294 26324 16346
rect 26336 16294 26388 16346
rect 26400 16294 26452 16346
rect 26464 16294 26516 16346
rect 26528 16294 26580 16346
rect 34713 16294 34765 16346
rect 34777 16294 34829 16346
rect 34841 16294 34893 16346
rect 34905 16294 34957 16346
rect 34969 16294 35021 16346
rect 5540 16192 5592 16244
rect 6460 16192 6512 16244
rect 6736 16235 6788 16244
rect 6736 16201 6745 16235
rect 6745 16201 6779 16235
rect 6779 16201 6788 16235
rect 6736 16192 6788 16201
rect 12256 16192 12308 16244
rect 13360 16192 13412 16244
rect 5724 16167 5776 16176
rect 5724 16133 5733 16167
rect 5733 16133 5767 16167
rect 5767 16133 5776 16167
rect 5724 16124 5776 16133
rect 6828 16124 6880 16176
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6644 16056 6696 16108
rect 7288 16124 7340 16176
rect 11520 16124 11572 16176
rect 7196 16056 7248 16108
rect 7472 16056 7524 16108
rect 10416 16099 10468 16108
rect 10416 16065 10425 16099
rect 10425 16065 10459 16099
rect 10459 16065 10468 16099
rect 10416 16056 10468 16065
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 7104 15988 7156 16040
rect 6460 15920 6512 15972
rect 19248 16192 19300 16244
rect 19524 16235 19576 16244
rect 19524 16201 19533 16235
rect 19533 16201 19567 16235
rect 19567 16201 19576 16235
rect 19524 16192 19576 16201
rect 20536 16192 20588 16244
rect 22652 16235 22704 16244
rect 14280 16167 14332 16176
rect 14280 16133 14289 16167
rect 14289 16133 14323 16167
rect 14323 16133 14332 16167
rect 14280 16124 14332 16133
rect 15200 16167 15252 16176
rect 15200 16133 15234 16167
rect 15234 16133 15252 16167
rect 15200 16124 15252 16133
rect 18236 16167 18288 16176
rect 18236 16133 18245 16167
rect 18245 16133 18279 16167
rect 18279 16133 18288 16167
rect 18236 16124 18288 16133
rect 21180 16124 21232 16176
rect 22652 16201 22661 16235
rect 22661 16201 22695 16235
rect 22695 16201 22704 16235
rect 22652 16192 22704 16201
rect 26056 16235 26108 16244
rect 26056 16201 26065 16235
rect 26065 16201 26099 16235
rect 26099 16201 26108 16235
rect 26056 16192 26108 16201
rect 17408 16099 17460 16108
rect 17408 16065 17417 16099
rect 17417 16065 17451 16099
rect 17451 16065 17460 16099
rect 17408 16056 17460 16065
rect 17684 16099 17736 16108
rect 17684 16065 17693 16099
rect 17693 16065 17727 16099
rect 17727 16065 17736 16099
rect 17684 16056 17736 16065
rect 20536 16056 20588 16108
rect 14740 15988 14792 16040
rect 19616 15988 19668 16040
rect 20904 16099 20956 16108
rect 20904 16065 20949 16099
rect 20949 16065 20956 16099
rect 21088 16099 21140 16108
rect 20904 16056 20956 16065
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 21916 16056 21968 16108
rect 25964 16124 26016 16176
rect 23112 16056 23164 16108
rect 25136 16099 25188 16108
rect 25136 16065 25145 16099
rect 25145 16065 25179 16099
rect 25179 16065 25188 16099
rect 25136 16056 25188 16065
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 26608 16056 26660 16108
rect 27712 16056 27764 16108
rect 29092 16192 29144 16244
rect 32588 16192 32640 16244
rect 33048 16192 33100 16244
rect 31392 16124 31444 16176
rect 33232 16124 33284 16176
rect 24400 15988 24452 16040
rect 29000 16056 29052 16108
rect 30288 16056 30340 16108
rect 33876 16056 33928 16108
rect 30104 15988 30156 16040
rect 32312 16031 32364 16040
rect 32312 15997 32321 16031
rect 32321 15997 32355 16031
rect 32355 15997 32364 16031
rect 32312 15988 32364 15997
rect 32220 15920 32272 15972
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 14464 15852 14516 15904
rect 20076 15852 20128 15904
rect 24584 15852 24636 15904
rect 28172 15852 28224 15904
rect 29460 15895 29512 15904
rect 29460 15861 29469 15895
rect 29469 15861 29503 15895
rect 29503 15861 29512 15895
rect 29460 15852 29512 15861
rect 5170 15750 5222 15802
rect 5234 15750 5286 15802
rect 5298 15750 5350 15802
rect 5362 15750 5414 15802
rect 5426 15750 5478 15802
rect 13611 15750 13663 15802
rect 13675 15750 13727 15802
rect 13739 15750 13791 15802
rect 13803 15750 13855 15802
rect 13867 15750 13919 15802
rect 22052 15750 22104 15802
rect 22116 15750 22168 15802
rect 22180 15750 22232 15802
rect 22244 15750 22296 15802
rect 22308 15750 22360 15802
rect 30493 15750 30545 15802
rect 30557 15750 30609 15802
rect 30621 15750 30673 15802
rect 30685 15750 30737 15802
rect 30749 15750 30801 15802
rect 4988 15648 5040 15700
rect 7748 15648 7800 15700
rect 11060 15648 11112 15700
rect 2964 15580 3016 15632
rect 14556 15580 14608 15632
rect 5080 15512 5132 15564
rect 6552 15512 6604 15564
rect 13452 15512 13504 15564
rect 4252 15444 4304 15496
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6460 15444 6512 15496
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 12624 15487 12676 15496
rect 12624 15453 12633 15487
rect 12633 15453 12667 15487
rect 12667 15453 12676 15487
rect 12624 15444 12676 15453
rect 14280 15444 14332 15496
rect 15660 15444 15712 15496
rect 16580 15580 16632 15632
rect 17408 15580 17460 15632
rect 16396 15512 16448 15564
rect 16212 15444 16264 15496
rect 25136 15648 25188 15700
rect 26056 15648 26108 15700
rect 31760 15648 31812 15700
rect 32312 15648 32364 15700
rect 33876 15691 33928 15700
rect 33876 15657 33885 15691
rect 33885 15657 33919 15691
rect 33919 15657 33928 15691
rect 33876 15648 33928 15657
rect 21916 15580 21968 15632
rect 19984 15512 20036 15564
rect 22560 15555 22612 15564
rect 22560 15521 22569 15555
rect 22569 15521 22603 15555
rect 22603 15521 22612 15555
rect 22560 15512 22612 15521
rect 18328 15444 18380 15496
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 24768 15512 24820 15564
rect 28172 15555 28224 15564
rect 28172 15521 28181 15555
rect 28181 15521 28215 15555
rect 28215 15521 28224 15555
rect 28172 15512 28224 15521
rect 29460 15512 29512 15564
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 27804 15444 27856 15496
rect 28448 15487 28500 15496
rect 28448 15453 28457 15487
rect 28457 15453 28491 15487
rect 28491 15453 28500 15487
rect 28448 15444 28500 15453
rect 33416 15487 33468 15496
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 33692 15487 33744 15496
rect 33692 15453 33701 15487
rect 33701 15453 33735 15487
rect 33735 15453 33744 15487
rect 33692 15444 33744 15453
rect 5540 15376 5592 15428
rect 4436 15308 4488 15360
rect 7196 15376 7248 15428
rect 12072 15376 12124 15428
rect 17316 15376 17368 15428
rect 17684 15419 17736 15428
rect 17684 15385 17693 15419
rect 17693 15385 17727 15419
rect 17727 15385 17736 15419
rect 17684 15376 17736 15385
rect 22376 15376 22428 15428
rect 23388 15419 23440 15428
rect 23388 15385 23397 15419
rect 23397 15385 23431 15419
rect 23431 15385 23440 15419
rect 23388 15376 23440 15385
rect 25136 15419 25188 15428
rect 25136 15385 25145 15419
rect 25145 15385 25179 15419
rect 25179 15385 25188 15419
rect 25136 15376 25188 15385
rect 33600 15376 33652 15428
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 20996 15308 21048 15360
rect 33048 15308 33100 15360
rect 9390 15206 9442 15258
rect 9454 15206 9506 15258
rect 9518 15206 9570 15258
rect 9582 15206 9634 15258
rect 9646 15206 9698 15258
rect 17831 15206 17883 15258
rect 17895 15206 17947 15258
rect 17959 15206 18011 15258
rect 18023 15206 18075 15258
rect 18087 15206 18139 15258
rect 26272 15206 26324 15258
rect 26336 15206 26388 15258
rect 26400 15206 26452 15258
rect 26464 15206 26516 15258
rect 26528 15206 26580 15258
rect 34713 15206 34765 15258
rect 34777 15206 34829 15258
rect 34841 15206 34893 15258
rect 34905 15206 34957 15258
rect 34969 15206 35021 15258
rect 5724 15104 5776 15156
rect 6368 15104 6420 15156
rect 18420 15104 18472 15156
rect 2964 15036 3016 15088
rect 6460 15036 6512 15088
rect 11980 15036 12032 15088
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 2688 14900 2740 14952
rect 3240 14832 3292 14884
rect 4528 14968 4580 15020
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 9036 14968 9088 14977
rect 9772 14968 9824 15020
rect 10324 14968 10376 15020
rect 10692 15011 10744 15020
rect 8944 14943 8996 14952
rect 8944 14909 8953 14943
rect 8953 14909 8987 14943
rect 8987 14909 8996 14943
rect 8944 14900 8996 14909
rect 9864 14900 9916 14952
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 12164 14968 12216 15020
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 13452 14968 13504 15020
rect 15660 14968 15712 15020
rect 16212 14968 16264 15020
rect 21824 15104 21876 15156
rect 22284 15147 22336 15156
rect 22284 15113 22293 15147
rect 22293 15113 22327 15147
rect 22327 15113 22336 15147
rect 22284 15104 22336 15113
rect 23388 15104 23440 15156
rect 25136 15104 25188 15156
rect 33600 15147 33652 15156
rect 33600 15113 33609 15147
rect 33609 15113 33643 15147
rect 33643 15113 33652 15147
rect 33600 15104 33652 15113
rect 19340 15036 19392 15088
rect 21916 15036 21968 15088
rect 26700 15036 26752 15088
rect 18236 15011 18288 15020
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 20352 14968 20404 15020
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 22468 14968 22520 15020
rect 23388 14968 23440 15020
rect 25136 15011 25188 15020
rect 25136 14977 25154 15011
rect 25154 14977 25188 15011
rect 25136 14968 25188 14977
rect 29920 14968 29972 15020
rect 18144 14900 18196 14952
rect 26424 14900 26476 14952
rect 16856 14832 16908 14884
rect 19616 14832 19668 14884
rect 22468 14832 22520 14884
rect 23204 14832 23256 14884
rect 29644 14875 29696 14884
rect 29644 14841 29653 14875
rect 29653 14841 29687 14875
rect 29687 14841 29696 14875
rect 29644 14832 29696 14841
rect 4252 14764 4304 14816
rect 6092 14764 6144 14816
rect 19708 14807 19760 14816
rect 19708 14773 19717 14807
rect 19717 14773 19751 14807
rect 19751 14773 19760 14807
rect 19708 14764 19760 14773
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 20904 14764 20956 14816
rect 22284 14764 22336 14816
rect 23296 14807 23348 14816
rect 23296 14773 23305 14807
rect 23305 14773 23339 14807
rect 23339 14773 23348 14807
rect 23296 14764 23348 14773
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 5170 14662 5222 14714
rect 5234 14662 5286 14714
rect 5298 14662 5350 14714
rect 5362 14662 5414 14714
rect 5426 14662 5478 14714
rect 13611 14662 13663 14714
rect 13675 14662 13727 14714
rect 13739 14662 13791 14714
rect 13803 14662 13855 14714
rect 13867 14662 13919 14714
rect 22052 14662 22104 14714
rect 22116 14662 22168 14714
rect 22180 14662 22232 14714
rect 22244 14662 22296 14714
rect 22308 14662 22360 14714
rect 30493 14662 30545 14714
rect 30557 14662 30609 14714
rect 30621 14662 30673 14714
rect 30685 14662 30737 14714
rect 30749 14662 30801 14714
rect 6828 14560 6880 14612
rect 7196 14603 7248 14612
rect 7196 14569 7205 14603
rect 7205 14569 7239 14603
rect 7239 14569 7248 14603
rect 7196 14560 7248 14569
rect 19432 14560 19484 14612
rect 8300 14492 8352 14544
rect 8484 14535 8536 14544
rect 8484 14501 8493 14535
rect 8493 14501 8527 14535
rect 8527 14501 8536 14535
rect 8484 14492 8536 14501
rect 9312 14492 9364 14544
rect 20720 14492 20772 14544
rect 22376 14560 22428 14612
rect 25780 14560 25832 14612
rect 26608 14560 26660 14612
rect 33232 14603 33284 14612
rect 23296 14492 23348 14544
rect 1400 14424 1452 14476
rect 17316 14467 17368 14476
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 3056 14356 3108 14408
rect 6368 14399 6420 14408
rect 2964 14331 3016 14340
rect 2964 14297 2973 14331
rect 2973 14297 3007 14331
rect 3007 14297 3016 14331
rect 2964 14288 3016 14297
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 7196 14356 7248 14408
rect 7932 14399 7984 14408
rect 7932 14365 7941 14399
rect 7941 14365 7975 14399
rect 7975 14365 7984 14399
rect 7932 14356 7984 14365
rect 11060 14356 11112 14408
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 6644 14288 6696 14340
rect 7840 14288 7892 14340
rect 8208 14331 8260 14340
rect 8208 14297 8217 14331
rect 8217 14297 8251 14331
rect 8251 14297 8260 14331
rect 8208 14288 8260 14297
rect 9772 14331 9824 14340
rect 6920 14220 6972 14272
rect 7472 14220 7524 14272
rect 8116 14220 8168 14272
rect 9772 14297 9781 14331
rect 9781 14297 9815 14331
rect 9815 14297 9824 14331
rect 9772 14288 9824 14297
rect 10692 14288 10744 14340
rect 12440 14288 12492 14340
rect 13728 14356 13780 14408
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 24584 14467 24636 14476
rect 17316 14424 17368 14433
rect 24584 14433 24593 14467
rect 24593 14433 24627 14467
rect 24627 14433 24636 14467
rect 24584 14424 24636 14433
rect 17684 14356 17736 14408
rect 18144 14356 18196 14408
rect 18420 14356 18472 14408
rect 13084 14331 13136 14340
rect 13084 14297 13093 14331
rect 13093 14297 13127 14331
rect 13127 14297 13136 14331
rect 13084 14288 13136 14297
rect 19340 14288 19392 14340
rect 19708 14356 19760 14408
rect 20996 14399 21048 14408
rect 20996 14365 21030 14399
rect 21030 14365 21048 14399
rect 20996 14356 21048 14365
rect 24860 14399 24912 14408
rect 24860 14365 24894 14399
rect 24894 14365 24912 14399
rect 24860 14356 24912 14365
rect 26424 14399 26476 14408
rect 26424 14365 26433 14399
rect 26433 14365 26467 14399
rect 26467 14365 26476 14399
rect 26424 14356 26476 14365
rect 26976 14356 27028 14408
rect 33232 14569 33241 14603
rect 33241 14569 33275 14603
rect 33275 14569 33284 14603
rect 33232 14560 33284 14569
rect 31760 14424 31812 14476
rect 32312 14424 32364 14476
rect 28816 14356 28868 14408
rect 30104 14356 30156 14408
rect 32128 14399 32180 14408
rect 32128 14365 32137 14399
rect 32137 14365 32171 14399
rect 32171 14365 32180 14399
rect 32128 14356 32180 14365
rect 22100 14288 22152 14340
rect 22192 14288 22244 14340
rect 23388 14288 23440 14340
rect 10232 14220 10284 14272
rect 19616 14263 19668 14272
rect 19616 14229 19625 14263
rect 19625 14229 19659 14263
rect 19659 14229 19668 14263
rect 19616 14220 19668 14229
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 21180 14220 21232 14272
rect 24768 14220 24820 14272
rect 29000 14288 29052 14340
rect 25596 14220 25648 14272
rect 27528 14220 27580 14272
rect 27620 14220 27672 14272
rect 31944 14220 31996 14272
rect 32772 14220 32824 14272
rect 9390 14118 9442 14170
rect 9454 14118 9506 14170
rect 9518 14118 9570 14170
rect 9582 14118 9634 14170
rect 9646 14118 9698 14170
rect 17831 14118 17883 14170
rect 17895 14118 17947 14170
rect 17959 14118 18011 14170
rect 18023 14118 18075 14170
rect 18087 14118 18139 14170
rect 26272 14118 26324 14170
rect 26336 14118 26388 14170
rect 26400 14118 26452 14170
rect 26464 14118 26516 14170
rect 26528 14118 26580 14170
rect 34713 14118 34765 14170
rect 34777 14118 34829 14170
rect 34841 14118 34893 14170
rect 34905 14118 34957 14170
rect 34969 14118 35021 14170
rect 1676 14016 1728 14068
rect 2964 14016 3016 14068
rect 3700 14016 3752 14068
rect 4436 13991 4488 14000
rect 4436 13957 4445 13991
rect 4445 13957 4479 13991
rect 4479 13957 4488 13991
rect 4436 13948 4488 13957
rect 3056 13880 3108 13932
rect 3608 13880 3660 13932
rect 5540 13880 5592 13932
rect 7932 14016 7984 14068
rect 8208 14016 8260 14068
rect 9956 14016 10008 14068
rect 6368 13948 6420 14000
rect 6644 13948 6696 14000
rect 7472 13948 7524 14000
rect 8392 13880 8444 13932
rect 11060 13948 11112 14000
rect 4160 13855 4212 13864
rect 4160 13821 4169 13855
rect 4169 13821 4203 13855
rect 4203 13821 4212 13855
rect 4160 13812 4212 13821
rect 5080 13812 5132 13864
rect 12440 14016 12492 14068
rect 12808 14016 12860 14068
rect 11980 13948 12032 14000
rect 13084 13948 13136 14000
rect 13728 13880 13780 13932
rect 16948 14016 17000 14068
rect 20168 14016 20220 14068
rect 20628 14016 20680 14068
rect 19432 13948 19484 14000
rect 20444 13948 20496 14000
rect 24032 13948 24084 14000
rect 24768 13948 24820 14000
rect 29000 14016 29052 14068
rect 29920 14016 29972 14068
rect 30104 14059 30156 14068
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 31944 14016 31996 14068
rect 32036 14016 32088 14068
rect 33692 14016 33744 14068
rect 28724 13991 28776 14000
rect 28724 13957 28733 13991
rect 28733 13957 28767 13991
rect 28767 13957 28776 13991
rect 28724 13948 28776 13957
rect 28908 13991 28960 14000
rect 28908 13957 28917 13991
rect 28917 13957 28951 13991
rect 28951 13957 28960 13991
rect 28908 13948 28960 13957
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 16856 13923 16908 13932
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 13268 13812 13320 13864
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 15200 13812 15252 13864
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 17684 13880 17736 13932
rect 18788 13923 18840 13932
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 22468 13880 22520 13932
rect 24584 13923 24636 13932
rect 20812 13812 20864 13864
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 25044 13880 25096 13932
rect 27712 13923 27764 13932
rect 26608 13812 26660 13864
rect 27344 13855 27396 13864
rect 27344 13821 27353 13855
rect 27353 13821 27387 13855
rect 27387 13821 27396 13855
rect 27344 13812 27396 13821
rect 27712 13889 27721 13923
rect 27721 13889 27755 13923
rect 27755 13889 27764 13923
rect 27712 13880 27764 13889
rect 27804 13923 27856 13932
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 29644 13923 29696 13932
rect 27804 13880 27856 13889
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 30380 13880 30432 13932
rect 25136 13744 25188 13796
rect 6828 13676 6880 13728
rect 28632 13812 28684 13864
rect 28908 13719 28960 13728
rect 28908 13685 28917 13719
rect 28917 13685 28951 13719
rect 28951 13685 28960 13719
rect 28908 13676 28960 13685
rect 29644 13676 29696 13728
rect 32036 13812 32088 13864
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 32772 13812 32824 13864
rect 33416 13676 33468 13728
rect 5170 13574 5222 13626
rect 5234 13574 5286 13626
rect 5298 13574 5350 13626
rect 5362 13574 5414 13626
rect 5426 13574 5478 13626
rect 13611 13574 13663 13626
rect 13675 13574 13727 13626
rect 13739 13574 13791 13626
rect 13803 13574 13855 13626
rect 13867 13574 13919 13626
rect 22052 13574 22104 13626
rect 22116 13574 22168 13626
rect 22180 13574 22232 13626
rect 22244 13574 22296 13626
rect 22308 13574 22360 13626
rect 30493 13574 30545 13626
rect 30557 13574 30609 13626
rect 30621 13574 30673 13626
rect 30685 13574 30737 13626
rect 30749 13574 30801 13626
rect 4160 13472 4212 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 4252 13404 4304 13456
rect 10508 13472 10560 13524
rect 3884 13268 3936 13320
rect 8300 13404 8352 13456
rect 9128 13379 9180 13388
rect 5080 13268 5132 13320
rect 3976 13200 4028 13252
rect 4068 13200 4120 13252
rect 8300 13311 8352 13320
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 3148 13132 3200 13184
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 8668 13200 8720 13252
rect 7472 13132 7524 13184
rect 8484 13132 8536 13184
rect 9864 13200 9916 13252
rect 9036 13132 9088 13184
rect 15384 13472 15436 13524
rect 15660 13515 15712 13524
rect 11152 13336 11204 13388
rect 11520 13336 11572 13388
rect 13084 13336 13136 13388
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 15660 13481 15669 13515
rect 15669 13481 15703 13515
rect 15703 13481 15712 13515
rect 15660 13472 15712 13481
rect 26976 13472 27028 13524
rect 32312 13472 32364 13524
rect 18328 13404 18380 13456
rect 15752 13268 15804 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 14096 13200 14148 13252
rect 15568 13200 15620 13252
rect 16856 13200 16908 13252
rect 17500 13200 17552 13252
rect 20536 13336 20588 13388
rect 22376 13336 22428 13388
rect 19800 13268 19852 13320
rect 26056 13311 26108 13320
rect 26056 13277 26065 13311
rect 26065 13277 26099 13311
rect 26099 13277 26108 13311
rect 26056 13268 26108 13277
rect 33600 13268 33652 13320
rect 18512 13200 18564 13252
rect 18236 13132 18288 13184
rect 9390 13030 9442 13082
rect 9454 13030 9506 13082
rect 9518 13030 9570 13082
rect 9582 13030 9634 13082
rect 9646 13030 9698 13082
rect 17831 13030 17883 13082
rect 17895 13030 17947 13082
rect 17959 13030 18011 13082
rect 18023 13030 18075 13082
rect 18087 13030 18139 13082
rect 26272 13030 26324 13082
rect 26336 13030 26388 13082
rect 26400 13030 26452 13082
rect 26464 13030 26516 13082
rect 26528 13030 26580 13082
rect 34713 13030 34765 13082
rect 34777 13030 34829 13082
rect 34841 13030 34893 13082
rect 34905 13030 34957 13082
rect 34969 13030 35021 13082
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 3976 12928 4028 12980
rect 9128 12928 9180 12980
rect 2412 12903 2464 12912
rect 2412 12869 2421 12903
rect 2421 12869 2455 12903
rect 2455 12869 2464 12903
rect 2412 12860 2464 12869
rect 3056 12860 3108 12912
rect 8668 12860 8720 12912
rect 9312 12860 9364 12912
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 11796 12928 11848 12980
rect 17592 12928 17644 12980
rect 22928 12971 22980 12980
rect 12992 12903 13044 12912
rect 12992 12869 13001 12903
rect 13001 12869 13035 12903
rect 13035 12869 13044 12903
rect 12992 12860 13044 12869
rect 14740 12903 14792 12912
rect 14740 12869 14749 12903
rect 14749 12869 14783 12903
rect 14783 12869 14792 12903
rect 14740 12860 14792 12869
rect 18328 12860 18380 12912
rect 15200 12792 15252 12844
rect 15568 12792 15620 12844
rect 3148 12724 3200 12776
rect 3608 12724 3660 12776
rect 16396 12792 16448 12844
rect 18052 12835 18104 12844
rect 10508 12656 10560 12708
rect 13176 12656 13228 12708
rect 16580 12724 16632 12776
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18420 12792 18472 12844
rect 18696 12792 18748 12844
rect 19616 12860 19668 12912
rect 19800 12792 19852 12844
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 28448 12928 28500 12980
rect 28540 12928 28592 12980
rect 32128 12928 32180 12980
rect 33232 12928 33284 12980
rect 24768 12860 24820 12912
rect 27528 12903 27580 12912
rect 27528 12869 27537 12903
rect 27537 12869 27571 12903
rect 27571 12869 27580 12903
rect 27528 12860 27580 12869
rect 28264 12860 28316 12912
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 22928 12792 22980 12844
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 27988 12792 28040 12844
rect 30288 12860 30340 12912
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 7564 12588 7616 12640
rect 14556 12588 14608 12640
rect 21088 12724 21140 12776
rect 23020 12724 23072 12776
rect 27620 12724 27672 12776
rect 29644 12792 29696 12844
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 33416 12792 33468 12844
rect 30196 12724 30248 12776
rect 19984 12588 20036 12640
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 23296 12656 23348 12708
rect 28080 12656 28132 12708
rect 28908 12656 28960 12708
rect 31024 12656 31076 12708
rect 28356 12631 28408 12640
rect 21088 12588 21140 12597
rect 28356 12597 28365 12631
rect 28365 12597 28399 12631
rect 28399 12597 28408 12631
rect 28356 12588 28408 12597
rect 5170 12486 5222 12538
rect 5234 12486 5286 12538
rect 5298 12486 5350 12538
rect 5362 12486 5414 12538
rect 5426 12486 5478 12538
rect 13611 12486 13663 12538
rect 13675 12486 13727 12538
rect 13739 12486 13791 12538
rect 13803 12486 13855 12538
rect 13867 12486 13919 12538
rect 22052 12486 22104 12538
rect 22116 12486 22168 12538
rect 22180 12486 22232 12538
rect 22244 12486 22296 12538
rect 22308 12486 22360 12538
rect 30493 12486 30545 12538
rect 30557 12486 30609 12538
rect 30621 12486 30673 12538
rect 30685 12486 30737 12538
rect 30749 12486 30801 12538
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 19800 12384 19852 12436
rect 20260 12384 20312 12436
rect 20812 12384 20864 12436
rect 21916 12384 21968 12436
rect 22744 12384 22796 12436
rect 23020 12427 23072 12436
rect 23020 12393 23029 12427
rect 23029 12393 23063 12427
rect 23063 12393 23072 12427
rect 23020 12384 23072 12393
rect 23388 12384 23440 12436
rect 24860 12384 24912 12436
rect 18328 12316 18380 12368
rect 23112 12316 23164 12368
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 2964 12112 3016 12164
rect 4068 12180 4120 12232
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 15752 12180 15804 12232
rect 16488 12180 16540 12232
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 18052 12248 18104 12300
rect 18788 12180 18840 12232
rect 21088 12248 21140 12300
rect 16948 12112 17000 12164
rect 18696 12112 18748 12164
rect 19616 12180 19668 12232
rect 20352 12180 20404 12232
rect 20536 12180 20588 12232
rect 22468 12180 22520 12232
rect 23296 12223 23348 12232
rect 23296 12189 23305 12223
rect 23305 12189 23339 12223
rect 23339 12189 23348 12223
rect 24676 12248 24728 12300
rect 23296 12180 23348 12189
rect 20260 12112 20312 12164
rect 20720 12112 20772 12164
rect 21272 12112 21324 12164
rect 22100 12112 22152 12164
rect 22192 12112 22244 12164
rect 22928 12112 22980 12164
rect 24860 12180 24912 12232
rect 28816 12316 28868 12368
rect 32128 12316 32180 12368
rect 27804 12180 27856 12232
rect 28540 12223 28592 12232
rect 28540 12189 28548 12223
rect 28548 12189 28582 12223
rect 28582 12189 28592 12223
rect 28540 12180 28592 12189
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 20168 12044 20220 12096
rect 22652 12044 22704 12096
rect 24584 12087 24636 12096
rect 24584 12053 24593 12087
rect 24593 12053 24627 12087
rect 24627 12053 24636 12087
rect 24584 12044 24636 12053
rect 24768 12044 24820 12096
rect 28448 12112 28500 12164
rect 31208 12044 31260 12096
rect 9390 11942 9442 11994
rect 9454 11942 9506 11994
rect 9518 11942 9570 11994
rect 9582 11942 9634 11994
rect 9646 11942 9698 11994
rect 17831 11942 17883 11994
rect 17895 11942 17947 11994
rect 17959 11942 18011 11994
rect 18023 11942 18075 11994
rect 18087 11942 18139 11994
rect 26272 11942 26324 11994
rect 26336 11942 26388 11994
rect 26400 11942 26452 11994
rect 26464 11942 26516 11994
rect 26528 11942 26580 11994
rect 34713 11942 34765 11994
rect 34777 11942 34829 11994
rect 34841 11942 34893 11994
rect 34905 11942 34957 11994
rect 34969 11942 35021 11994
rect 22192 11840 22244 11892
rect 22376 11883 22428 11892
rect 22376 11849 22385 11883
rect 22385 11849 22419 11883
rect 22419 11849 22428 11883
rect 22376 11840 22428 11849
rect 22836 11840 22888 11892
rect 13268 11704 13320 11756
rect 15200 11772 15252 11824
rect 15752 11815 15804 11824
rect 15752 11781 15761 11815
rect 15761 11781 15795 11815
rect 15795 11781 15804 11815
rect 15752 11772 15804 11781
rect 16764 11772 16816 11824
rect 14556 11704 14608 11756
rect 15292 11704 15344 11756
rect 16488 11704 16540 11756
rect 16580 11704 16632 11756
rect 22468 11772 22520 11824
rect 24584 11772 24636 11824
rect 24768 11840 24820 11892
rect 28724 11840 28776 11892
rect 30840 11840 30892 11892
rect 31208 11883 31260 11892
rect 31208 11849 31217 11883
rect 31217 11849 31251 11883
rect 31251 11849 31260 11883
rect 31208 11840 31260 11849
rect 32220 11840 32272 11892
rect 33600 11840 33652 11892
rect 20904 11704 20956 11756
rect 21088 11704 21140 11756
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 22652 11747 22704 11756
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 18420 11679 18472 11688
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 19984 11636 20036 11688
rect 23020 11704 23072 11756
rect 28356 11772 28408 11824
rect 30380 11772 30432 11824
rect 25964 11704 26016 11756
rect 23848 11679 23900 11688
rect 18512 11568 18564 11620
rect 21364 11568 21416 11620
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 28080 11704 28132 11756
rect 30196 11704 30248 11756
rect 32128 11704 32180 11756
rect 22100 11500 22152 11552
rect 22376 11500 22428 11552
rect 23388 11500 23440 11552
rect 26056 11543 26108 11552
rect 26056 11509 26065 11543
rect 26065 11509 26099 11543
rect 26099 11509 26108 11543
rect 26056 11500 26108 11509
rect 33416 11636 33468 11688
rect 28540 11568 28592 11620
rect 28724 11500 28776 11552
rect 31576 11543 31628 11552
rect 31576 11509 31585 11543
rect 31585 11509 31619 11543
rect 31619 11509 31628 11543
rect 31576 11500 31628 11509
rect 32312 11543 32364 11552
rect 32312 11509 32321 11543
rect 32321 11509 32355 11543
rect 32355 11509 32364 11543
rect 32312 11500 32364 11509
rect 5170 11398 5222 11450
rect 5234 11398 5286 11450
rect 5298 11398 5350 11450
rect 5362 11398 5414 11450
rect 5426 11398 5478 11450
rect 13611 11398 13663 11450
rect 13675 11398 13727 11450
rect 13739 11398 13791 11450
rect 13803 11398 13855 11450
rect 13867 11398 13919 11450
rect 22052 11398 22104 11450
rect 22116 11398 22168 11450
rect 22180 11398 22232 11450
rect 22244 11398 22296 11450
rect 22308 11398 22360 11450
rect 30493 11398 30545 11450
rect 30557 11398 30609 11450
rect 30621 11398 30673 11450
rect 30685 11398 30737 11450
rect 30749 11398 30801 11450
rect 4528 11296 4580 11348
rect 11244 11296 11296 11348
rect 12256 11296 12308 11348
rect 20536 11339 20588 11348
rect 20536 11305 20545 11339
rect 20545 11305 20579 11339
rect 20579 11305 20588 11339
rect 20536 11296 20588 11305
rect 20904 11296 20956 11348
rect 15844 11228 15896 11280
rect 12164 11160 12216 11212
rect 19524 11228 19576 11280
rect 21088 11228 21140 11280
rect 4528 11092 4580 11144
rect 7196 11092 7248 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 11060 11092 11112 11144
rect 11980 11092 12032 11144
rect 12532 11092 12584 11144
rect 12900 11092 12952 11144
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 18420 11160 18472 11212
rect 27988 11296 28040 11348
rect 28356 11296 28408 11348
rect 31208 11296 31260 11348
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 20076 11135 20128 11144
rect 20076 11101 20083 11135
rect 20083 11101 20128 11135
rect 20076 11092 20128 11101
rect 20168 11135 20220 11144
rect 20168 11101 20177 11135
rect 20177 11101 20211 11135
rect 20211 11101 20220 11135
rect 20168 11092 20220 11101
rect 21180 11135 21232 11144
rect 21180 11101 21189 11135
rect 21189 11101 21223 11135
rect 21223 11101 21232 11135
rect 21180 11092 21232 11101
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 25044 11228 25096 11280
rect 25780 11228 25832 11280
rect 26148 11160 26200 11212
rect 3792 11024 3844 11076
rect 5632 11024 5684 11076
rect 9312 11024 9364 11076
rect 4160 10999 4212 11008
rect 4160 10965 4185 10999
rect 4185 10965 4212 10999
rect 4344 10999 4396 11008
rect 4160 10956 4212 10965
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 7380 10956 7432 11008
rect 9772 10956 9824 11008
rect 11244 10956 11296 11008
rect 12440 11024 12492 11076
rect 12624 11067 12676 11076
rect 12624 11033 12633 11067
rect 12633 11033 12667 11067
rect 12667 11033 12676 11067
rect 12624 11024 12676 11033
rect 13452 11067 13504 11076
rect 13452 11033 13461 11067
rect 13461 11033 13495 11067
rect 13495 11033 13504 11067
rect 13452 11024 13504 11033
rect 16672 11067 16724 11076
rect 16672 11033 16681 11067
rect 16681 11033 16715 11067
rect 16715 11033 16724 11067
rect 16672 11024 16724 11033
rect 20536 11024 20588 11076
rect 20904 11024 20956 11076
rect 24584 11092 24636 11144
rect 26056 11135 26108 11144
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 29368 11092 29420 11144
rect 30932 11160 30984 11212
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 32220 11092 32272 11144
rect 12716 10956 12768 11008
rect 20444 10956 20496 11008
rect 24860 11024 24912 11076
rect 27712 11024 27764 11076
rect 31576 11024 31628 11076
rect 27344 10999 27396 11008
rect 27344 10965 27353 10999
rect 27353 10965 27387 10999
rect 27387 10965 27396 10999
rect 27344 10956 27396 10965
rect 29736 10999 29788 11008
rect 29736 10965 29745 10999
rect 29745 10965 29779 10999
rect 29779 10965 29788 10999
rect 29736 10956 29788 10965
rect 9390 10854 9442 10906
rect 9454 10854 9506 10906
rect 9518 10854 9570 10906
rect 9582 10854 9634 10906
rect 9646 10854 9698 10906
rect 17831 10854 17883 10906
rect 17895 10854 17947 10906
rect 17959 10854 18011 10906
rect 18023 10854 18075 10906
rect 18087 10854 18139 10906
rect 26272 10854 26324 10906
rect 26336 10854 26388 10906
rect 26400 10854 26452 10906
rect 26464 10854 26516 10906
rect 26528 10854 26580 10906
rect 34713 10854 34765 10906
rect 34777 10854 34829 10906
rect 34841 10854 34893 10906
rect 34905 10854 34957 10906
rect 34969 10854 35021 10906
rect 8116 10752 8168 10804
rect 8668 10752 8720 10804
rect 2964 10684 3016 10736
rect 3056 10616 3108 10668
rect 6736 10684 6788 10736
rect 6920 10684 6972 10736
rect 7380 10684 7432 10736
rect 7564 10727 7616 10736
rect 7564 10693 7573 10727
rect 7573 10693 7607 10727
rect 7607 10693 7616 10727
rect 7564 10684 7616 10693
rect 8576 10684 8628 10736
rect 9772 10752 9824 10804
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 10048 10752 10100 10804
rect 25504 10752 25556 10804
rect 28172 10795 28224 10804
rect 28172 10761 28181 10795
rect 28181 10761 28215 10795
rect 28215 10761 28224 10795
rect 28172 10752 28224 10761
rect 28724 10752 28776 10804
rect 33600 10752 33652 10804
rect 9404 10684 9456 10736
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 12900 10727 12952 10736
rect 12900 10693 12909 10727
rect 12909 10693 12943 10727
rect 12943 10693 12952 10727
rect 12900 10684 12952 10693
rect 13268 10727 13320 10736
rect 13268 10693 13277 10727
rect 13277 10693 13311 10727
rect 13311 10693 13320 10727
rect 13268 10684 13320 10693
rect 18236 10727 18288 10736
rect 18236 10693 18245 10727
rect 18245 10693 18279 10727
rect 18279 10693 18288 10727
rect 18236 10684 18288 10693
rect 19984 10727 20036 10736
rect 19984 10693 19993 10727
rect 19993 10693 20027 10727
rect 20027 10693 20036 10727
rect 19984 10684 20036 10693
rect 27344 10684 27396 10736
rect 30840 10727 30892 10736
rect 30840 10693 30849 10727
rect 30849 10693 30883 10727
rect 30883 10693 30892 10727
rect 30840 10684 30892 10693
rect 3884 10616 3936 10668
rect 4252 10616 4304 10668
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 6552 10548 6604 10600
rect 3516 10480 3568 10532
rect 12164 10616 12216 10668
rect 12440 10616 12492 10668
rect 25688 10616 25740 10668
rect 25872 10659 25924 10668
rect 25872 10625 25881 10659
rect 25881 10625 25915 10659
rect 25915 10625 25924 10659
rect 25872 10616 25924 10625
rect 25964 10659 26016 10668
rect 25964 10625 25973 10659
rect 25973 10625 26007 10659
rect 26007 10625 26016 10659
rect 26148 10659 26200 10668
rect 25964 10616 26016 10625
rect 26148 10625 26156 10659
rect 26156 10625 26190 10659
rect 26190 10625 26200 10659
rect 26148 10616 26200 10625
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 27712 10659 27764 10668
rect 27712 10625 27719 10659
rect 27719 10625 27764 10659
rect 27712 10616 27764 10625
rect 27896 10659 27948 10668
rect 27896 10625 27905 10659
rect 27905 10625 27939 10659
rect 27939 10625 27948 10659
rect 27896 10616 27948 10625
rect 28356 10616 28408 10668
rect 28908 10616 28960 10668
rect 29920 10616 29972 10668
rect 32312 10684 32364 10736
rect 27712 10480 27764 10532
rect 2780 10412 2832 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 10140 10455 10192 10464
rect 10140 10421 10149 10455
rect 10149 10421 10183 10455
rect 10183 10421 10192 10455
rect 10140 10412 10192 10421
rect 14372 10412 14424 10464
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 25964 10412 26016 10464
rect 28448 10548 28500 10600
rect 32220 10548 32272 10600
rect 31024 10455 31076 10464
rect 31024 10421 31033 10455
rect 31033 10421 31067 10455
rect 31067 10421 31076 10455
rect 31024 10412 31076 10421
rect 32312 10412 32364 10464
rect 5170 10310 5222 10362
rect 5234 10310 5286 10362
rect 5298 10310 5350 10362
rect 5362 10310 5414 10362
rect 5426 10310 5478 10362
rect 13611 10310 13663 10362
rect 13675 10310 13727 10362
rect 13739 10310 13791 10362
rect 13803 10310 13855 10362
rect 13867 10310 13919 10362
rect 22052 10310 22104 10362
rect 22116 10310 22168 10362
rect 22180 10310 22232 10362
rect 22244 10310 22296 10362
rect 22308 10310 22360 10362
rect 30493 10310 30545 10362
rect 30557 10310 30609 10362
rect 30621 10310 30673 10362
rect 30685 10310 30737 10362
rect 30749 10310 30801 10362
rect 3056 10208 3108 10260
rect 4068 10208 4120 10260
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 7564 10208 7616 10260
rect 8116 10208 8168 10260
rect 8668 10208 8720 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 25320 10208 25372 10260
rect 26148 10208 26200 10260
rect 26240 10208 26292 10260
rect 32220 10208 32272 10260
rect 3884 10072 3936 10124
rect 4252 10072 4304 10124
rect 8944 10140 8996 10192
rect 10048 10140 10100 10192
rect 27620 10140 27672 10192
rect 7196 10115 7248 10124
rect 2136 9911 2188 9920
rect 2136 9877 2145 9911
rect 2145 9877 2179 9911
rect 2179 9877 2188 9911
rect 2136 9868 2188 9877
rect 2780 10004 2832 10056
rect 4344 10004 4396 10056
rect 7196 10081 7205 10115
rect 7205 10081 7239 10115
rect 7239 10081 7248 10115
rect 7196 10072 7248 10081
rect 10324 10072 10376 10124
rect 19248 10072 19300 10124
rect 6828 10004 6880 10056
rect 7472 10047 7524 10056
rect 7472 10013 7506 10047
rect 7506 10013 7524 10047
rect 7472 10004 7524 10013
rect 17316 10047 17368 10056
rect 3976 9979 4028 9988
rect 3976 9945 3985 9979
rect 3985 9945 4019 9979
rect 4019 9945 4028 9979
rect 3976 9936 4028 9945
rect 5632 9979 5684 9988
rect 5632 9945 5666 9979
rect 5666 9945 5684 9979
rect 5632 9936 5684 9945
rect 11520 9979 11572 9988
rect 11520 9945 11554 9979
rect 11554 9945 11572 9979
rect 11520 9936 11572 9945
rect 11796 9936 11848 9988
rect 3332 9868 3384 9920
rect 8116 9868 8168 9920
rect 13360 9868 13412 9920
rect 16580 9868 16632 9920
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 20628 10047 20680 10056
rect 20628 10013 20637 10047
rect 20637 10013 20671 10047
rect 20671 10013 20680 10047
rect 20628 10004 20680 10013
rect 23848 10072 23900 10124
rect 28724 10115 28776 10124
rect 28724 10081 28733 10115
rect 28733 10081 28767 10115
rect 28767 10081 28776 10115
rect 28724 10072 28776 10081
rect 28908 10072 28960 10124
rect 17224 9979 17276 9988
rect 17224 9945 17233 9979
rect 17233 9945 17267 9979
rect 17267 9945 17276 9979
rect 21088 10047 21140 10056
rect 21088 10013 21102 10047
rect 21102 10013 21136 10047
rect 21136 10013 21140 10047
rect 24860 10047 24912 10056
rect 21088 10004 21140 10013
rect 24860 10013 24894 10047
rect 24894 10013 24912 10047
rect 24860 10004 24912 10013
rect 29736 10004 29788 10056
rect 29920 10047 29972 10056
rect 29920 10013 29929 10047
rect 29929 10013 29963 10047
rect 29963 10013 29972 10047
rect 29920 10004 29972 10013
rect 30288 10047 30340 10056
rect 30288 10013 30297 10047
rect 30297 10013 30331 10047
rect 30331 10013 30340 10047
rect 30288 10004 30340 10013
rect 33416 10047 33468 10056
rect 33416 10013 33425 10047
rect 33425 10013 33459 10047
rect 33459 10013 33468 10047
rect 33416 10004 33468 10013
rect 33692 10047 33744 10056
rect 33692 10013 33701 10047
rect 33701 10013 33735 10047
rect 33735 10013 33744 10047
rect 33692 10004 33744 10013
rect 17224 9936 17276 9945
rect 20444 9868 20496 9920
rect 20628 9868 20680 9920
rect 20812 9868 20864 9920
rect 29000 9936 29052 9988
rect 32220 9868 32272 9920
rect 33692 9868 33744 9920
rect 33876 9911 33928 9920
rect 33876 9877 33885 9911
rect 33885 9877 33919 9911
rect 33919 9877 33928 9911
rect 33876 9868 33928 9877
rect 9390 9766 9442 9818
rect 9454 9766 9506 9818
rect 9518 9766 9570 9818
rect 9582 9766 9634 9818
rect 9646 9766 9698 9818
rect 17831 9766 17883 9818
rect 17895 9766 17947 9818
rect 17959 9766 18011 9818
rect 18023 9766 18075 9818
rect 18087 9766 18139 9818
rect 26272 9766 26324 9818
rect 26336 9766 26388 9818
rect 26400 9766 26452 9818
rect 26464 9766 26516 9818
rect 26528 9766 26580 9818
rect 34713 9766 34765 9818
rect 34777 9766 34829 9818
rect 34841 9766 34893 9818
rect 34905 9766 34957 9818
rect 34969 9766 35021 9818
rect 4344 9664 4396 9716
rect 8576 9707 8628 9716
rect 8576 9673 8585 9707
rect 8585 9673 8619 9707
rect 8619 9673 8628 9707
rect 8576 9664 8628 9673
rect 10140 9664 10192 9716
rect 17132 9664 17184 9716
rect 27712 9707 27764 9716
rect 27712 9673 27721 9707
rect 27721 9673 27755 9707
rect 27755 9673 27764 9707
rect 27712 9664 27764 9673
rect 2504 9596 2556 9648
rect 3608 9596 3660 9648
rect 3976 9596 4028 9648
rect 7472 9639 7524 9648
rect 7472 9605 7506 9639
rect 7506 9605 7524 9639
rect 7472 9596 7524 9605
rect 17500 9596 17552 9648
rect 3148 9528 3200 9580
rect 4528 9571 4580 9580
rect 3056 9460 3108 9512
rect 2596 9324 2648 9376
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 4528 9537 4537 9571
rect 4537 9537 4571 9571
rect 4571 9537 4580 9571
rect 4528 9528 4580 9537
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4068 9460 4120 9512
rect 6828 9528 6880 9580
rect 11796 9528 11848 9580
rect 17408 9528 17460 9580
rect 17776 9571 17828 9580
rect 17776 9537 17785 9571
rect 17785 9537 17819 9571
rect 17819 9537 17828 9571
rect 17776 9528 17828 9537
rect 17868 9571 17920 9580
rect 17868 9537 17877 9571
rect 17877 9537 17911 9571
rect 17911 9537 17920 9571
rect 17868 9528 17920 9537
rect 18512 9571 18564 9580
rect 10784 9460 10836 9512
rect 17684 9460 17736 9512
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 12716 9392 12768 9444
rect 18328 9392 18380 9444
rect 18788 9528 18840 9580
rect 19340 9528 19392 9580
rect 19524 9596 19576 9648
rect 20352 9596 20404 9648
rect 20996 9596 21048 9648
rect 25688 9596 25740 9648
rect 31392 9639 31444 9648
rect 31392 9605 31401 9639
rect 31401 9605 31435 9639
rect 31435 9605 31444 9639
rect 31392 9596 31444 9605
rect 32312 9639 32364 9648
rect 32312 9605 32321 9639
rect 32321 9605 32355 9639
rect 32355 9605 32364 9639
rect 32312 9596 32364 9605
rect 20628 9571 20680 9580
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 18512 9324 18564 9376
rect 19248 9460 19300 9512
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 25964 9528 26016 9580
rect 27804 9528 27856 9580
rect 28908 9528 28960 9580
rect 30196 9528 30248 9580
rect 23664 9460 23716 9512
rect 29368 9460 29420 9512
rect 19800 9392 19852 9444
rect 19892 9392 19944 9444
rect 19340 9324 19392 9376
rect 21088 9392 21140 9444
rect 21180 9392 21232 9444
rect 27252 9392 27304 9444
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 20536 9324 20588 9376
rect 28816 9324 28868 9376
rect 31760 9367 31812 9376
rect 31760 9333 31769 9367
rect 31769 9333 31803 9367
rect 31803 9333 31812 9367
rect 31760 9324 31812 9333
rect 33692 9324 33744 9376
rect 5170 9222 5222 9274
rect 5234 9222 5286 9274
rect 5298 9222 5350 9274
rect 5362 9222 5414 9274
rect 5426 9222 5478 9274
rect 13611 9222 13663 9274
rect 13675 9222 13727 9274
rect 13739 9222 13791 9274
rect 13803 9222 13855 9274
rect 13867 9222 13919 9274
rect 22052 9222 22104 9274
rect 22116 9222 22168 9274
rect 22180 9222 22232 9274
rect 22244 9222 22296 9274
rect 22308 9222 22360 9274
rect 30493 9222 30545 9274
rect 30557 9222 30609 9274
rect 30621 9222 30673 9274
rect 30685 9222 30737 9274
rect 30749 9222 30801 9274
rect 2136 9120 2188 9172
rect 2688 9120 2740 9172
rect 12532 9120 12584 9172
rect 17224 9120 17276 9172
rect 20812 9120 20864 9172
rect 22836 9120 22888 9172
rect 27436 9120 27488 9172
rect 32220 9120 32272 9172
rect 2504 9052 2556 9104
rect 3700 9052 3752 9104
rect 2964 8984 3016 9036
rect 6828 8984 6880 9036
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 20996 8984 21048 9036
rect 4344 8916 4396 8968
rect 11060 8959 11112 8968
rect 11060 8925 11094 8959
rect 11094 8925 11112 8959
rect 11060 8916 11112 8925
rect 15108 8916 15160 8968
rect 16304 8916 16356 8968
rect 19524 8916 19576 8968
rect 19892 8959 19944 8968
rect 19892 8925 19901 8959
rect 19901 8925 19935 8959
rect 19935 8925 19944 8959
rect 19892 8916 19944 8925
rect 20444 8916 20496 8968
rect 22836 8959 22888 8968
rect 22836 8925 22845 8959
rect 22845 8925 22879 8959
rect 22879 8925 22888 8959
rect 22836 8916 22888 8925
rect 24584 8959 24636 8968
rect 2872 8848 2924 8900
rect 16580 8848 16632 8900
rect 17408 8848 17460 8900
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 17224 8780 17276 8832
rect 17868 8848 17920 8900
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 23664 8848 23716 8900
rect 28816 8959 28868 8968
rect 28816 8925 28825 8959
rect 28825 8925 28859 8959
rect 28859 8925 28868 8959
rect 30380 9052 30432 9104
rect 28816 8916 28868 8925
rect 29092 8916 29144 8968
rect 30196 8959 30248 8968
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 32312 8916 32364 8968
rect 30288 8848 30340 8900
rect 33876 8848 33928 8900
rect 17776 8780 17828 8832
rect 20444 8780 20496 8832
rect 21824 8780 21876 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 25780 8780 25832 8832
rect 28908 8780 28960 8832
rect 29000 8780 29052 8832
rect 29184 8823 29236 8832
rect 29184 8789 29193 8823
rect 29193 8789 29227 8823
rect 29227 8789 29236 8823
rect 29184 8780 29236 8789
rect 29736 8823 29788 8832
rect 29736 8789 29745 8823
rect 29745 8789 29779 8823
rect 29779 8789 29788 8823
rect 29736 8780 29788 8789
rect 9390 8678 9442 8730
rect 9454 8678 9506 8730
rect 9518 8678 9570 8730
rect 9582 8678 9634 8730
rect 9646 8678 9698 8730
rect 17831 8678 17883 8730
rect 17895 8678 17947 8730
rect 17959 8678 18011 8730
rect 18023 8678 18075 8730
rect 18087 8678 18139 8730
rect 26272 8678 26324 8730
rect 26336 8678 26388 8730
rect 26400 8678 26452 8730
rect 26464 8678 26516 8730
rect 26528 8678 26580 8730
rect 34713 8678 34765 8730
rect 34777 8678 34829 8730
rect 34841 8678 34893 8730
rect 34905 8678 34957 8730
rect 34969 8678 35021 8730
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 17684 8576 17736 8628
rect 12072 8508 12124 8560
rect 17316 8508 17368 8560
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 2780 8440 2832 8492
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 17040 8440 17092 8492
rect 20904 8576 20956 8628
rect 22560 8576 22612 8628
rect 23664 8619 23716 8628
rect 18512 8508 18564 8560
rect 20996 8508 21048 8560
rect 22744 8551 22796 8560
rect 22744 8517 22753 8551
rect 22753 8517 22787 8551
rect 22787 8517 22796 8551
rect 22744 8508 22796 8517
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 25688 8576 25740 8628
rect 25872 8619 25924 8628
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 28908 8576 28960 8628
rect 25044 8508 25096 8560
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 20536 8440 20588 8492
rect 21088 8440 21140 8492
rect 24952 8440 25004 8492
rect 25780 8440 25832 8492
rect 26056 8440 26108 8492
rect 29092 8508 29144 8560
rect 30288 8576 30340 8628
rect 31392 8576 31444 8628
rect 29736 8440 29788 8492
rect 30196 8440 30248 8492
rect 30840 8483 30892 8492
rect 18328 8372 18380 8424
rect 19892 8372 19944 8424
rect 21272 8372 21324 8424
rect 25044 8415 25096 8424
rect 25044 8381 25053 8415
rect 25053 8381 25087 8415
rect 25087 8381 25096 8415
rect 25044 8372 25096 8381
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 31760 8508 31812 8560
rect 32128 8440 32180 8492
rect 32312 8483 32364 8492
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 19708 8304 19760 8356
rect 21180 8304 21232 8356
rect 24032 8304 24084 8356
rect 8208 8236 8260 8288
rect 16672 8236 16724 8288
rect 18512 8236 18564 8288
rect 21732 8236 21784 8288
rect 28080 8236 28132 8288
rect 5170 8134 5222 8186
rect 5234 8134 5286 8186
rect 5298 8134 5350 8186
rect 5362 8134 5414 8186
rect 5426 8134 5478 8186
rect 13611 8134 13663 8186
rect 13675 8134 13727 8186
rect 13739 8134 13791 8186
rect 13803 8134 13855 8186
rect 13867 8134 13919 8186
rect 22052 8134 22104 8186
rect 22116 8134 22168 8186
rect 22180 8134 22232 8186
rect 22244 8134 22296 8186
rect 22308 8134 22360 8186
rect 30493 8134 30545 8186
rect 30557 8134 30609 8186
rect 30621 8134 30673 8186
rect 30685 8134 30737 8186
rect 30749 8134 30801 8186
rect 18236 8032 18288 8084
rect 28080 8032 28132 8084
rect 32312 8032 32364 8084
rect 8208 7828 8260 7880
rect 7380 7803 7432 7812
rect 7380 7769 7389 7803
rect 7389 7769 7423 7803
rect 7423 7769 7432 7803
rect 7380 7760 7432 7769
rect 8116 7760 8168 7812
rect 20720 7828 20772 7880
rect 24032 7828 24084 7880
rect 33692 7871 33744 7880
rect 33692 7837 33701 7871
rect 33701 7837 33735 7871
rect 33735 7837 33744 7871
rect 33692 7828 33744 7837
rect 10232 7760 10284 7812
rect 15936 7760 15988 7812
rect 20812 7760 20864 7812
rect 28080 7803 28132 7812
rect 28080 7769 28089 7803
rect 28089 7769 28123 7803
rect 28123 7769 28132 7803
rect 28080 7760 28132 7769
rect 28356 7760 28408 7812
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 20444 7692 20496 7744
rect 23388 7692 23440 7744
rect 30380 7692 30432 7744
rect 9390 7590 9442 7642
rect 9454 7590 9506 7642
rect 9518 7590 9570 7642
rect 9582 7590 9634 7642
rect 9646 7590 9698 7642
rect 17831 7590 17883 7642
rect 17895 7590 17947 7642
rect 17959 7590 18011 7642
rect 18023 7590 18075 7642
rect 18087 7590 18139 7642
rect 26272 7590 26324 7642
rect 26336 7590 26388 7642
rect 26400 7590 26452 7642
rect 26464 7590 26516 7642
rect 26528 7590 26580 7642
rect 34713 7590 34765 7642
rect 34777 7590 34829 7642
rect 34841 7590 34893 7642
rect 34905 7590 34957 7642
rect 34969 7590 35021 7642
rect 10508 7488 10560 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 17408 7488 17460 7540
rect 19524 7531 19576 7540
rect 5632 7420 5684 7472
rect 7380 7420 7432 7472
rect 10232 7420 10284 7472
rect 15200 7420 15252 7472
rect 16672 7420 16724 7472
rect 3792 7352 3844 7404
rect 8392 7352 8444 7404
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 17592 7420 17644 7472
rect 19524 7497 19533 7531
rect 19533 7497 19567 7531
rect 19567 7497 19576 7531
rect 19524 7488 19576 7497
rect 20536 7488 20588 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 20996 7488 21048 7540
rect 25964 7531 26016 7540
rect 25964 7497 25973 7531
rect 25973 7497 26007 7531
rect 26007 7497 26016 7531
rect 25964 7488 26016 7497
rect 29092 7531 29144 7540
rect 29092 7497 29101 7531
rect 29101 7497 29135 7531
rect 29135 7497 29144 7531
rect 29092 7488 29144 7497
rect 20444 7463 20496 7472
rect 20444 7429 20453 7463
rect 20453 7429 20487 7463
rect 20487 7429 20496 7463
rect 20444 7420 20496 7429
rect 20904 7420 20956 7472
rect 23388 7463 23440 7472
rect 17684 7395 17736 7404
rect 11060 7284 11112 7336
rect 11244 7284 11296 7336
rect 13084 7284 13136 7336
rect 17040 7284 17092 7336
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 17868 7352 17920 7404
rect 22376 7352 22428 7404
rect 23388 7429 23397 7463
rect 23397 7429 23431 7463
rect 23431 7429 23440 7463
rect 23388 7420 23440 7429
rect 25044 7463 25096 7472
rect 25044 7429 25053 7463
rect 25053 7429 25087 7463
rect 25087 7429 25096 7463
rect 25044 7420 25096 7429
rect 29368 7420 29420 7472
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 15108 7148 15160 7200
rect 15660 7148 15712 7200
rect 19432 7148 19484 7200
rect 21732 7216 21784 7268
rect 23756 7284 23808 7336
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 30380 7395 30432 7404
rect 30380 7361 30389 7395
rect 30389 7361 30423 7395
rect 30423 7361 30432 7395
rect 30380 7352 30432 7361
rect 24032 7284 24084 7336
rect 24584 7284 24636 7336
rect 20720 7148 20772 7200
rect 25596 7191 25648 7200
rect 25596 7157 25605 7191
rect 25605 7157 25639 7191
rect 25639 7157 25648 7191
rect 25596 7148 25648 7157
rect 5170 7046 5222 7098
rect 5234 7046 5286 7098
rect 5298 7046 5350 7098
rect 5362 7046 5414 7098
rect 5426 7046 5478 7098
rect 13611 7046 13663 7098
rect 13675 7046 13727 7098
rect 13739 7046 13791 7098
rect 13803 7046 13855 7098
rect 13867 7046 13919 7098
rect 22052 7046 22104 7098
rect 22116 7046 22168 7098
rect 22180 7046 22232 7098
rect 22244 7046 22296 7098
rect 22308 7046 22360 7098
rect 30493 7046 30545 7098
rect 30557 7046 30609 7098
rect 30621 7046 30673 7098
rect 30685 7046 30737 7098
rect 30749 7046 30801 7098
rect 2596 6944 2648 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 3148 6808 3200 6860
rect 3792 6808 3844 6860
rect 4344 6808 4396 6860
rect 5080 6808 5132 6860
rect 5724 6783 5776 6792
rect 5724 6749 5758 6783
rect 5758 6749 5776 6783
rect 5724 6740 5776 6749
rect 2872 6672 2924 6724
rect 8300 6808 8352 6860
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 15108 6808 15160 6860
rect 10416 6740 10468 6792
rect 10508 6740 10560 6792
rect 11244 6740 11296 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 11060 6672 11112 6724
rect 6920 6604 6972 6656
rect 8300 6604 8352 6656
rect 12808 6672 12860 6724
rect 15660 6740 15712 6792
rect 17224 6740 17276 6792
rect 17868 6876 17920 6928
rect 20352 6944 20404 6996
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 22652 6808 22704 6860
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 19524 6740 19576 6792
rect 19708 6783 19760 6792
rect 19708 6749 19742 6783
rect 19742 6749 19760 6783
rect 19708 6740 19760 6749
rect 21824 6740 21876 6792
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 24032 6783 24084 6792
rect 24032 6749 24041 6783
rect 24041 6749 24075 6783
rect 24075 6749 24084 6783
rect 24032 6740 24084 6749
rect 28908 6783 28960 6792
rect 28908 6749 28926 6783
rect 28926 6749 28960 6783
rect 28908 6740 28960 6749
rect 29092 6740 29144 6792
rect 29828 6740 29880 6792
rect 17500 6672 17552 6724
rect 24952 6672 25004 6724
rect 25044 6672 25096 6724
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 18328 6604 18380 6656
rect 22836 6604 22888 6656
rect 23572 6647 23624 6656
rect 23572 6613 23581 6647
rect 23581 6613 23615 6647
rect 23615 6613 23624 6647
rect 23572 6604 23624 6613
rect 25872 6604 25924 6656
rect 28264 6672 28316 6724
rect 29276 6672 29328 6724
rect 27896 6604 27948 6656
rect 9390 6502 9442 6554
rect 9454 6502 9506 6554
rect 9518 6502 9570 6554
rect 9582 6502 9634 6554
rect 9646 6502 9698 6554
rect 17831 6502 17883 6554
rect 17895 6502 17947 6554
rect 17959 6502 18011 6554
rect 18023 6502 18075 6554
rect 18087 6502 18139 6554
rect 26272 6502 26324 6554
rect 26336 6502 26388 6554
rect 26400 6502 26452 6554
rect 26464 6502 26516 6554
rect 26528 6502 26580 6554
rect 34713 6502 34765 6554
rect 34777 6502 34829 6554
rect 34841 6502 34893 6554
rect 34905 6502 34957 6554
rect 34969 6502 35021 6554
rect 2872 6400 2924 6452
rect 6920 6443 6972 6452
rect 6920 6409 6929 6443
rect 6929 6409 6963 6443
rect 6963 6409 6972 6443
rect 6920 6400 6972 6409
rect 12532 6400 12584 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 28264 6400 28316 6452
rect 30840 6400 30892 6452
rect 3792 6332 3844 6384
rect 7012 6332 7064 6384
rect 13636 6332 13688 6384
rect 20720 6332 20772 6384
rect 23572 6332 23624 6384
rect 29184 6332 29236 6384
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 4068 6196 4120 6248
rect 6092 6196 6144 6248
rect 12440 6196 12492 6248
rect 19524 6196 19576 6248
rect 29828 6239 29880 6248
rect 18420 6128 18472 6180
rect 22652 6128 22704 6180
rect 3976 6060 4028 6112
rect 19984 6060 20036 6112
rect 24676 6060 24728 6112
rect 29828 6205 29837 6239
rect 29837 6205 29871 6239
rect 29871 6205 29880 6239
rect 29828 6196 29880 6205
rect 28816 6128 28868 6180
rect 5170 5958 5222 6010
rect 5234 5958 5286 6010
rect 5298 5958 5350 6010
rect 5362 5958 5414 6010
rect 5426 5958 5478 6010
rect 13611 5958 13663 6010
rect 13675 5958 13727 6010
rect 13739 5958 13791 6010
rect 13803 5958 13855 6010
rect 13867 5958 13919 6010
rect 22052 5958 22104 6010
rect 22116 5958 22168 6010
rect 22180 5958 22232 6010
rect 22244 5958 22296 6010
rect 22308 5958 22360 6010
rect 30493 5958 30545 6010
rect 30557 5958 30609 6010
rect 30621 5958 30673 6010
rect 30685 5958 30737 6010
rect 30749 5958 30801 6010
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 29276 5856 29328 5908
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 5632 5720 5684 5772
rect 24676 5652 24728 5704
rect 25596 5652 25648 5704
rect 29000 5788 29052 5840
rect 29368 5652 29420 5704
rect 4712 5584 4764 5636
rect 4068 5516 4120 5568
rect 8208 5584 8260 5636
rect 27896 5584 27948 5636
rect 6092 5559 6144 5568
rect 6092 5525 6101 5559
rect 6101 5525 6135 5559
rect 6135 5525 6144 5559
rect 6092 5516 6144 5525
rect 9390 5414 9442 5466
rect 9454 5414 9506 5466
rect 9518 5414 9570 5466
rect 9582 5414 9634 5466
rect 9646 5414 9698 5466
rect 17831 5414 17883 5466
rect 17895 5414 17947 5466
rect 17959 5414 18011 5466
rect 18023 5414 18075 5466
rect 18087 5414 18139 5466
rect 26272 5414 26324 5466
rect 26336 5414 26388 5466
rect 26400 5414 26452 5466
rect 26464 5414 26516 5466
rect 26528 5414 26580 5466
rect 34713 5414 34765 5466
rect 34777 5414 34829 5466
rect 34841 5414 34893 5466
rect 34905 5414 34957 5466
rect 34969 5414 35021 5466
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6092 5312 6144 5364
rect 10508 5355 10560 5364
rect 2964 5244 3016 5296
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 4712 5244 4764 5296
rect 9312 5244 9364 5296
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 13176 5312 13228 5364
rect 19524 5355 19576 5364
rect 12440 5244 12492 5296
rect 5632 5108 5684 5160
rect 6552 5108 6604 5160
rect 9864 5176 9916 5228
rect 10876 5176 10928 5228
rect 11796 5176 11848 5228
rect 10692 5108 10744 5160
rect 11704 5151 11756 5160
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 7196 5040 7248 5092
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 18236 5287 18288 5296
rect 18236 5253 18245 5287
rect 18245 5253 18279 5287
rect 18279 5253 18288 5287
rect 18236 5244 18288 5253
rect 23388 5287 23440 5296
rect 23388 5253 23397 5287
rect 23397 5253 23431 5287
rect 23431 5253 23440 5287
rect 23388 5244 23440 5253
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 17408 5176 17460 5228
rect 25780 5219 25832 5228
rect 25780 5185 25789 5219
rect 25789 5185 25823 5219
rect 25823 5185 25832 5219
rect 25780 5176 25832 5185
rect 26608 5108 26660 5160
rect 8116 4972 8168 5024
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 11244 4972 11296 5024
rect 11980 4972 12032 5024
rect 25044 5040 25096 5092
rect 14280 4972 14332 5024
rect 14924 4972 14976 5024
rect 25688 4972 25740 5024
rect 5170 4870 5222 4922
rect 5234 4870 5286 4922
rect 5298 4870 5350 4922
rect 5362 4870 5414 4922
rect 5426 4870 5478 4922
rect 13611 4870 13663 4922
rect 13675 4870 13727 4922
rect 13739 4870 13791 4922
rect 13803 4870 13855 4922
rect 13867 4870 13919 4922
rect 22052 4870 22104 4922
rect 22116 4870 22168 4922
rect 22180 4870 22232 4922
rect 22244 4870 22296 4922
rect 22308 4870 22360 4922
rect 30493 4870 30545 4922
rect 30557 4870 30609 4922
rect 30621 4870 30673 4922
rect 30685 4870 30737 4922
rect 30749 4870 30801 4922
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11980 4811 12032 4820
rect 11980 4777 11989 4811
rect 11989 4777 12023 4811
rect 12023 4777 12032 4811
rect 11980 4768 12032 4777
rect 5080 4632 5132 4684
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 8944 4632 8996 4684
rect 7472 4607 7524 4616
rect 7472 4573 7506 4607
rect 7506 4573 7524 4607
rect 7472 4564 7524 4573
rect 10508 4564 10560 4616
rect 20720 4700 20772 4752
rect 24676 4743 24728 4752
rect 24676 4709 24685 4743
rect 24685 4709 24719 4743
rect 24719 4709 24728 4743
rect 24676 4700 24728 4709
rect 14188 4632 14240 4684
rect 12440 4564 12492 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 20444 4675 20496 4684
rect 20444 4641 20453 4675
rect 20453 4641 20487 4675
rect 20487 4641 20496 4675
rect 20444 4632 20496 4641
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 15844 4564 15896 4616
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 19984 4564 20036 4616
rect 20904 4564 20956 4616
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 25872 4564 25924 4573
rect 11796 4496 11848 4548
rect 26148 4539 26200 4548
rect 26148 4505 26182 4539
rect 26182 4505 26200 4539
rect 26148 4496 26200 4505
rect 9772 4428 9824 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16304 4428 16356 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 18236 4428 18288 4480
rect 19064 4428 19116 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 20812 4428 20864 4480
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 22100 4428 22152 4480
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 26792 4428 26844 4480
rect 9390 4326 9442 4378
rect 9454 4326 9506 4378
rect 9518 4326 9570 4378
rect 9582 4326 9634 4378
rect 9646 4326 9698 4378
rect 17831 4326 17883 4378
rect 17895 4326 17947 4378
rect 17959 4326 18011 4378
rect 18023 4326 18075 4378
rect 18087 4326 18139 4378
rect 26272 4326 26324 4378
rect 26336 4326 26388 4378
rect 26400 4326 26452 4378
rect 26464 4326 26516 4378
rect 26528 4326 26580 4378
rect 34713 4326 34765 4378
rect 34777 4326 34829 4378
rect 34841 4326 34893 4378
rect 34905 4326 34957 4378
rect 34969 4326 35021 4378
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 7472 4156 7524 4208
rect 7932 4156 7984 4208
rect 8944 4088 8996 4140
rect 9864 4224 9916 4276
rect 9956 4224 10008 4276
rect 22468 4224 22520 4276
rect 26148 4267 26200 4276
rect 26148 4233 26157 4267
rect 26157 4233 26191 4267
rect 26191 4233 26200 4267
rect 26148 4224 26200 4233
rect 13360 4199 13412 4208
rect 13360 4165 13369 4199
rect 13369 4165 13403 4199
rect 13403 4165 13412 4199
rect 13360 4156 13412 4165
rect 15568 4156 15620 4208
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 10508 4131 10560 4140
rect 9772 4088 9824 4097
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10876 4131 10928 4140
rect 10600 4088 10652 4097
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 14004 4088 14056 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 17408 4088 17460 4140
rect 17500 4088 17552 4140
rect 17960 4131 18012 4140
rect 17960 4097 17994 4131
rect 17994 4097 18012 4131
rect 17960 4088 18012 4097
rect 19708 4088 19760 4140
rect 20904 4088 20956 4140
rect 21180 4131 21232 4140
rect 21180 4097 21198 4131
rect 21198 4097 21232 4131
rect 21180 4088 21232 4097
rect 21548 4088 21600 4140
rect 22100 4088 22152 4140
rect 22284 4131 22336 4140
rect 22284 4097 22318 4131
rect 22318 4097 22336 4131
rect 25872 4156 25924 4208
rect 22284 4088 22336 4097
rect 24584 4131 24636 4140
rect 24584 4097 24618 4131
rect 24618 4097 24636 4131
rect 24584 4088 24636 4097
rect 26608 4131 26660 4140
rect 26608 4097 26617 4131
rect 26617 4097 26651 4131
rect 26651 4097 26660 4131
rect 26608 4088 26660 4097
rect 27068 4088 27120 4140
rect 28080 4156 28132 4208
rect 27804 4088 27856 4140
rect 11244 4020 11296 4072
rect 14188 4020 14240 4072
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16672 3884 16724 3936
rect 19064 3927 19116 3936
rect 19064 3893 19073 3927
rect 19073 3893 19107 3927
rect 19107 3893 19116 3927
rect 19064 3884 19116 3893
rect 21088 3884 21140 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 26608 3884 26660 3936
rect 28356 3884 28408 3936
rect 5170 3782 5222 3834
rect 5234 3782 5286 3834
rect 5298 3782 5350 3834
rect 5362 3782 5414 3834
rect 5426 3782 5478 3834
rect 13611 3782 13663 3834
rect 13675 3782 13727 3834
rect 13739 3782 13791 3834
rect 13803 3782 13855 3834
rect 13867 3782 13919 3834
rect 22052 3782 22104 3834
rect 22116 3782 22168 3834
rect 22180 3782 22232 3834
rect 22244 3782 22296 3834
rect 22308 3782 22360 3834
rect 30493 3782 30545 3834
rect 30557 3782 30609 3834
rect 30621 3782 30673 3834
rect 30685 3782 30737 3834
rect 30749 3782 30801 3834
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 14004 3680 14056 3732
rect 16856 3680 16908 3732
rect 20812 3723 20864 3732
rect 20812 3689 20821 3723
rect 20821 3689 20855 3723
rect 20855 3689 20864 3723
rect 20812 3680 20864 3689
rect 22376 3680 22428 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 27804 3723 27856 3732
rect 27804 3689 27813 3723
rect 27813 3689 27847 3723
rect 27847 3689 27856 3723
rect 27804 3680 27856 3689
rect 26792 3655 26844 3664
rect 26792 3621 26801 3655
rect 26801 3621 26835 3655
rect 26835 3621 26844 3655
rect 26792 3612 26844 3621
rect 8208 3544 8260 3596
rect 10876 3544 10928 3596
rect 16672 3587 16724 3596
rect 16672 3553 16681 3587
rect 16681 3553 16715 3587
rect 16715 3553 16724 3587
rect 16672 3544 16724 3553
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 26148 3544 26200 3596
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 10600 3476 10652 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 12992 3476 13044 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 23388 3476 23440 3528
rect 25688 3519 25740 3528
rect 25688 3485 25706 3519
rect 25706 3485 25740 3519
rect 25688 3476 25740 3485
rect 25872 3476 25924 3528
rect 26608 3476 26660 3528
rect 27620 3612 27672 3664
rect 27160 3544 27212 3596
rect 14740 3408 14792 3460
rect 16948 3451 17000 3460
rect 16948 3417 16982 3451
rect 16982 3417 17000 3451
rect 16948 3408 17000 3417
rect 19800 3408 19852 3460
rect 25780 3408 25832 3460
rect 28356 3476 28408 3528
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 18236 3340 18288 3392
rect 9390 3238 9442 3290
rect 9454 3238 9506 3290
rect 9518 3238 9570 3290
rect 9582 3238 9634 3290
rect 9646 3238 9698 3290
rect 17831 3238 17883 3290
rect 17895 3238 17947 3290
rect 17959 3238 18011 3290
rect 18023 3238 18075 3290
rect 18087 3238 18139 3290
rect 26272 3238 26324 3290
rect 26336 3238 26388 3290
rect 26400 3238 26452 3290
rect 26464 3238 26516 3290
rect 26528 3238 26580 3290
rect 34713 3238 34765 3290
rect 34777 3238 34829 3290
rect 34841 3238 34893 3290
rect 34905 3238 34957 3290
rect 34969 3238 35021 3290
rect 12348 3136 12400 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14740 3179 14792 3188
rect 14740 3145 14749 3179
rect 14749 3145 14783 3179
rect 14783 3145 14792 3179
rect 14740 3136 14792 3145
rect 15660 3136 15712 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 17132 3136 17184 3188
rect 18236 3136 18288 3188
rect 19432 3136 19484 3188
rect 21180 3136 21232 3188
rect 29828 3136 29880 3188
rect 21088 3111 21140 3120
rect 10876 3000 10928 3052
rect 21088 3077 21097 3111
rect 21097 3077 21131 3111
rect 21131 3077 21140 3111
rect 21088 3068 21140 3077
rect 30380 3111 30432 3120
rect 30380 3077 30389 3111
rect 30389 3077 30423 3111
rect 30423 3077 30432 3111
rect 30380 3068 30432 3077
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 20720 3000 20772 3052
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 15476 2932 15528 2984
rect 20444 2932 20496 2984
rect 22744 3000 22796 3052
rect 26792 3000 26844 3052
rect 27620 3000 27672 3052
rect 25044 2932 25096 2984
rect 26148 2932 26200 2984
rect 25780 2796 25832 2848
rect 26240 2796 26292 2848
rect 26608 2796 26660 2848
rect 5170 2694 5222 2746
rect 5234 2694 5286 2746
rect 5298 2694 5350 2746
rect 5362 2694 5414 2746
rect 5426 2694 5478 2746
rect 13611 2694 13663 2746
rect 13675 2694 13727 2746
rect 13739 2694 13791 2746
rect 13803 2694 13855 2746
rect 13867 2694 13919 2746
rect 22052 2694 22104 2746
rect 22116 2694 22168 2746
rect 22180 2694 22232 2746
rect 22244 2694 22296 2746
rect 22308 2694 22360 2746
rect 30493 2694 30545 2746
rect 30557 2694 30609 2746
rect 30621 2694 30673 2746
rect 30685 2694 30737 2746
rect 30749 2694 30801 2746
rect 1216 2320 1268 2372
rect 2504 2320 2556 2372
rect 3792 2320 3844 2372
rect 15936 2592 15988 2644
rect 10140 2524 10192 2576
rect 5080 2320 5132 2372
rect 6368 2388 6420 2440
rect 7564 2320 7616 2372
rect 14372 2456 14424 2508
rect 18236 2456 18288 2508
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8944 2388 8996 2440
rect 10232 2388 10284 2440
rect 11520 2388 11572 2440
rect 12808 2388 12860 2440
rect 14004 2388 14056 2440
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16304 2388 16356 2440
rect 19064 2388 19116 2440
rect 20812 2388 20864 2440
rect 21088 2388 21140 2440
rect 23388 2388 23440 2440
rect 25044 2431 25096 2440
rect 25044 2397 25053 2431
rect 25053 2397 25087 2431
rect 25087 2397 25096 2431
rect 25044 2388 25096 2397
rect 26240 2431 26292 2440
rect 26240 2397 26249 2431
rect 26249 2397 26283 2431
rect 26283 2397 26292 2431
rect 27620 2431 27672 2440
rect 26240 2388 26292 2397
rect 27620 2397 27629 2431
rect 27629 2397 27663 2431
rect 27663 2397 27672 2431
rect 27620 2388 27672 2397
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 29552 2388 29604 2440
rect 30840 2388 30892 2440
rect 32128 2388 32180 2440
rect 33416 2388 33468 2440
rect 14096 2320 14148 2372
rect 15384 2320 15436 2372
rect 16672 2320 16724 2372
rect 18236 2320 18288 2372
rect 19248 2320 19300 2372
rect 20536 2320 20588 2372
rect 21824 2320 21876 2372
rect 23112 2320 23164 2372
rect 24400 2320 24452 2372
rect 25688 2320 25740 2372
rect 26976 2320 27028 2372
rect 28264 2320 28316 2372
rect 34612 2252 34664 2304
rect 9390 2150 9442 2202
rect 9454 2150 9506 2202
rect 9518 2150 9570 2202
rect 9582 2150 9634 2202
rect 9646 2150 9698 2202
rect 17831 2150 17883 2202
rect 17895 2150 17947 2202
rect 17959 2150 18011 2202
rect 18023 2150 18075 2202
rect 18087 2150 18139 2202
rect 26272 2150 26324 2202
rect 26336 2150 26388 2202
rect 26400 2150 26452 2202
rect 26464 2150 26516 2202
rect 26528 2150 26580 2202
rect 34713 2150 34765 2202
rect 34777 2150 34829 2202
rect 34841 2150 34893 2202
rect 34905 2150 34957 2202
rect 34969 2150 35021 2202
<< metal2 >>
rect 1766 35306 1822 36000
rect 1412 35278 1822 35306
rect 1412 14482 1440 35278
rect 1766 35200 1822 35278
rect 4710 35306 4766 36000
rect 7654 35306 7710 36000
rect 4710 35278 4936 35306
rect 4710 35200 4766 35278
rect 4908 33590 4936 35278
rect 7654 35278 7880 35306
rect 7654 35200 7710 35278
rect 7852 33590 7880 35278
rect 10598 35200 10654 36000
rect 13542 35306 13598 36000
rect 13542 35278 13768 35306
rect 13542 35200 13598 35278
rect 9390 33756 9698 33765
rect 9390 33754 9396 33756
rect 9452 33754 9476 33756
rect 9532 33754 9556 33756
rect 9612 33754 9636 33756
rect 9692 33754 9698 33756
rect 9452 33702 9454 33754
rect 9634 33702 9636 33754
rect 9390 33700 9396 33702
rect 9452 33700 9476 33702
rect 9532 33700 9556 33702
rect 9612 33700 9636 33702
rect 9692 33700 9698 33702
rect 9390 33691 9698 33700
rect 10612 33590 10640 35200
rect 4896 33584 4948 33590
rect 4896 33526 4948 33532
rect 7840 33584 7892 33590
rect 7840 33526 7892 33532
rect 10600 33584 10652 33590
rect 13740 33572 13768 35278
rect 16486 35200 16542 36000
rect 19430 35200 19486 36000
rect 22374 35306 22430 36000
rect 25318 35306 25374 36000
rect 28262 35306 28318 36000
rect 31206 35306 31262 36000
rect 34150 35306 34206 36000
rect 22374 35278 22692 35306
rect 22374 35200 22430 35278
rect 13820 33584 13872 33590
rect 13740 33544 13820 33572
rect 10600 33526 10652 33532
rect 16500 33572 16528 35200
rect 17831 33756 18139 33765
rect 17831 33754 17837 33756
rect 17893 33754 17917 33756
rect 17973 33754 17997 33756
rect 18053 33754 18077 33756
rect 18133 33754 18139 33756
rect 17893 33702 17895 33754
rect 18075 33702 18077 33754
rect 17831 33700 17837 33702
rect 17893 33700 17917 33702
rect 17973 33700 17997 33702
rect 18053 33700 18077 33702
rect 18133 33700 18139 33702
rect 17831 33691 18139 33700
rect 19444 33590 19472 35200
rect 22664 33590 22692 35278
rect 25318 35278 25636 35306
rect 25318 35200 25374 35278
rect 25608 33590 25636 35278
rect 28262 35278 28580 35306
rect 28262 35200 28318 35278
rect 26272 33756 26580 33765
rect 26272 33754 26278 33756
rect 26334 33754 26358 33756
rect 26414 33754 26438 33756
rect 26494 33754 26518 33756
rect 26574 33754 26580 33756
rect 26334 33702 26336 33754
rect 26516 33702 26518 33754
rect 26272 33700 26278 33702
rect 26334 33700 26358 33702
rect 26414 33700 26438 33702
rect 26494 33700 26518 33702
rect 26574 33700 26580 33702
rect 26272 33691 26580 33700
rect 28552 33590 28580 35278
rect 31206 35278 31524 35306
rect 31206 35200 31262 35278
rect 31496 33590 31524 35278
rect 34150 35278 34284 35306
rect 34150 35200 34206 35278
rect 34256 33590 34284 35278
rect 34713 33756 35021 33765
rect 34713 33754 34719 33756
rect 34775 33754 34799 33756
rect 34855 33754 34879 33756
rect 34935 33754 34959 33756
rect 35015 33754 35021 33756
rect 34775 33702 34777 33754
rect 34957 33702 34959 33754
rect 34713 33700 34719 33702
rect 34775 33700 34799 33702
rect 34855 33700 34879 33702
rect 34935 33700 34959 33702
rect 35015 33700 35021 33702
rect 34713 33691 35021 33700
rect 16580 33584 16632 33590
rect 16500 33544 16580 33572
rect 13820 33526 13872 33532
rect 16580 33526 16632 33532
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 22652 33584 22704 33590
rect 22652 33526 22704 33532
rect 25596 33584 25648 33590
rect 25596 33526 25648 33532
rect 28540 33584 28592 33590
rect 28540 33526 28592 33532
rect 31484 33584 31536 33590
rect 31484 33526 31536 33532
rect 34244 33584 34296 33590
rect 34244 33526 34296 33532
rect 8024 33380 8076 33386
rect 8024 33322 8076 33328
rect 12256 33380 12308 33386
rect 12256 33322 12308 33328
rect 14280 33380 14332 33386
rect 14280 33322 14332 33328
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 20260 33380 20312 33386
rect 20260 33322 20312 33328
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 31300 33380 31352 33386
rect 31300 33322 31352 33328
rect 33324 33380 33376 33386
rect 33324 33322 33376 33328
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 5000 31754 5028 33254
rect 5170 33212 5478 33221
rect 5170 33210 5176 33212
rect 5232 33210 5256 33212
rect 5312 33210 5336 33212
rect 5392 33210 5416 33212
rect 5472 33210 5478 33212
rect 5232 33158 5234 33210
rect 5414 33158 5416 33210
rect 5170 33156 5176 33158
rect 5232 33156 5256 33158
rect 5312 33156 5336 33158
rect 5392 33156 5416 33158
rect 5472 33156 5478 33158
rect 5170 33147 5478 33156
rect 5170 32124 5478 32133
rect 5170 32122 5176 32124
rect 5232 32122 5256 32124
rect 5312 32122 5336 32124
rect 5392 32122 5416 32124
rect 5472 32122 5478 32124
rect 5232 32070 5234 32122
rect 5414 32070 5416 32122
rect 5170 32068 5176 32070
rect 5232 32068 5256 32070
rect 5312 32068 5336 32070
rect 5392 32068 5416 32070
rect 5472 32068 5478 32070
rect 5170 32059 5478 32068
rect 4908 31726 5028 31754
rect 3332 25288 3384 25294
rect 3332 25230 3384 25236
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4252 25288 4304 25294
rect 4252 25230 4304 25236
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2792 24410 2820 24686
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2688 24336 2740 24342
rect 2884 24290 2912 25094
rect 2688 24278 2740 24284
rect 2700 24138 2728 24278
rect 2792 24274 2912 24290
rect 2964 24336 3016 24342
rect 2964 24278 3016 24284
rect 2780 24268 2912 24274
rect 2832 24262 2912 24268
rect 2780 24210 2832 24216
rect 2320 24132 2372 24138
rect 2320 24074 2372 24080
rect 2688 24132 2740 24138
rect 2688 24074 2740 24080
rect 2332 23866 2360 24074
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2884 23322 2912 24262
rect 2976 24206 3004 24278
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2976 21486 3004 24142
rect 3344 23798 3372 25230
rect 3884 24812 3936 24818
rect 3884 24754 3936 24760
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 3332 23792 3384 23798
rect 3332 23734 3384 23740
rect 3436 23322 3464 24074
rect 3700 23724 3752 23730
rect 3700 23666 3752 23672
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3712 22574 3740 23666
rect 3896 23526 3924 24754
rect 4080 24682 4108 25230
rect 4160 25220 4212 25226
rect 4160 25162 4212 25168
rect 4172 24818 4200 25162
rect 4160 24812 4212 24818
rect 4160 24754 4212 24760
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3068 20398 3096 21286
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3160 20466 3188 20742
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2412 20324 2464 20330
rect 2412 20266 2464 20272
rect 2424 19922 2452 20266
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1872 19514 1900 19790
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 2976 19446 3004 20198
rect 3252 19922 3280 20878
rect 3620 20534 3648 21286
rect 3712 20942 3740 22510
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2700 17134 2728 17546
rect 2976 17270 3004 18838
rect 3344 18766 3372 19722
rect 3436 18766 3464 20334
rect 3712 19854 3740 20878
rect 3700 19848 3752 19854
rect 3698 19816 3700 19825
rect 3752 19816 3754 19825
rect 3698 19751 3754 19760
rect 3896 19378 3924 23462
rect 4172 23186 4200 24754
rect 4264 23526 4292 25230
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4344 24404 4396 24410
rect 4344 24346 4396 24352
rect 4356 24070 4384 24346
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4252 23520 4304 23526
rect 4252 23462 4304 23468
rect 4264 23322 4292 23462
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3988 21554 4016 22918
rect 4356 22642 4384 24006
rect 4724 23662 4752 24686
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4344 22636 4396 22642
rect 4344 22578 4396 22584
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 20058 4016 20402
rect 4080 20398 4108 21354
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4172 20058 4200 21490
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4158 19952 4214 19961
rect 4158 19887 4214 19896
rect 4172 19854 4200 19887
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3252 17678 3280 18634
rect 3528 17814 3556 19314
rect 4264 19174 4292 19722
rect 4540 19514 4568 20402
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4632 19378 4660 23462
rect 4724 22982 4752 23598
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4908 22234 4936 31726
rect 8036 31686 8064 33322
rect 12072 33108 12124 33114
rect 12072 33050 12124 33056
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 9390 32668 9698 32677
rect 9390 32666 9396 32668
rect 9452 32666 9476 32668
rect 9532 32666 9556 32668
rect 9612 32666 9636 32668
rect 9692 32666 9698 32668
rect 9452 32614 9454 32666
rect 9634 32614 9636 32666
rect 9390 32612 9396 32614
rect 9452 32612 9476 32614
rect 9532 32612 9556 32614
rect 9612 32612 9636 32614
rect 9692 32612 9698 32614
rect 9390 32603 9698 32612
rect 8576 32292 8628 32298
rect 8576 32234 8628 32240
rect 8588 31822 8616 32234
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 8760 31952 8812 31958
rect 8760 31894 8812 31900
rect 8576 31816 8628 31822
rect 8576 31758 8628 31764
rect 8024 31680 8076 31686
rect 8024 31622 8076 31628
rect 5170 31036 5478 31045
rect 5170 31034 5176 31036
rect 5232 31034 5256 31036
rect 5312 31034 5336 31036
rect 5392 31034 5416 31036
rect 5472 31034 5478 31036
rect 5232 30982 5234 31034
rect 5414 30982 5416 31034
rect 5170 30980 5176 30982
rect 5232 30980 5256 30982
rect 5312 30980 5336 30982
rect 5392 30980 5416 30982
rect 5472 30980 5478 30982
rect 5170 30971 5478 30980
rect 5170 29948 5478 29957
rect 5170 29946 5176 29948
rect 5232 29946 5256 29948
rect 5312 29946 5336 29948
rect 5392 29946 5416 29948
rect 5472 29946 5478 29948
rect 5232 29894 5234 29946
rect 5414 29894 5416 29946
rect 5170 29892 5176 29894
rect 5232 29892 5256 29894
rect 5312 29892 5336 29894
rect 5392 29892 5416 29894
rect 5472 29892 5478 29894
rect 5170 29883 5478 29892
rect 5170 28860 5478 28869
rect 5170 28858 5176 28860
rect 5232 28858 5256 28860
rect 5312 28858 5336 28860
rect 5392 28858 5416 28860
rect 5472 28858 5478 28860
rect 5232 28806 5234 28858
rect 5414 28806 5416 28858
rect 5170 28804 5176 28806
rect 5232 28804 5256 28806
rect 5312 28804 5336 28806
rect 5392 28804 5416 28806
rect 5472 28804 5478 28806
rect 5170 28795 5478 28804
rect 8772 28014 8800 31894
rect 9864 31884 9916 31890
rect 9864 31826 9916 31832
rect 9390 31580 9698 31589
rect 9390 31578 9396 31580
rect 9452 31578 9476 31580
rect 9532 31578 9556 31580
rect 9612 31578 9636 31580
rect 9692 31578 9698 31580
rect 9452 31526 9454 31578
rect 9634 31526 9636 31578
rect 9390 31524 9396 31526
rect 9452 31524 9476 31526
rect 9532 31524 9556 31526
rect 9612 31524 9636 31526
rect 9692 31524 9698 31526
rect 9390 31515 9698 31524
rect 9876 31482 9904 31826
rect 10060 31754 10088 32166
rect 10152 31822 10180 32710
rect 10520 32434 10548 32846
rect 12084 32502 12112 33050
rect 12268 32570 12296 33322
rect 13611 33212 13919 33221
rect 13611 33210 13617 33212
rect 13673 33210 13697 33212
rect 13753 33210 13777 33212
rect 13833 33210 13857 33212
rect 13913 33210 13919 33212
rect 13673 33158 13675 33210
rect 13855 33158 13857 33210
rect 13611 33156 13617 33158
rect 13673 33156 13697 33158
rect 13753 33156 13777 33158
rect 13833 33156 13857 33158
rect 13913 33156 13919 33158
rect 13611 33147 13919 33156
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 12256 32564 12308 32570
rect 12256 32506 12308 32512
rect 13280 32502 13308 32710
rect 14292 32570 14320 33322
rect 16868 32910 16896 33322
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 14280 32564 14332 32570
rect 14280 32506 14332 32512
rect 12072 32496 12124 32502
rect 12072 32438 12124 32444
rect 13268 32496 13320 32502
rect 13268 32438 13320 32444
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 11428 32428 11480 32434
rect 11428 32370 11480 32376
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 10060 31414 10088 31690
rect 9772 31408 9824 31414
rect 9772 31350 9824 31356
rect 10048 31408 10100 31414
rect 10048 31350 10100 31356
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30938 9444 31214
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9390 30492 9698 30501
rect 9390 30490 9396 30492
rect 9452 30490 9476 30492
rect 9532 30490 9556 30492
rect 9612 30490 9636 30492
rect 9692 30490 9698 30492
rect 9452 30438 9454 30490
rect 9634 30438 9636 30490
rect 9390 30436 9396 30438
rect 9452 30436 9476 30438
rect 9532 30436 9556 30438
rect 9612 30436 9636 30438
rect 9692 30436 9698 30438
rect 9390 30427 9698 30436
rect 9036 29776 9088 29782
rect 9036 29718 9088 29724
rect 9048 29170 9076 29718
rect 9312 29504 9364 29510
rect 9312 29446 9364 29452
rect 9324 29170 9352 29446
rect 9390 29404 9698 29413
rect 9390 29402 9396 29404
rect 9452 29402 9476 29404
rect 9532 29402 9556 29404
rect 9612 29402 9636 29404
rect 9692 29402 9698 29404
rect 9452 29350 9454 29402
rect 9634 29350 9636 29402
rect 9390 29348 9396 29350
rect 9452 29348 9476 29350
rect 9532 29348 9556 29350
rect 9612 29348 9636 29350
rect 9692 29348 9698 29350
rect 9390 29339 9698 29348
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 8944 28960 8996 28966
rect 8944 28902 8996 28908
rect 8956 28218 8984 28902
rect 9048 28490 9076 29106
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 9324 28422 9352 29106
rect 9508 28626 9536 29106
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 8944 28212 8996 28218
rect 8944 28154 8996 28160
rect 8956 28014 8984 28154
rect 9140 28082 9168 28358
rect 9390 28316 9698 28325
rect 9390 28314 9396 28316
rect 9452 28314 9476 28316
rect 9532 28314 9556 28316
rect 9612 28314 9636 28316
rect 9692 28314 9698 28316
rect 9452 28262 9454 28314
rect 9634 28262 9636 28314
rect 9390 28260 9396 28262
rect 9452 28260 9476 28262
rect 9532 28260 9556 28262
rect 9612 28260 9636 28262
rect 9692 28260 9698 28262
rect 9390 28251 9698 28260
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 9784 28014 9812 31350
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 10060 30938 10088 31214
rect 10244 30938 10272 31282
rect 10336 31142 10364 32370
rect 10520 31890 10548 32370
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10508 31884 10560 31890
rect 10508 31826 10560 31832
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10048 30932 10100 30938
rect 10048 30874 10100 30880
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10336 30734 10364 31078
rect 10520 30802 10548 31826
rect 10612 31414 10640 32166
rect 11440 31822 11468 32370
rect 12348 32360 12400 32366
rect 12348 32302 12400 32308
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 11428 31816 11480 31822
rect 11428 31758 11480 31764
rect 10600 31408 10652 31414
rect 10600 31350 10652 31356
rect 10600 31272 10652 31278
rect 10600 31214 10652 31220
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 10140 30728 10192 30734
rect 10140 30670 10192 30676
rect 10324 30728 10376 30734
rect 10324 30670 10376 30676
rect 9968 29510 9996 30670
rect 10152 29578 10180 30670
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 8760 28008 8812 28014
rect 8760 27950 8812 27956
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 5170 27772 5478 27781
rect 5170 27770 5176 27772
rect 5232 27770 5256 27772
rect 5312 27770 5336 27772
rect 5392 27770 5416 27772
rect 5472 27770 5478 27772
rect 5232 27718 5234 27770
rect 5414 27718 5416 27770
rect 5170 27716 5176 27718
rect 5232 27716 5256 27718
rect 5312 27716 5336 27718
rect 5392 27716 5416 27718
rect 5472 27716 5478 27718
rect 5170 27707 5478 27716
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 8220 26994 8248 27338
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 8772 26790 8800 27950
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9036 27532 9088 27538
rect 9036 27474 9088 27480
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 5170 26684 5478 26693
rect 5170 26682 5176 26684
rect 5232 26682 5256 26684
rect 5312 26682 5336 26684
rect 5392 26682 5416 26684
rect 5472 26682 5478 26684
rect 5232 26630 5234 26682
rect 5414 26630 5416 26682
rect 5170 26628 5176 26630
rect 5232 26628 5256 26630
rect 5312 26628 5336 26630
rect 5392 26628 5416 26630
rect 5472 26628 5478 26630
rect 5170 26619 5478 26628
rect 9048 26314 9076 27474
rect 9140 27470 9168 27814
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 9140 26926 9168 26998
rect 9128 26920 9180 26926
rect 9128 26862 9180 26868
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9036 26308 9088 26314
rect 9036 26250 9088 26256
rect 9232 25838 9260 26726
rect 9324 26518 9352 27814
rect 9600 27470 9628 27814
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9390 27228 9698 27237
rect 9390 27226 9396 27228
rect 9452 27226 9476 27228
rect 9532 27226 9556 27228
rect 9612 27226 9636 27228
rect 9692 27226 9698 27228
rect 9452 27174 9454 27226
rect 9634 27174 9636 27226
rect 9390 27172 9396 27174
rect 9452 27172 9476 27174
rect 9532 27172 9556 27174
rect 9612 27172 9636 27174
rect 9692 27172 9698 27174
rect 9390 27163 9698 27172
rect 9784 26994 9812 27814
rect 10336 27062 10364 30670
rect 10612 30598 10640 31214
rect 10692 31204 10744 31210
rect 10692 31146 10744 31152
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10428 29510 10456 29582
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 10612 28966 10640 30534
rect 10704 29714 10732 31146
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10704 29578 10732 29650
rect 10692 29572 10744 29578
rect 10692 29514 10744 29520
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10704 28558 10732 29514
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11348 28218 11376 28494
rect 11336 28212 11388 28218
rect 11336 28154 11388 28160
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 11164 26450 11192 26726
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9324 25906 9352 26182
rect 9390 26140 9698 26149
rect 9390 26138 9396 26140
rect 9452 26138 9476 26140
rect 9532 26138 9556 26140
rect 9612 26138 9636 26140
rect 9692 26138 9698 26140
rect 9452 26086 9454 26138
rect 9634 26086 9636 26138
rect 9390 26084 9396 26086
rect 9452 26084 9476 26086
rect 9532 26084 9556 26086
rect 9612 26084 9636 26086
rect 9692 26084 9698 26086
rect 9390 26075 9698 26084
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9588 25832 9640 25838
rect 9864 25832 9916 25838
rect 9640 25792 9864 25820
rect 9588 25774 9640 25780
rect 9864 25774 9916 25780
rect 5170 25596 5478 25605
rect 5170 25594 5176 25596
rect 5232 25594 5256 25596
rect 5312 25594 5336 25596
rect 5392 25594 5416 25596
rect 5472 25594 5478 25596
rect 5232 25542 5234 25594
rect 5414 25542 5416 25594
rect 5170 25540 5176 25542
rect 5232 25540 5256 25542
rect 5312 25540 5336 25542
rect 5392 25540 5416 25542
rect 5472 25540 5478 25542
rect 5170 25531 5478 25540
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 4988 24676 5040 24682
rect 4988 24618 5040 24624
rect 5000 24154 5028 24618
rect 5092 24274 5120 24822
rect 5170 24508 5478 24517
rect 5170 24506 5176 24508
rect 5232 24506 5256 24508
rect 5312 24506 5336 24508
rect 5392 24506 5416 24508
rect 5472 24506 5478 24508
rect 5232 24454 5234 24506
rect 5414 24454 5416 24506
rect 5170 24452 5176 24454
rect 5232 24452 5256 24454
rect 5312 24452 5336 24454
rect 5392 24452 5416 24454
rect 5472 24452 5478 24454
rect 5170 24443 5478 24452
rect 5080 24268 5132 24274
rect 5080 24210 5132 24216
rect 5552 24206 5580 25094
rect 6840 24818 6868 25230
rect 7852 24818 7880 25230
rect 9390 25052 9698 25061
rect 9390 25050 9396 25052
rect 9452 25050 9476 25052
rect 9532 25050 9556 25052
rect 9612 25050 9636 25052
rect 9692 25050 9698 25052
rect 9452 24998 9454 25050
rect 9634 24998 9636 25050
rect 9390 24996 9396 24998
rect 9452 24996 9476 24998
rect 9532 24996 9556 24998
rect 9612 24996 9636 24998
rect 9692 24996 9698 24998
rect 9390 24987 9698 24996
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 7840 24812 7892 24818
rect 7892 24772 7972 24800
rect 7840 24754 7892 24760
rect 6840 24410 6868 24754
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 5540 24200 5592 24206
rect 5000 24126 5120 24154
rect 5540 24142 5592 24148
rect 5092 23730 5120 24126
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5828 23798 5856 24006
rect 5816 23792 5868 23798
rect 5816 23734 5868 23740
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 5092 23050 5120 23666
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 5170 23420 5478 23429
rect 5170 23418 5176 23420
rect 5232 23418 5256 23420
rect 5312 23418 5336 23420
rect 5392 23418 5416 23420
rect 5472 23418 5478 23420
rect 5232 23366 5234 23418
rect 5414 23366 5416 23418
rect 5170 23364 5176 23366
rect 5232 23364 5256 23366
rect 5312 23364 5336 23366
rect 5392 23364 5416 23366
rect 5472 23364 5478 23366
rect 5170 23355 5478 23364
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 5092 22438 5120 22986
rect 6748 22982 6776 23598
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5170 22332 5478 22341
rect 5170 22330 5176 22332
rect 5232 22330 5256 22332
rect 5312 22330 5336 22332
rect 5392 22330 5416 22332
rect 5472 22330 5478 22332
rect 5232 22278 5234 22330
rect 5414 22278 5416 22330
rect 5170 22276 5176 22278
rect 5232 22276 5256 22278
rect 5312 22276 5336 22278
rect 5392 22276 5416 22278
rect 5472 22276 5478 22278
rect 5170 22267 5478 22276
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 6748 22094 6776 22918
rect 6564 22066 6776 22094
rect 5170 21244 5478 21253
rect 5170 21242 5176 21244
rect 5232 21242 5256 21244
rect 5312 21242 5336 21244
rect 5392 21242 5416 21244
rect 5472 21242 5478 21244
rect 5232 21190 5234 21242
rect 5414 21190 5416 21242
rect 5170 21188 5176 21190
rect 5232 21188 5256 21190
rect 5312 21188 5336 21190
rect 5392 21188 5416 21190
rect 5472 21188 5478 21190
rect 5170 21179 5478 21188
rect 5170 20156 5478 20165
rect 5170 20154 5176 20156
rect 5232 20154 5256 20156
rect 5312 20154 5336 20156
rect 5392 20154 5416 20156
rect 5472 20154 5478 20156
rect 5232 20102 5234 20154
rect 5414 20102 5416 20154
rect 5170 20100 5176 20102
rect 5232 20100 5256 20102
rect 5312 20100 5336 20102
rect 5392 20100 5416 20102
rect 5472 20100 5478 20102
rect 5170 20091 5478 20100
rect 5354 19952 5410 19961
rect 5354 19887 5410 19896
rect 5368 19854 5396 19887
rect 5356 19848 5408 19854
rect 4894 19816 4950 19825
rect 5356 19790 5408 19796
rect 4894 19751 4950 19760
rect 5080 19780 5132 19786
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4908 19258 4936 19751
rect 5080 19722 5132 19728
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5092 19514 5120 19722
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5276 19258 5304 19722
rect 6564 19718 6592 22066
rect 6932 21894 6960 24210
rect 7748 24132 7800 24138
rect 7748 24074 7800 24080
rect 7760 23866 7788 24074
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7116 23322 7144 23598
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7116 22710 7144 23054
rect 7208 23050 7236 23666
rect 7380 23248 7432 23254
rect 7380 23190 7432 23196
rect 7392 23118 7420 23190
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7208 22030 7236 22986
rect 7576 22778 7604 23054
rect 7760 23050 7788 23802
rect 7944 23662 7972 24772
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8496 23798 8524 24686
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 8576 24132 8628 24138
rect 8628 24092 8708 24120
rect 8576 24074 8628 24080
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7748 23044 7800 23050
rect 7748 22986 7800 22992
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7944 22658 7972 23598
rect 8300 23588 8352 23594
rect 8300 23530 8352 23536
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 23186 8064 23462
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 8312 22710 8340 23530
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 7484 22642 7972 22658
rect 8300 22704 8352 22710
rect 8300 22646 8352 22652
rect 7472 22636 7972 22642
rect 7524 22630 7972 22636
rect 7472 22578 7524 22584
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 4908 19230 5304 19258
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2700 16794 2728 17070
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 3068 16522 3096 17478
rect 3160 16776 3188 17478
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4264 16794 4292 17138
rect 3240 16788 3292 16794
rect 3160 16748 3240 16776
rect 3240 16730 3292 16736
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2976 15094 3004 15574
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1688 14074 1716 14894
rect 2700 14414 2728 14894
rect 3068 14414 3096 16458
rect 3252 14890 3280 16730
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4264 15502 4292 16526
rect 5000 15706 5028 19230
rect 5170 19068 5478 19077
rect 5170 19066 5176 19068
rect 5232 19066 5256 19068
rect 5312 19066 5336 19068
rect 5392 19066 5416 19068
rect 5472 19066 5478 19068
rect 5232 19014 5234 19066
rect 5414 19014 5416 19066
rect 5170 19012 5176 19014
rect 5232 19012 5256 19014
rect 5312 19012 5336 19014
rect 5392 19012 5416 19014
rect 5472 19012 5478 19014
rect 5170 19003 5478 19012
rect 5170 17980 5478 17989
rect 5170 17978 5176 17980
rect 5232 17978 5256 17980
rect 5312 17978 5336 17980
rect 5392 17978 5416 17980
rect 5472 17978 5478 17980
rect 5232 17926 5234 17978
rect 5414 17926 5416 17978
rect 5170 17924 5176 17926
rect 5232 17924 5256 17926
rect 5312 17924 5336 17926
rect 5392 17924 5416 17926
rect 5472 17924 5478 17926
rect 5170 17915 5478 17924
rect 6564 17678 6592 19654
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6656 18290 6684 19314
rect 7116 18834 7144 19926
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7208 18698 7236 21830
rect 7484 21010 7512 21966
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7300 20466 7328 20878
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19786 7328 20402
rect 7392 19854 7420 20742
rect 7484 20058 7512 20946
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 20058 7696 20878
rect 8312 20602 8340 22646
rect 8404 22574 8432 23054
rect 8496 22710 8524 23734
rect 8680 23118 8708 24092
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 9324 23066 9352 24142
rect 9390 23964 9698 23973
rect 9390 23962 9396 23964
rect 9452 23962 9476 23964
rect 9532 23962 9556 23964
rect 9612 23962 9636 23964
rect 9692 23962 9698 23964
rect 9452 23910 9454 23962
rect 9634 23910 9636 23962
rect 9390 23908 9396 23910
rect 9452 23908 9476 23910
rect 9532 23908 9556 23910
rect 9612 23908 9636 23910
rect 9692 23908 9698 23910
rect 9390 23899 9698 23908
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9508 23526 9536 23598
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9508 23186 9536 23462
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9404 23112 9456 23118
rect 9324 23060 9404 23066
rect 9324 23054 9456 23060
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8404 21894 8432 22510
rect 8680 22506 8708 23054
rect 9324 23038 9444 23054
rect 9772 23044 9824 23050
rect 9324 22778 9352 23038
rect 9772 22986 9824 22992
rect 9390 22876 9698 22885
rect 9390 22874 9396 22876
rect 9452 22874 9476 22876
rect 9532 22874 9556 22876
rect 9612 22874 9636 22876
rect 9692 22874 9698 22876
rect 9452 22822 9454 22874
rect 9634 22822 9636 22874
rect 9390 22820 9396 22822
rect 9452 22820 9476 22822
rect 9532 22820 9556 22822
rect 9612 22820 9636 22822
rect 9692 22820 9698 22822
rect 9390 22811 9698 22820
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 8668 22500 8720 22506
rect 8668 22442 8720 22448
rect 9220 22432 9272 22438
rect 9220 22374 9272 22380
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 5170 16892 5478 16901
rect 5170 16890 5176 16892
rect 5232 16890 5256 16892
rect 5312 16890 5336 16892
rect 5392 16890 5416 16892
rect 5472 16890 5478 16892
rect 5232 16838 5234 16890
rect 5414 16838 5416 16890
rect 5170 16836 5176 16838
rect 5232 16836 5256 16838
rect 5312 16836 5336 16838
rect 5392 16836 5416 16838
rect 5472 16836 5478 16838
rect 5170 16827 5478 16836
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 5092 15570 5120 16458
rect 6380 16454 6408 17614
rect 6564 17218 6592 17614
rect 6472 17190 6592 17218
rect 6472 16590 6500 17190
rect 6656 17134 6684 18226
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6748 17882 6776 18158
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6932 17338 6960 18158
rect 7116 17542 7144 18294
rect 7300 18154 7328 19722
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6644 17128 6696 17134
rect 6564 17088 6644 17116
rect 6564 16794 6592 17088
rect 6644 17070 6696 17076
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6472 16250 6500 16526
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 5170 15804 5478 15813
rect 5170 15802 5176 15804
rect 5232 15802 5256 15804
rect 5312 15802 5336 15804
rect 5392 15802 5416 15804
rect 5472 15802 5478 15804
rect 5232 15750 5234 15802
rect 5414 15750 5416 15802
rect 5170 15748 5176 15750
rect 5232 15748 5256 15750
rect 5312 15748 5336 15750
rect 5392 15748 5416 15750
rect 5472 15748 5478 15750
rect 5170 15739 5478 15748
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2976 14074 3004 14282
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3068 13938 3096 14350
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 2424 12918 2452 13126
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 3068 12442 3096 12854
rect 3160 12782 3188 13126
rect 3620 12782 3648 13874
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3712 12730 3740 14010
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13530 4200 13806
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4264 13462 4292 14758
rect 4448 14006 4476 15302
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3896 12986 3924 13262
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3988 12986 4016 13194
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3160 12322 3188 12718
rect 3620 12458 3648 12718
rect 3712 12702 3924 12730
rect 3620 12430 3832 12458
rect 3068 12294 3188 12322
rect 3068 12238 3096 12294
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2976 10742 3004 12106
rect 3804 11082 3832 12430
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10062 2820 10406
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2148 9178 2176 9862
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2516 9110 2544 9590
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2608 8498 2636 9318
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2700 8634 2728 9114
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2792 8498 2820 9998
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 8906 2912 9318
rect 2976 9042 3004 10678
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 3068 10266 3096 10610
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3068 9518 3096 10202
rect 3344 9926 3372 10542
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3528 9602 3556 10474
rect 3160 9586 3556 9602
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3148 9580 3556 9586
rect 3200 9574 3556 9580
rect 3148 9522 3200 9528
rect 3528 9518 3556 9574
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 7002 2636 7142
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2884 6458 2912 6666
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2976 6322 3004 8978
rect 3068 8634 3096 9454
rect 3620 8634 3648 9590
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3712 8498 3740 9046
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3804 7410 3832 11018
rect 3896 10674 3924 12702
rect 4080 12238 4108 13194
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4160 11008 4212 11014
rect 4264 10996 4292 13398
rect 4540 12850 4568 14962
rect 5092 13870 5120 15506
rect 5552 15434 5580 16186
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5736 15162 5764 16118
rect 6472 15978 6500 16186
rect 6564 16114 6592 16390
rect 6656 16114 6684 16662
rect 6748 16250 6776 17138
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6564 15570 6592 16050
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6460 15496 6512 15502
rect 6656 15450 6684 16050
rect 6748 15502 6776 16186
rect 6840 16182 6868 17138
rect 7116 16674 7144 17478
rect 7484 17202 7512 19994
rect 7760 19990 7788 20470
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 7748 19984 7800 19990
rect 7748 19926 7800 19932
rect 7852 19718 7880 20266
rect 8036 19854 8064 20402
rect 8496 19854 8524 20402
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18970 7696 19314
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7196 16720 7248 16726
rect 7116 16668 7196 16674
rect 7116 16662 7248 16668
rect 7116 16646 7236 16662
rect 7288 16652 7340 16658
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 7116 16046 7144 16646
rect 7288 16594 7340 16600
rect 7300 16182 7328 16594
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 6512 15444 6684 15450
rect 6460 15438 6684 15444
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 6104 14822 6132 15438
rect 6472 15422 6684 15438
rect 7208 15434 7236 16050
rect 7196 15428 7248 15434
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 5170 14716 5478 14725
rect 5170 14714 5176 14716
rect 5232 14714 5256 14716
rect 5312 14714 5336 14716
rect 5392 14714 5416 14716
rect 5472 14714 5478 14716
rect 5232 14662 5234 14714
rect 5414 14662 5416 14714
rect 5170 14660 5176 14662
rect 5232 14660 5256 14662
rect 5312 14660 5336 14662
rect 5392 14660 5416 14662
rect 5472 14660 5478 14662
rect 5170 14651 5478 14660
rect 6380 14414 6408 15098
rect 6472 15094 6500 15422
rect 7196 15370 7248 15376
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6460 15088 6512 15094
rect 6460 15030 6512 15036
rect 6840 14618 6868 15302
rect 7208 14618 7236 15370
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 14006 6408 14350
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6656 14006 6684 14282
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13326 5120 13806
rect 5170 13628 5478 13637
rect 5170 13626 5176 13628
rect 5232 13626 5256 13628
rect 5312 13626 5336 13628
rect 5392 13626 5416 13628
rect 5472 13626 5478 13628
rect 5232 13574 5234 13626
rect 5414 13574 5416 13626
rect 5170 13572 5176 13574
rect 5232 13572 5256 13574
rect 5312 13572 5336 13574
rect 5392 13572 5416 13574
rect 5472 13572 5478 13574
rect 5170 13563 5478 13572
rect 5552 13530 5580 13874
rect 6840 13734 6868 14554
rect 7208 14414 7236 14554
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7484 14278 7512 16050
rect 7760 15910 7788 17138
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15706 7788 15846
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7852 14346 7880 19654
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8128 18698 8156 19110
rect 8496 18902 8524 19790
rect 8956 19786 8984 20334
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8956 19378 8984 19722
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 8128 18290 8156 18634
rect 8956 18426 8984 19314
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 17066 8156 18226
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4540 11354 4568 12786
rect 5170 12540 5478 12549
rect 5170 12538 5176 12540
rect 5232 12538 5256 12540
rect 5312 12538 5336 12540
rect 5392 12538 5416 12540
rect 5472 12538 5478 12540
rect 5232 12486 5234 12538
rect 5414 12486 5416 12538
rect 5170 12484 5176 12486
rect 5232 12484 5256 12486
rect 5312 12484 5336 12486
rect 5392 12484 5416 12486
rect 5472 12484 5478 12486
rect 5170 12475 5478 12484
rect 6932 12434 6960 14214
rect 7484 14006 7512 14214
rect 7944 14074 7972 14350
rect 8128 14278 8156 17002
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8220 16726 8248 16934
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 9048 15026 9076 21830
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18834 9168 19110
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9232 17270 9260 22374
rect 9324 22030 9352 22714
rect 9784 22710 9812 22986
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9876 22234 9904 23190
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9390 21788 9698 21797
rect 9390 21786 9396 21788
rect 9452 21786 9476 21788
rect 9532 21786 9556 21788
rect 9612 21786 9636 21788
rect 9692 21786 9698 21788
rect 9452 21734 9454 21786
rect 9634 21734 9636 21786
rect 9390 21732 9396 21734
rect 9452 21732 9476 21734
rect 9532 21732 9556 21734
rect 9612 21732 9636 21734
rect 9692 21732 9698 21734
rect 9390 21723 9698 21732
rect 9390 20700 9698 20709
rect 9390 20698 9396 20700
rect 9452 20698 9476 20700
rect 9532 20698 9556 20700
rect 9612 20698 9636 20700
rect 9692 20698 9698 20700
rect 9452 20646 9454 20698
rect 9634 20646 9636 20698
rect 9390 20644 9396 20646
rect 9452 20644 9476 20646
rect 9532 20644 9556 20646
rect 9612 20644 9636 20646
rect 9692 20644 9698 20646
rect 9390 20635 9698 20644
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9390 19612 9698 19621
rect 9390 19610 9396 19612
rect 9452 19610 9476 19612
rect 9532 19610 9556 19612
rect 9612 19610 9636 19612
rect 9692 19610 9698 19612
rect 9452 19558 9454 19610
rect 9634 19558 9636 19610
rect 9390 19556 9396 19558
rect 9452 19556 9476 19558
rect 9532 19556 9556 19558
rect 9612 19556 9636 19558
rect 9692 19556 9698 19558
rect 9390 19547 9698 19556
rect 9784 19378 9812 19722
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9390 18524 9698 18533
rect 9390 18522 9396 18524
rect 9452 18522 9476 18524
rect 9532 18522 9556 18524
rect 9612 18522 9636 18524
rect 9692 18522 9698 18524
rect 9452 18470 9454 18522
rect 9634 18470 9636 18522
rect 9390 18468 9396 18470
rect 9452 18468 9476 18470
rect 9532 18468 9556 18470
rect 9612 18468 9636 18470
rect 9692 18468 9698 18470
rect 9390 18459 9698 18468
rect 9968 17542 9996 19790
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9390 17436 9698 17445
rect 9390 17434 9396 17436
rect 9452 17434 9476 17436
rect 9532 17434 9556 17436
rect 9612 17434 9636 17436
rect 9692 17434 9698 17436
rect 9452 17382 9454 17434
rect 9634 17382 9636 17434
rect 9390 17380 9396 17382
rect 9452 17380 9476 17382
rect 9532 17380 9556 17382
rect 9612 17380 9636 17382
rect 9692 17380 9698 17382
rect 9390 17371 9698 17380
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9390 16348 9698 16357
rect 9390 16346 9396 16348
rect 9452 16346 9476 16348
rect 9532 16346 9556 16348
rect 9612 16346 9636 16348
rect 9692 16346 9698 16348
rect 9452 16294 9454 16346
rect 9634 16294 9636 16346
rect 9390 16292 9396 16294
rect 9452 16292 9476 16294
rect 9532 16292 9556 16294
rect 9612 16292 9636 16294
rect 9692 16292 9698 16294
rect 9390 16283 9698 16292
rect 9390 15260 9698 15269
rect 9390 15258 9396 15260
rect 9452 15258 9476 15260
rect 9532 15258 9556 15260
rect 9612 15258 9636 15260
rect 9692 15258 9698 15260
rect 9452 15206 9454 15258
rect 9634 15206 9636 15258
rect 9390 15204 9396 15206
rect 9452 15204 9476 15206
rect 9532 15204 9556 15206
rect 9612 15204 9636 15206
rect 9692 15204 9698 15206
rect 9390 15195 9698 15204
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 8944 14952 8996 14958
rect 8944 14894 8996 14900
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 6932 12406 7052 12434
rect 5170 11452 5478 11461
rect 5170 11450 5176 11452
rect 5232 11450 5256 11452
rect 5312 11450 5336 11452
rect 5392 11450 5416 11452
rect 5472 11450 5478 11452
rect 5232 11398 5234 11450
rect 5414 11398 5416 11450
rect 5170 11396 5176 11398
rect 5232 11396 5256 11398
rect 5312 11396 5336 11398
rect 5392 11396 5416 11398
rect 5472 11396 5478 11398
rect 5170 11387 5478 11396
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4212 10968 4292 10996
rect 4160 10950 4212 10956
rect 4264 10674 4292 10968
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 3896 10130 3924 10610
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3988 9654 4016 9930
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4080 9518 4108 10202
rect 4264 10130 4292 10610
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4356 10062 4384 10950
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9722 4384 9998
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4356 8974 4384 9658
rect 4540 9586 4568 11086
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5170 10364 5478 10373
rect 5170 10362 5176 10364
rect 5232 10362 5256 10364
rect 5312 10362 5336 10364
rect 5392 10362 5416 10364
rect 5472 10362 5478 10364
rect 5232 10310 5234 10362
rect 5414 10310 5416 10362
rect 5170 10308 5176 10310
rect 5232 10308 5256 10310
rect 5312 10308 5336 10310
rect 5392 10308 5416 10310
rect 5472 10308 5478 10310
rect 5170 10299 5478 10308
rect 5644 9994 5672 11018
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10742 6960 10950
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 5170 9276 5478 9285
rect 5170 9274 5176 9276
rect 5232 9274 5256 9276
rect 5312 9274 5336 9276
rect 5392 9274 5416 9276
rect 5472 9274 5478 9276
rect 5232 9222 5234 9274
rect 5414 9222 5416 9274
rect 5170 9220 5176 9222
rect 5232 9220 5256 9222
rect 5312 9220 5336 9222
rect 5392 9220 5416 9222
rect 5472 9220 5478 9222
rect 5170 9211 5478 9220
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3804 6866 3832 7346
rect 4356 6866 4384 8774
rect 5170 8188 5478 8197
rect 5170 8186 5176 8188
rect 5232 8186 5256 8188
rect 5312 8186 5336 8188
rect 5392 8186 5416 8188
rect 5472 8186 5478 8188
rect 5232 8134 5234 8186
rect 5414 8134 5416 8186
rect 5170 8132 5176 8134
rect 5232 8132 5256 8134
rect 5312 8132 5336 8134
rect 5392 8132 5416 8134
rect 5472 8132 5478 8134
rect 5170 8123 5478 8132
rect 5644 7478 5672 9930
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5170 7100 5478 7109
rect 5170 7098 5176 7100
rect 5232 7098 5256 7100
rect 5312 7098 5336 7100
rect 5392 7098 5416 7100
rect 5472 7098 5478 7100
rect 5232 7046 5234 7098
rect 5414 7046 5416 7098
rect 5170 7044 5176 7046
rect 5232 7044 5256 7046
rect 5312 7044 5336 7046
rect 5392 7044 5416 7046
rect 5472 7044 5478 7046
rect 5170 7035 5478 7044
rect 5644 6882 5672 7414
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 5080 6860 5132 6866
rect 5644 6854 5764 6882
rect 5080 6802 5132 6808
rect 3160 6322 3188 6802
rect 3804 6390 3832 6802
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2976 5302 3004 6258
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4080 5574 4108 6190
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 4080 5234 4108 5510
rect 4724 5302 4752 5578
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 5092 4690 5120 6802
rect 5736 6798 5764 6854
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5170 6012 5478 6021
rect 5170 6010 5176 6012
rect 5232 6010 5256 6012
rect 5312 6010 5336 6012
rect 5392 6010 5416 6012
rect 5472 6010 5478 6012
rect 5232 5958 5234 6010
rect 5414 5958 5416 6010
rect 5170 5956 5176 5958
rect 5232 5956 5256 5958
rect 5312 5956 5336 5958
rect 5392 5956 5416 5958
rect 5472 5956 5478 5958
rect 5170 5947 5478 5956
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5644 5370 5672 5714
rect 6104 5574 6132 6190
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6104 5370 6132 5510
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 5644 5166 5672 5306
rect 6564 5166 6592 10542
rect 6748 10266 6776 10678
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9586 6868 9998
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9042 6868 9522
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6458 6960 6598
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7024 6390 7052 12406
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10130 7236 11086
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10742 7420 10950
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7484 10062 7512 13126
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 10742 7604 12582
rect 8128 10810 8156 14214
rect 8220 14074 8248 14282
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8312 13462 8340 14486
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 10266 8156 10406
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7484 9654 7512 9998
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7392 7478 7420 7754
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 5170 4924 5478 4933
rect 5170 4922 5176 4924
rect 5232 4922 5256 4924
rect 5312 4922 5336 4924
rect 5392 4922 5416 4924
rect 5472 4922 5478 4924
rect 5232 4870 5234 4922
rect 5414 4870 5416 4922
rect 5170 4868 5176 4870
rect 5232 4868 5256 4870
rect 5312 4868 5336 4870
rect 5392 4868 5416 4870
rect 5472 4868 5478 4870
rect 5170 4859 5478 4868
rect 7208 4690 7236 5034
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7484 4622 7512 9590
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7484 4214 7512 4558
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 5170 3836 5478 3845
rect 5170 3834 5176 3836
rect 5232 3834 5256 3836
rect 5312 3834 5336 3836
rect 5392 3834 5416 3836
rect 5472 3834 5478 3836
rect 5232 3782 5234 3834
rect 5414 3782 5416 3834
rect 5170 3780 5176 3782
rect 5232 3780 5256 3782
rect 5312 3780 5336 3782
rect 5392 3780 5416 3782
rect 5472 3780 5478 3782
rect 5170 3771 5478 3780
rect 5170 2748 5478 2757
rect 5170 2746 5176 2748
rect 5232 2746 5256 2748
rect 5312 2746 5336 2748
rect 5392 2746 5416 2748
rect 5472 2746 5478 2748
rect 5232 2694 5234 2746
rect 5414 2694 5416 2746
rect 5170 2692 5176 2694
rect 5232 2692 5256 2694
rect 5312 2692 5336 2694
rect 5392 2692 5416 2694
rect 5472 2692 5478 2694
rect 5170 2683 5478 2692
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 1228 800 1256 2314
rect 2516 800 2544 2314
rect 3804 800 3832 2314
rect 5092 800 5120 2314
rect 6380 800 6408 2382
rect 7576 2378 7604 10202
rect 8128 9926 8156 10202
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8208 8288 8260 8294
rect 8312 8242 8340 13262
rect 8260 8236 8340 8242
rect 8208 8230 8340 8236
rect 8220 8214 8340 8230
rect 8220 7886 8248 8214
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 5030 8156 7754
rect 8220 5642 8248 7822
rect 8404 7410 8432 13874
rect 8496 13190 8524 14486
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8680 12918 8708 13194
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8588 9722 8616 10678
rect 8680 10266 8708 10746
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8956 10198 8984 14894
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 10962 9076 13126
rect 9140 12986 9168 13330
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9324 12918 9352 14486
rect 9784 14346 9812 14962
rect 9876 14958 9904 17138
rect 9968 16590 9996 17478
rect 10060 17202 10088 23122
rect 10244 22234 10272 23258
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10336 22778 10364 22918
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10428 22642 10456 22918
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10336 20942 10364 22374
rect 10428 22094 10456 22578
rect 10428 22066 10548 22094
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10244 20466 10272 20742
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10244 19786 10272 20402
rect 10336 20398 10364 20878
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10336 19854 10364 20334
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10152 17134 10180 19178
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10244 18766 10272 19110
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16590 10088 16934
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9390 14172 9698 14181
rect 9390 14170 9396 14172
rect 9452 14170 9476 14172
rect 9532 14170 9556 14172
rect 9612 14170 9636 14172
rect 9692 14170 9698 14172
rect 9452 14118 9454 14170
rect 9634 14118 9636 14170
rect 9390 14116 9396 14118
rect 9452 14116 9476 14118
rect 9532 14116 9556 14118
rect 9612 14116 9636 14118
rect 9692 14116 9698 14118
rect 9390 14107 9698 14116
rect 9956 14068 10008 14074
rect 10152 14056 10180 17070
rect 10244 14278 10272 18022
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10336 15026 10364 17274
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16114 10456 16390
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10008 14028 10180 14056
rect 9956 14010 10008 14016
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9876 13258 9904 13806
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9390 13084 9698 13093
rect 9390 13082 9396 13084
rect 9452 13082 9476 13084
rect 9532 13082 9556 13084
rect 9612 13082 9636 13084
rect 9692 13082 9698 13084
rect 9452 13030 9454 13082
rect 9634 13030 9636 13082
rect 9390 13028 9396 13030
rect 9452 13028 9476 13030
rect 9532 13028 9556 13030
rect 9612 13028 9636 13030
rect 9692 13028 9698 13030
rect 9390 13019 9698 13028
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9324 11082 9352 12854
rect 9390 11996 9698 12005
rect 9390 11994 9396 11996
rect 9452 11994 9476 11996
rect 9532 11994 9556 11996
rect 9612 11994 9636 11996
rect 9692 11994 9698 11996
rect 9452 11942 9454 11994
rect 9634 11942 9636 11994
rect 9390 11940 9396 11942
rect 9452 11940 9476 11942
rect 9532 11940 9556 11942
rect 9612 11940 9636 11942
rect 9692 11940 9698 11942
rect 9390 11931 9698 11940
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9772 11008 9824 11014
rect 9048 10934 9352 10962
rect 9772 10950 9824 10956
rect 9324 10724 9352 10934
rect 9390 10908 9698 10917
rect 9390 10906 9396 10908
rect 9452 10906 9476 10908
rect 9532 10906 9556 10908
rect 9612 10906 9636 10908
rect 9692 10906 9698 10908
rect 9452 10854 9454 10906
rect 9634 10854 9636 10906
rect 9390 10852 9396 10854
rect 9452 10852 9476 10854
rect 9532 10852 9556 10854
rect 9612 10852 9636 10854
rect 9692 10852 9698 10854
rect 9390 10843 9698 10852
rect 9784 10810 9812 10950
rect 9968 10810 9996 14010
rect 10520 13530 10548 22066
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 20942 10732 21830
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10704 19786 10732 20878
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10796 19378 10824 22714
rect 11716 22642 11744 31894
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11808 28626 11836 29106
rect 11796 28620 11848 28626
rect 11796 28562 11848 28568
rect 11900 24206 11928 32166
rect 12360 31822 12388 32302
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12636 29510 12664 31282
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12912 29646 12940 29990
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12624 29504 12676 29510
rect 12624 29446 12676 29452
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12636 29170 12664 29446
rect 12820 29170 12848 29446
rect 12912 29306 12940 29582
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12624 29164 12676 29170
rect 12624 29106 12676 29112
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12544 28082 12572 28562
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12360 25974 12388 27338
rect 12452 26994 12480 27950
rect 12544 27538 12572 28018
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12636 27402 12664 29106
rect 12820 28558 12848 29106
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 13096 28422 13124 28494
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 13084 28416 13136 28422
rect 13084 28358 13136 28364
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12636 27062 12664 27338
rect 12912 27130 12940 28358
rect 13096 28218 13124 28358
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12624 27056 12676 27062
rect 12624 26998 12676 27004
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 26738 12480 26930
rect 12624 26784 12676 26790
rect 12452 26710 12572 26738
rect 12624 26726 12676 26732
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12452 25974 12480 26522
rect 12544 26314 12572 26710
rect 12636 26382 12664 26726
rect 12912 26586 12940 27066
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12808 26444 12860 26450
rect 12808 26386 12860 26392
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12544 26042 12572 26250
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12268 25294 12296 25842
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12728 25294 12756 25638
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12268 24954 12296 25230
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12820 24818 12848 26386
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 25362 13124 25638
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 11900 23050 11928 24142
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 23662 12296 24074
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 22234 11744 22578
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 10980 22094 11008 22170
rect 10980 22066 11100 22094
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10980 20806 11008 21422
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 19922 11008 20742
rect 11072 20466 11100 22066
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 11532 19310 11560 19654
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10704 18766 10732 19110
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 11072 18290 11100 19246
rect 11624 19122 11652 22034
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21622 11744 21898
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11808 21554 11836 22510
rect 11980 22500 12032 22506
rect 11980 22442 12032 22448
rect 11992 21554 12020 22442
rect 12084 22098 12112 23054
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11532 19094 11652 19122
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11532 17746 11560 19094
rect 11808 18290 11836 21490
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 16726 11008 17478
rect 11532 17134 11560 17682
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10980 16114 11008 16662
rect 11072 16590 11100 16730
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11072 15706 11100 16526
rect 11164 16522 11192 16934
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 16114 11192 16458
rect 11532 16182 11560 17070
rect 12084 16590 12112 18294
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12176 17610 12204 18158
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12268 17354 12296 23598
rect 12452 22642 12480 24142
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12636 22642 12664 24006
rect 12912 23730 12940 24006
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13188 23662 13216 32166
rect 13611 32124 13919 32133
rect 13611 32122 13617 32124
rect 13673 32122 13697 32124
rect 13753 32122 13777 32124
rect 13833 32122 13857 32124
rect 13913 32122 13919 32124
rect 13673 32070 13675 32122
rect 13855 32070 13857 32122
rect 13611 32068 13617 32070
rect 13673 32068 13697 32070
rect 13753 32068 13777 32070
rect 13833 32068 13857 32070
rect 13913 32068 13919 32070
rect 13611 32059 13919 32068
rect 16120 32020 16172 32026
rect 16120 31962 16172 31968
rect 16132 31822 16160 31962
rect 14004 31816 14056 31822
rect 14004 31758 14056 31764
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13280 30938 13308 31214
rect 13611 31036 13919 31045
rect 13611 31034 13617 31036
rect 13673 31034 13697 31036
rect 13753 31034 13777 31036
rect 13833 31034 13857 31036
rect 13913 31034 13919 31036
rect 13673 30982 13675 31034
rect 13855 30982 13857 31034
rect 13611 30980 13617 30982
rect 13673 30980 13697 30982
rect 13753 30980 13777 30982
rect 13833 30980 13857 30982
rect 13913 30980 13919 30982
rect 13611 30971 13919 30980
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 14016 30598 14044 31758
rect 14292 31482 14320 31758
rect 14280 31476 14332 31482
rect 14280 31418 14332 31424
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 14108 30734 14136 31282
rect 14660 31278 14688 31758
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15580 31414 15608 31690
rect 15752 31680 15804 31686
rect 15752 31622 15804 31628
rect 15568 31408 15620 31414
rect 15568 31350 15620 31356
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14292 30258 14320 31078
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 13611 29948 13919 29957
rect 13611 29946 13617 29948
rect 13673 29946 13697 29948
rect 13753 29946 13777 29948
rect 13833 29946 13857 29948
rect 13913 29946 13919 29948
rect 13673 29894 13675 29946
rect 13855 29894 13857 29946
rect 13611 29892 13617 29894
rect 13673 29892 13697 29894
rect 13753 29892 13777 29894
rect 13833 29892 13857 29894
rect 13913 29892 13919 29894
rect 13611 29883 13919 29892
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13464 28694 13492 29106
rect 13611 28860 13919 28869
rect 13611 28858 13617 28860
rect 13673 28858 13697 28860
rect 13753 28858 13777 28860
rect 13833 28858 13857 28860
rect 13913 28858 13919 28860
rect 13673 28806 13675 28858
rect 13855 28806 13857 28858
rect 13611 28804 13617 28806
rect 13673 28804 13697 28806
rect 13753 28804 13777 28806
rect 13833 28804 13857 28806
rect 13913 28804 13919 28806
rect 13611 28795 13919 28804
rect 13452 28688 13504 28694
rect 13452 28630 13504 28636
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 13280 28082 13308 28494
rect 13464 28490 13492 28630
rect 13452 28484 13504 28490
rect 13452 28426 13504 28432
rect 13464 28150 13492 28426
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 14292 28082 14320 29514
rect 14568 29306 14596 30670
rect 14556 29300 14608 29306
rect 14556 29242 14608 29248
rect 14660 29186 14688 31214
rect 14844 30870 14872 31282
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14844 29850 14872 30806
rect 15488 30734 15516 31282
rect 15764 31278 15792 31622
rect 16132 31482 16160 31758
rect 16120 31476 16172 31482
rect 16120 31418 16172 31424
rect 15752 31272 15804 31278
rect 15752 31214 15804 31220
rect 15764 30802 15792 31214
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 14936 30258 14964 30670
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14936 29306 14964 30194
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14924 29300 14976 29306
rect 14924 29242 14976 29248
rect 14568 29158 14688 29186
rect 14568 28558 14596 29158
rect 15028 29102 15056 29582
rect 15108 29572 15160 29578
rect 15108 29514 15160 29520
rect 15120 29238 15148 29514
rect 15108 29232 15160 29238
rect 15108 29174 15160 29180
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 15028 28626 15056 29038
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 13611 27772 13919 27781
rect 13611 27770 13617 27772
rect 13673 27770 13697 27772
rect 13753 27770 13777 27772
rect 13833 27770 13857 27772
rect 13913 27770 13919 27772
rect 13673 27718 13675 27770
rect 13855 27718 13857 27770
rect 13611 27716 13617 27718
rect 13673 27716 13697 27718
rect 13753 27716 13777 27718
rect 13833 27716 13857 27718
rect 13913 27716 13919 27718
rect 13611 27707 13919 27716
rect 14016 27538 14044 28018
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13740 26994 13768 27338
rect 13832 27062 13860 27406
rect 14292 27062 14320 28018
rect 14568 28014 14596 28494
rect 15028 28150 15056 28562
rect 15120 28558 15148 29174
rect 15568 29164 15620 29170
rect 15568 29106 15620 29112
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15396 28218 15424 28494
rect 15384 28212 15436 28218
rect 15384 28154 15436 28160
rect 15016 28144 15068 28150
rect 15016 28086 15068 28092
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 14280 27056 14332 27062
rect 14280 26998 14332 27004
rect 13452 26988 13504 26994
rect 13452 26930 13504 26936
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 13360 26580 13412 26586
rect 13360 26522 13412 26528
rect 13372 25974 13400 26522
rect 13464 26450 13492 26930
rect 13611 26684 13919 26693
rect 13611 26682 13617 26684
rect 13673 26682 13697 26684
rect 13753 26682 13777 26684
rect 13833 26682 13857 26684
rect 13913 26682 13919 26684
rect 13673 26630 13675 26682
rect 13855 26630 13857 26682
rect 13611 26628 13617 26630
rect 13673 26628 13697 26630
rect 13753 26628 13777 26630
rect 13833 26628 13857 26630
rect 13913 26628 13919 26630
rect 13611 26619 13919 26628
rect 13452 26444 13504 26450
rect 13452 26386 13504 26392
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13360 25968 13412 25974
rect 13360 25910 13412 25916
rect 13464 25906 13492 26250
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 14464 25764 14516 25770
rect 14464 25706 14516 25712
rect 13611 25596 13919 25605
rect 13611 25594 13617 25596
rect 13673 25594 13697 25596
rect 13753 25594 13777 25596
rect 13833 25594 13857 25596
rect 13913 25594 13919 25596
rect 13673 25542 13675 25594
rect 13855 25542 13857 25594
rect 13611 25540 13617 25542
rect 13673 25540 13697 25542
rect 13753 25540 13777 25542
rect 13833 25540 13857 25542
rect 13913 25540 13919 25542
rect 13611 25531 13919 25540
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13464 24274 13492 25094
rect 13611 24508 13919 24517
rect 13611 24506 13617 24508
rect 13673 24506 13697 24508
rect 13753 24506 13777 24508
rect 13833 24506 13857 24508
rect 13913 24506 13919 24508
rect 13673 24454 13675 24506
rect 13855 24454 13857 24506
rect 13611 24452 13617 24454
rect 13673 24452 13697 24454
rect 13753 24452 13777 24454
rect 13833 24452 13857 24454
rect 13913 24452 13919 24454
rect 13611 24443 13919 24452
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13280 23730 13308 24142
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12912 22030 12940 22442
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 22030 13032 22374
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12728 21690 12756 21966
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12360 18698 12388 21490
rect 12912 21146 12940 21966
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18766 12480 19314
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12360 18358 12388 18634
rect 12452 18426 12480 18702
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12176 17326 12296 17354
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 14346 10732 14962
rect 11072 14414 11100 15642
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10520 12714 10548 13466
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9404 10736 9456 10742
rect 9324 10696 9404 10724
rect 9404 10678 9456 10684
rect 10060 10198 10088 10746
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9390 9820 9698 9829
rect 9390 9818 9396 9820
rect 9452 9818 9476 9820
rect 9532 9818 9556 9820
rect 9612 9818 9636 9820
rect 9692 9818 9698 9820
rect 9452 9766 9454 9818
rect 9634 9766 9636 9818
rect 9390 9764 9396 9766
rect 9452 9764 9476 9766
rect 9532 9764 9556 9766
rect 9612 9764 9636 9766
rect 9692 9764 9698 9766
rect 9390 9755 9698 9764
rect 10152 9722 10180 10406
rect 10336 10130 10364 11086
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 9390 8732 9698 8741
rect 9390 8730 9396 8732
rect 9452 8730 9476 8732
rect 9532 8730 9556 8732
rect 9612 8730 9636 8732
rect 9692 8730 9698 8732
rect 9452 8678 9454 8730
rect 9634 8678 9636 8730
rect 9390 8676 9396 8678
rect 9452 8676 9476 8678
rect 9532 8676 9556 8678
rect 9612 8676 9636 8678
rect 9692 8676 9698 8678
rect 9390 8667 9698 8676
rect 9390 7644 9698 7653
rect 9390 7642 9396 7644
rect 9452 7642 9476 7644
rect 9532 7642 9556 7644
rect 9612 7642 9636 7644
rect 9692 7642 9698 7644
rect 9452 7590 9454 7642
rect 9634 7590 9636 7642
rect 9390 7588 9396 7590
rect 9452 7588 9476 7590
rect 9532 7588 9556 7590
rect 9612 7588 9636 7590
rect 9692 7588 9698 7590
rect 9390 7579 9698 7588
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6866 8340 7142
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8312 6662 8340 6802
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 3738 7972 4150
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8128 3534 8156 4966
rect 8220 3602 8248 5578
rect 8956 4690 8984 7346
rect 9390 6556 9698 6565
rect 9390 6554 9396 6556
rect 9452 6554 9476 6556
rect 9532 6554 9556 6556
rect 9612 6554 9636 6556
rect 9692 6554 9698 6556
rect 9452 6502 9454 6554
rect 9634 6502 9636 6554
rect 9390 6500 9396 6502
rect 9452 6500 9476 6502
rect 9532 6500 9556 6502
rect 9612 6500 9636 6502
rect 9692 6500 9698 6502
rect 9390 6491 9698 6500
rect 9390 5468 9698 5477
rect 9390 5466 9396 5468
rect 9452 5466 9476 5468
rect 9532 5466 9556 5468
rect 9612 5466 9636 5468
rect 9692 5466 9698 5468
rect 9452 5414 9454 5466
rect 9634 5414 9636 5466
rect 9390 5412 9396 5414
rect 9452 5412 9476 5414
rect 9532 5412 9556 5414
rect 9612 5412 9636 5414
rect 9692 5412 9698 5414
rect 9390 5403 9698 5412
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 4146 8984 4626
rect 9324 4282 9352 5238
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9390 4380 9698 4389
rect 9390 4378 9396 4380
rect 9452 4378 9476 4380
rect 9532 4378 9556 4380
rect 9612 4378 9636 4380
rect 9692 4378 9698 4380
rect 9452 4326 9454 4378
rect 9634 4326 9636 4378
rect 9390 4324 9396 4326
rect 9452 4324 9476 4326
rect 9532 4324 9556 4326
rect 9612 4324 9636 4326
rect 9692 4324 9698 4326
rect 9390 4315 9698 4324
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9784 4146 9812 4422
rect 9876 4282 9904 5170
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4282 9996 4966
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 9390 3292 9698 3301
rect 9390 3290 9396 3292
rect 9452 3290 9476 3292
rect 9532 3290 9556 3292
rect 9612 3290 9636 3292
rect 9692 3290 9698 3292
rect 9452 3238 9454 3290
rect 9634 3238 9636 3290
rect 9390 3236 9396 3238
rect 9452 3236 9476 3238
rect 9532 3236 9556 3238
rect 9612 3236 9636 3238
rect 9692 3236 9698 3238
rect 9390 3227 9698 3236
rect 10152 2582 10180 9658
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 10244 7478 10272 7754
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10520 6882 10548 7482
rect 10428 6854 10548 6882
rect 10704 6866 10732 14282
rect 11072 14006 11100 14350
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11164 13394 11192 14894
rect 11992 14006 12020 15030
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 11072 8974 11100 11086
rect 11256 11014 11284 11290
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 7342 11100 8910
rect 11256 7342 11284 10950
rect 11532 9994 11560 13330
rect 11808 13326 11836 13806
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11808 12986 11836 13262
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11992 11150 12020 13942
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11808 9586 11836 9930
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 10692 6860 10744 6866
rect 10428 6798 10456 6854
rect 10692 6802 10744 6808
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 5370 10548 6734
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10704 5166 10732 6802
rect 11072 6730 11100 7278
rect 11256 6798 11284 7278
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10888 4826 10916 5170
rect 11256 5030 11284 6734
rect 11716 5166 11744 6734
rect 11808 5234 11836 9522
rect 12084 8566 12112 15370
rect 12176 15026 12204 17326
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12268 16794 12296 17206
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12452 16658 12480 18090
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12268 11370 12296 16186
rect 12452 14346 12480 16594
rect 12636 15502 12664 16934
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 14074 12480 14282
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12728 12434 12756 19790
rect 12912 17610 12940 20266
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 13004 17542 13032 18226
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 14074 12848 14350
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 13004 12918 13032 17478
rect 13188 17270 13216 23598
rect 13280 22658 13308 23666
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 13611 23420 13919 23429
rect 13611 23418 13617 23420
rect 13673 23418 13697 23420
rect 13753 23418 13777 23420
rect 13833 23418 13857 23420
rect 13913 23418 13919 23420
rect 13673 23366 13675 23418
rect 13855 23366 13857 23418
rect 13611 23364 13617 23366
rect 13673 23364 13697 23366
rect 13753 23364 13777 23366
rect 13833 23364 13857 23366
rect 13913 23364 13919 23366
rect 13611 23355 13919 23364
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 13280 22642 13492 22658
rect 13280 22636 13504 22642
rect 13280 22630 13452 22636
rect 13372 22166 13400 22630
rect 13452 22578 13504 22584
rect 13611 22332 13919 22341
rect 13611 22330 13617 22332
rect 13673 22330 13697 22332
rect 13753 22330 13777 22332
rect 13833 22330 13857 22332
rect 13913 22330 13919 22332
rect 13673 22278 13675 22330
rect 13855 22278 13857 22330
rect 13611 22276 13617 22278
rect 13673 22276 13697 22278
rect 13753 22276 13777 22278
rect 13833 22276 13857 22278
rect 13913 22276 13919 22278
rect 13611 22267 13919 22276
rect 13360 22160 13412 22166
rect 13360 22102 13412 22108
rect 13372 20398 13400 22102
rect 14016 21554 14044 23054
rect 14200 22574 14228 23530
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13611 21244 13919 21253
rect 13611 21242 13617 21244
rect 13673 21242 13697 21244
rect 13753 21242 13777 21244
rect 13833 21242 13857 21244
rect 13913 21242 13919 21244
rect 13673 21190 13675 21242
rect 13855 21190 13857 21242
rect 13611 21188 13617 21190
rect 13673 21188 13697 21190
rect 13753 21188 13777 21190
rect 13833 21188 13857 21190
rect 13913 21188 13919 21190
rect 13611 21179 13919 21188
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 13372 19854 13400 20334
rect 13464 19854 13492 20878
rect 14200 20602 14228 22510
rect 14476 20942 14504 25706
rect 14568 24206 14596 27950
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14752 23662 14780 25978
rect 15028 24698 15056 28086
rect 15488 28082 15516 28494
rect 15580 28150 15608 29106
rect 15764 28490 15792 29106
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15568 28144 15620 28150
rect 15568 28086 15620 28092
rect 15476 28076 15528 28082
rect 15476 28018 15528 28024
rect 15488 25226 15516 28018
rect 15764 26994 15792 28426
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 15948 25294 15976 28358
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16040 27606 16068 28086
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 16040 27470 16068 27542
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24818 15240 25094
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15028 24670 15148 24698
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14752 23050 14780 23598
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22642 14688 22918
rect 14752 22710 14780 22986
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14200 20398 14228 20538
rect 14384 20534 14412 20742
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 13611 20156 13919 20165
rect 13611 20154 13617 20156
rect 13673 20154 13697 20156
rect 13753 20154 13777 20156
rect 13833 20154 13857 20156
rect 13913 20154 13919 20156
rect 13673 20102 13675 20154
rect 13855 20102 13857 20154
rect 13611 20100 13617 20102
rect 13673 20100 13697 20102
rect 13753 20100 13777 20102
rect 13833 20100 13857 20102
rect 13913 20100 13919 20102
rect 13611 20091 13919 20100
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13372 16250 13400 19314
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13464 15570 13492 19790
rect 13611 19068 13919 19077
rect 13611 19066 13617 19068
rect 13673 19066 13697 19068
rect 13753 19066 13777 19068
rect 13833 19066 13857 19068
rect 13913 19066 13919 19068
rect 13673 19014 13675 19066
rect 13855 19014 13857 19066
rect 13611 19012 13617 19014
rect 13673 19012 13697 19014
rect 13753 19012 13777 19014
rect 13833 19012 13857 19014
rect 13913 19012 13919 19014
rect 13611 19003 13919 19012
rect 13611 17980 13919 17989
rect 13611 17978 13617 17980
rect 13673 17978 13697 17980
rect 13753 17978 13777 17980
rect 13833 17978 13857 17980
rect 13913 17978 13919 17980
rect 13673 17926 13675 17978
rect 13855 17926 13857 17978
rect 13611 17924 13617 17926
rect 13673 17924 13697 17926
rect 13753 17924 13777 17926
rect 13833 17924 13857 17926
rect 13913 17924 13919 17926
rect 13611 17915 13919 17924
rect 14384 17338 14412 19790
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 13611 16892 13919 16901
rect 13611 16890 13617 16892
rect 13673 16890 13697 16892
rect 13753 16890 13777 16892
rect 13833 16890 13857 16892
rect 13913 16890 13919 16892
rect 13673 16838 13675 16890
rect 13855 16838 13857 16890
rect 13611 16836 13617 16838
rect 13673 16836 13697 16838
rect 13753 16836 13777 16838
rect 13833 16836 13857 16838
rect 13913 16836 13919 16838
rect 13611 16827 13919 16836
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 14292 16182 14320 16458
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 13611 15804 13919 15813
rect 13611 15802 13617 15804
rect 13673 15802 13697 15804
rect 13753 15802 13777 15804
rect 13833 15802 13857 15804
rect 13913 15802 13919 15804
rect 13673 15750 13675 15802
rect 13855 15750 13857 15802
rect 13611 15748 13617 15750
rect 13673 15748 13697 15750
rect 13753 15748 13777 15750
rect 13833 15748 13857 15750
rect 13913 15748 13919 15750
rect 13611 15739 13919 15748
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 14292 15502 14320 16118
rect 14476 15910 14504 16390
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14568 15638 14596 19790
rect 14660 18970 14688 20334
rect 14752 19990 14780 20334
rect 14844 19990 14872 24142
rect 15028 23866 15056 24550
rect 15120 24342 15148 24670
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15028 23118 15056 23802
rect 15304 23662 15332 24890
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 23866 15424 24754
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15488 24070 15516 24618
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15212 23186 15240 23598
rect 15396 23254 15424 23802
rect 15488 23730 15516 24006
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15384 23248 15436 23254
rect 15384 23190 15436 23196
rect 15488 23186 15516 23462
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 15580 22642 15608 24074
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15488 22522 15516 22578
rect 15672 22522 15700 25230
rect 16120 25152 16172 25158
rect 16120 25094 16172 25100
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15856 23730 15884 24142
rect 16132 23866 16160 25094
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15488 22494 15700 22522
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16040 20466 16068 21490
rect 16224 20534 16252 32778
rect 16776 32366 16804 32778
rect 17831 32668 18139 32677
rect 17831 32666 17837 32668
rect 17893 32666 17917 32668
rect 17973 32666 17997 32668
rect 18053 32666 18077 32668
rect 18133 32666 18139 32668
rect 17893 32614 17895 32666
rect 18075 32614 18077 32666
rect 17831 32612 17837 32614
rect 17893 32612 17917 32614
rect 17973 32612 17997 32614
rect 18053 32612 18077 32614
rect 18133 32612 18139 32614
rect 17831 32603 18139 32612
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16316 30666 16344 31282
rect 16304 30660 16356 30666
rect 16304 30602 16356 30608
rect 16304 27396 16356 27402
rect 16304 27338 16356 27344
rect 16316 25838 16344 27338
rect 16396 26988 16448 26994
rect 16396 26930 16448 26936
rect 16304 25832 16356 25838
rect 16304 25774 16356 25780
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 16316 24818 16344 25366
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16408 24206 16436 26930
rect 16672 26920 16724 26926
rect 16672 26862 16724 26868
rect 16684 26586 16712 26862
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 25974 16712 26522
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16488 25832 16540 25838
rect 16488 25774 16540 25780
rect 16500 24410 16528 25774
rect 16684 25498 16712 25910
rect 16672 25492 16724 25498
rect 16672 25434 16724 25440
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16408 22234 16436 22578
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15672 20058 15700 20402
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 14832 19984 14884 19990
rect 14832 19926 14884 19932
rect 15856 19854 15884 20198
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15660 19780 15712 19786
rect 15660 19722 15712 19728
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14752 18766 14780 19246
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 14752 18358 14780 18702
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 15212 17678 15240 18566
rect 15396 17882 15424 18702
rect 15672 18290 15700 19722
rect 16040 19446 16068 20402
rect 16028 19440 16080 19446
rect 16028 19382 16080 19388
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15764 18426 15792 18634
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 16040 18358 16068 19382
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15396 17202 15424 17818
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15948 16794 15976 17070
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14752 16046 14780 16594
rect 15212 16182 15240 16662
rect 15384 16584 15436 16590
rect 15488 16572 15516 16730
rect 15436 16544 15516 16572
rect 15384 16526 15436 16532
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 14006 13124 14282
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12728 12406 12848 12434
rect 12268 11354 12572 11370
rect 12256 11348 12572 11354
rect 12308 11342 12572 11348
rect 12256 11290 12308 11296
rect 12268 11259 12296 11290
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12176 10674 12204 11154
rect 12544 11150 12572 11342
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12452 10674 12480 11018
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12544 9178 12572 10678
rect 12636 10266 12664 11018
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 9450 12756 10950
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6458 12572 7142
rect 12820 6730 12848 12406
rect 13096 11150 13124 13330
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12912 10742 12940 11086
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13096 7002 13124 7278
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5302 12480 6190
rect 13188 5370 13216 12650
rect 13280 11762 13308 13806
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13280 10742 13308 11698
rect 13464 11082 13492 14962
rect 13611 14716 13919 14725
rect 13611 14714 13617 14716
rect 13673 14714 13697 14716
rect 13753 14714 13777 14716
rect 13833 14714 13857 14716
rect 13913 14714 13919 14716
rect 13673 14662 13675 14714
rect 13855 14662 13857 14714
rect 13611 14660 13617 14662
rect 13673 14660 13697 14662
rect 13753 14660 13777 14662
rect 13833 14660 13857 14662
rect 13913 14660 13919 14662
rect 13611 14651 13919 14660
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13938 13768 14350
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13611 13628 13919 13637
rect 13611 13626 13617 13628
rect 13673 13626 13697 13628
rect 13753 13626 13777 13628
rect 13833 13626 13857 13628
rect 13913 13626 13919 13628
rect 13673 13574 13675 13626
rect 13855 13574 13857 13626
rect 13611 13572 13617 13574
rect 13673 13572 13697 13574
rect 13753 13572 13777 13574
rect 13833 13572 13857 13574
rect 13913 13572 13919 13574
rect 13611 13563 13919 13572
rect 14108 13258 14136 13806
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14752 12918 14780 15982
rect 16408 15570 16436 22170
rect 16500 21554 16528 24346
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16684 18970 16712 20266
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16684 18426 16712 18906
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 16590 16620 17478
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 15672 15026 15700 15438
rect 16224 15026 16252 15438
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15108 13320 15160 13326
rect 15212 13274 15240 13806
rect 15396 13530 15424 13874
rect 15672 13530 15700 14962
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15752 13320 15804 13326
rect 15160 13268 15332 13274
rect 15108 13262 15332 13268
rect 15752 13262 15804 13268
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 15120 13246 15332 13262
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 13611 12540 13919 12549
rect 13611 12538 13617 12540
rect 13673 12538 13697 12540
rect 13753 12538 13777 12540
rect 13833 12538 13857 12540
rect 13913 12538 13919 12540
rect 13673 12486 13675 12538
rect 13855 12486 13857 12538
rect 13611 12484 13617 12486
rect 13673 12484 13697 12486
rect 13753 12484 13777 12486
rect 13833 12484 13857 12486
rect 13913 12484 13919 12486
rect 13611 12475 13919 12484
rect 14568 12238 14596 12582
rect 15212 12238 15240 12786
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 14568 11762 14596 12174
rect 15212 11830 15240 12174
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15304 11762 15332 13246
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15580 12850 15608 13194
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15764 12238 15792 13262
rect 16408 12850 16436 13262
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16592 12782 16620 15574
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 15764 11830 15792 12174
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 16500 11762 16528 12174
rect 16592 11762 16620 12718
rect 16776 12434 16804 32302
rect 16856 31952 16908 31958
rect 16856 31894 16908 31900
rect 16868 30734 16896 31894
rect 17132 31884 17184 31890
rect 17132 31826 17184 31832
rect 17144 31346 17172 31826
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 17328 31482 17356 31758
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17040 31136 17092 31142
rect 17040 31078 17092 31084
rect 17052 30734 17080 31078
rect 17420 30938 17448 32302
rect 17880 31822 17908 32370
rect 18248 32026 18276 32370
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 17868 31816 17920 31822
rect 17696 31776 17868 31804
rect 17696 31346 17724 31776
rect 17868 31758 17920 31764
rect 17831 31580 18139 31589
rect 17831 31578 17837 31580
rect 17893 31578 17917 31580
rect 17973 31578 17997 31580
rect 18053 31578 18077 31580
rect 18133 31578 18139 31580
rect 17893 31526 17895 31578
rect 18075 31526 18077 31578
rect 17831 31524 17837 31526
rect 17893 31524 17917 31526
rect 17973 31524 17997 31526
rect 18053 31524 18077 31526
rect 18133 31524 18139 31526
rect 17831 31515 18139 31524
rect 19352 31414 19380 32846
rect 19536 32502 19564 33322
rect 20272 33046 20300 33322
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20260 33040 20312 33046
rect 20260 32982 20312 32988
rect 20456 32978 20484 33254
rect 22052 33212 22360 33221
rect 22052 33210 22058 33212
rect 22114 33210 22138 33212
rect 22194 33210 22218 33212
rect 22274 33210 22298 33212
rect 22354 33210 22360 33212
rect 22114 33158 22116 33210
rect 22296 33158 22298 33210
rect 22052 33156 22058 33158
rect 22114 33156 22138 33158
rect 22194 33156 22218 33158
rect 22274 33156 22298 33158
rect 22354 33156 22360 33158
rect 22052 33147 22360 33156
rect 20444 32972 20496 32978
rect 20444 32914 20496 32920
rect 20628 32972 20680 32978
rect 20628 32914 20680 32920
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 19524 32496 19576 32502
rect 19524 32438 19576 32444
rect 20640 32026 20668 32914
rect 22836 32904 22888 32910
rect 22836 32846 22888 32852
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21284 32366 21312 32710
rect 22020 32434 22048 32710
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 21272 32360 21324 32366
rect 21272 32302 21324 32308
rect 21088 32292 21140 32298
rect 21088 32234 21140 32240
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 19340 31408 19392 31414
rect 19340 31350 19392 31356
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 17831 30492 18139 30501
rect 17831 30490 17837 30492
rect 17893 30490 17917 30492
rect 17973 30490 17997 30492
rect 18053 30490 18077 30492
rect 18133 30490 18139 30492
rect 17893 30438 17895 30490
rect 18075 30438 18077 30490
rect 17831 30436 17837 30438
rect 17893 30436 17917 30438
rect 17973 30436 17997 30438
rect 18053 30436 18077 30438
rect 18133 30436 18139 30438
rect 17831 30427 18139 30436
rect 18800 30326 18828 30602
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 17831 29404 18139 29413
rect 17831 29402 17837 29404
rect 17893 29402 17917 29404
rect 17973 29402 17997 29404
rect 18053 29402 18077 29404
rect 18133 29402 18139 29404
rect 17893 29350 17895 29402
rect 18075 29350 18077 29402
rect 17831 29348 17837 29350
rect 17893 29348 17917 29350
rect 17973 29348 17997 29350
rect 18053 29348 18077 29350
rect 18133 29348 18139 29350
rect 17831 29339 18139 29348
rect 19260 28490 19288 29582
rect 19524 29504 19576 29510
rect 19524 29446 19576 29452
rect 19536 29170 19564 29446
rect 20180 29306 20208 30194
rect 20364 29646 20392 31282
rect 20548 31278 20576 31894
rect 21100 31890 21128 32234
rect 22052 32124 22360 32133
rect 22052 32122 22058 32124
rect 22114 32122 22138 32124
rect 22194 32122 22218 32124
rect 22274 32122 22298 32124
rect 22354 32122 22360 32124
rect 22114 32070 22116 32122
rect 22296 32070 22298 32122
rect 22052 32068 22058 32070
rect 22114 32068 22138 32070
rect 22194 32068 22218 32070
rect 22274 32068 22298 32070
rect 22354 32068 22360 32070
rect 22052 32059 22360 32068
rect 22480 31958 22508 32370
rect 22848 32230 22876 32846
rect 24596 32434 24624 32914
rect 25424 32842 25452 33322
rect 30493 33212 30801 33221
rect 30493 33210 30499 33212
rect 30555 33210 30579 33212
rect 30635 33210 30659 33212
rect 30715 33210 30739 33212
rect 30795 33210 30801 33212
rect 30555 33158 30557 33210
rect 30737 33158 30739 33210
rect 30493 33156 30499 33158
rect 30555 33156 30579 33158
rect 30635 33156 30659 33158
rect 30715 33156 30739 33158
rect 30795 33156 30801 33158
rect 30493 33147 30801 33156
rect 25412 32836 25464 32842
rect 25412 32778 25464 32784
rect 26272 32668 26580 32677
rect 26272 32666 26278 32668
rect 26334 32666 26358 32668
rect 26414 32666 26438 32668
rect 26494 32666 26518 32668
rect 26574 32666 26580 32668
rect 26334 32614 26336 32666
rect 26516 32614 26518 32666
rect 26272 32612 26278 32614
rect 26334 32612 26358 32614
rect 26414 32612 26438 32614
rect 26494 32612 26518 32614
rect 26574 32612 26580 32614
rect 26272 32603 26580 32612
rect 31312 32434 31340 33322
rect 33336 32434 33364 33322
rect 34713 32668 35021 32677
rect 34713 32666 34719 32668
rect 34775 32666 34799 32668
rect 34855 32666 34879 32668
rect 34935 32666 34959 32668
rect 35015 32666 35021 32668
rect 34775 32614 34777 32666
rect 34957 32614 34959 32666
rect 34713 32612 34719 32614
rect 34775 32612 34799 32614
rect 34855 32612 34879 32614
rect 34935 32612 34959 32614
rect 35015 32612 35021 32614
rect 34713 32603 35021 32612
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 28080 32428 28132 32434
rect 28080 32370 28132 32376
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22468 31952 22520 31958
rect 22468 31894 22520 31900
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20824 31482 20852 31758
rect 21100 31754 21128 31826
rect 22848 31822 22876 32166
rect 23216 32026 23244 32370
rect 23388 32360 23440 32366
rect 23388 32302 23440 32308
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 21180 31816 21232 31822
rect 21180 31758 21232 31764
rect 21364 31816 21416 31822
rect 22836 31816 22888 31822
rect 21364 31758 21416 31764
rect 22664 31776 22836 31804
rect 21088 31748 21140 31754
rect 21088 31690 21140 31696
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20548 29714 20576 31214
rect 21008 30938 21036 31282
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20536 29708 20588 29714
rect 20536 29650 20588 29656
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19524 29164 19576 29170
rect 20364 29152 20392 29582
rect 20548 29238 20576 29650
rect 20536 29232 20588 29238
rect 20536 29174 20588 29180
rect 20640 29170 20668 29990
rect 20824 29714 20852 30194
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20732 29170 20760 29582
rect 20444 29164 20496 29170
rect 20364 29124 20444 29152
rect 19524 29106 19576 29112
rect 20444 29106 20496 29112
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 17831 28316 18139 28325
rect 17831 28314 17837 28316
rect 17893 28314 17917 28316
rect 17973 28314 17997 28316
rect 18053 28314 18077 28316
rect 18133 28314 18139 28316
rect 17893 28262 17895 28314
rect 18075 28262 18077 28314
rect 17831 28260 17837 28262
rect 17893 28260 17917 28262
rect 17973 28260 17997 28262
rect 18053 28260 18077 28262
rect 18133 28260 18139 28262
rect 17831 28251 18139 28260
rect 19260 28082 19288 28426
rect 19352 28150 19380 29106
rect 20732 28966 20760 29106
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20732 28694 20760 28902
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20732 28558 20760 28630
rect 20824 28626 20852 29650
rect 20916 29578 20944 30194
rect 20904 29572 20956 29578
rect 20904 29514 20956 29520
rect 20812 28620 20864 28626
rect 20812 28562 20864 28568
rect 20916 28558 20944 29514
rect 21192 28762 21220 31758
rect 21376 31278 21404 31758
rect 22664 31346 22692 31776
rect 22836 31758 22888 31764
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 22756 31346 22784 31622
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22744 31340 22796 31346
rect 22744 31282 22796 31288
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 21364 31272 21416 31278
rect 21364 31214 21416 31220
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21376 29306 21404 31214
rect 21468 30734 21496 31214
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21468 29510 21496 30670
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21456 29504 21508 29510
rect 21456 29446 21508 29452
rect 21364 29300 21416 29306
rect 21364 29242 21416 29248
rect 21652 29238 21680 29514
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 19812 28218 19840 28494
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 17831 27228 18139 27237
rect 17831 27226 17837 27228
rect 17893 27226 17917 27228
rect 17973 27226 17997 27228
rect 18053 27226 18077 27228
rect 18133 27226 18139 27228
rect 17893 27174 17895 27226
rect 18075 27174 18077 27226
rect 17831 27172 17837 27174
rect 17893 27172 17917 27174
rect 17973 27172 17997 27174
rect 18053 27172 18077 27174
rect 18133 27172 18139 27174
rect 17831 27163 18139 27172
rect 18248 27130 18276 27406
rect 18236 27124 18288 27130
rect 18236 27066 18288 27072
rect 18248 26450 18276 27066
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 16868 26042 16896 26250
rect 17831 26140 18139 26149
rect 17831 26138 17837 26140
rect 17893 26138 17917 26140
rect 17973 26138 17997 26140
rect 18053 26138 18077 26140
rect 18133 26138 18139 26140
rect 17893 26086 17895 26138
rect 18075 26086 18077 26138
rect 17831 26084 17837 26086
rect 17893 26084 17917 26086
rect 17973 26084 17997 26086
rect 18053 26084 18077 26086
rect 18133 26084 18139 26086
rect 17831 26075 18139 26084
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17052 24954 17080 25842
rect 17831 25052 18139 25061
rect 17831 25050 17837 25052
rect 17893 25050 17917 25052
rect 17973 25050 17997 25052
rect 18053 25050 18077 25052
rect 18133 25050 18139 25052
rect 17893 24998 17895 25050
rect 18075 24998 18077 25050
rect 17831 24996 17837 24998
rect 17893 24996 17917 24998
rect 17973 24996 17997 24998
rect 18053 24996 18077 24998
rect 18133 24996 18139 24998
rect 17831 24987 18139 24996
rect 17040 24948 17092 24954
rect 17040 24890 17092 24896
rect 18248 24818 18276 26250
rect 18340 25702 18368 26930
rect 18972 26512 19024 26518
rect 18972 26454 19024 26460
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17144 23730 17172 24006
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17144 22642 17172 23666
rect 17328 23186 17356 24686
rect 18052 24608 18104 24614
rect 18052 24550 18104 24556
rect 17960 24200 18012 24206
rect 18064 24188 18092 24550
rect 18012 24160 18092 24188
rect 17960 24142 18012 24148
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17132 22636 17184 22642
rect 17132 22578 17184 22584
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16868 17270 16896 21286
rect 17328 21146 17356 23122
rect 17604 23118 17632 24006
rect 17831 23964 18139 23973
rect 17831 23962 17837 23964
rect 17893 23962 17917 23964
rect 17973 23962 17997 23964
rect 18053 23962 18077 23964
rect 18133 23962 18139 23964
rect 17893 23910 17895 23962
rect 18075 23910 18077 23962
rect 17831 23908 17837 23910
rect 17893 23908 17917 23910
rect 17973 23908 17997 23910
rect 18053 23908 18077 23910
rect 18133 23908 18139 23910
rect 17831 23899 18139 23908
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17831 22876 18139 22885
rect 17831 22874 17837 22876
rect 17893 22874 17917 22876
rect 17973 22874 17997 22876
rect 18053 22874 18077 22876
rect 18133 22874 18139 22876
rect 17893 22822 17895 22874
rect 18075 22822 18077 22874
rect 17831 22820 17837 22822
rect 17893 22820 17917 22822
rect 17973 22820 17997 22822
rect 18053 22820 18077 22822
rect 18133 22820 18139 22822
rect 17831 22811 18139 22820
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 22166 18000 22374
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 18064 22030 18092 22442
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17831 21788 18139 21797
rect 17831 21786 17837 21788
rect 17893 21786 17917 21788
rect 17973 21786 17997 21788
rect 18053 21786 18077 21788
rect 18133 21786 18139 21788
rect 17893 21734 17895 21786
rect 18075 21734 18077 21786
rect 17831 21732 17837 21734
rect 17893 21732 17917 21734
rect 17973 21732 17997 21734
rect 18053 21732 18077 21734
rect 18133 21732 18139 21734
rect 17831 21723 18139 21732
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 18340 20942 18368 25638
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18432 22030 18460 23598
rect 18708 23322 18736 24074
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18708 22642 18736 23258
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 17831 20700 18139 20709
rect 17831 20698 17837 20700
rect 17893 20698 17917 20700
rect 17973 20698 17997 20700
rect 18053 20698 18077 20700
rect 18133 20698 18139 20700
rect 17893 20646 17895 20698
rect 18075 20646 18077 20698
rect 17831 20644 17837 20646
rect 17893 20644 17917 20646
rect 17973 20644 17997 20646
rect 18053 20644 18077 20646
rect 18133 20644 18139 20646
rect 17831 20635 18139 20644
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 17144 19378 17172 19722
rect 17831 19612 18139 19621
rect 17831 19610 17837 19612
rect 17893 19610 17917 19612
rect 17973 19610 17997 19612
rect 18053 19610 18077 19612
rect 18133 19610 18139 19612
rect 17893 19558 17895 19610
rect 18075 19558 18077 19610
rect 17831 19556 17837 19558
rect 17893 19556 17917 19558
rect 17973 19556 17997 19558
rect 18053 19556 18077 19558
rect 18133 19556 18139 19558
rect 17831 19547 18139 19556
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 13938 16896 14826
rect 16960 14074 16988 18566
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16868 13258 16896 13874
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 17144 12434 17172 19314
rect 17831 18524 18139 18533
rect 17831 18522 17837 18524
rect 17893 18522 17917 18524
rect 17973 18522 17997 18524
rect 18053 18522 18077 18524
rect 18133 18522 18139 18524
rect 17893 18470 17895 18522
rect 18075 18470 18077 18522
rect 17831 18468 17837 18470
rect 17893 18468 17917 18470
rect 17973 18468 17997 18470
rect 18053 18468 18077 18470
rect 18133 18468 18139 18470
rect 17831 18459 18139 18468
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17236 16590 17264 17138
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17328 16522 17356 17546
rect 17512 17134 17540 17614
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 16658 17540 17070
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17328 16232 17356 16458
rect 16776 12406 16896 12434
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 13611 11452 13919 11461
rect 13611 11450 13617 11452
rect 13673 11450 13697 11452
rect 13753 11450 13777 11452
rect 13833 11450 13857 11452
rect 13913 11450 13919 11452
rect 13673 11398 13675 11450
rect 13855 11398 13857 11450
rect 13611 11396 13617 11398
rect 13673 11396 13697 11398
rect 13753 11396 13777 11398
rect 13833 11396 13857 11398
rect 13913 11396 13919 11398
rect 13611 11387 13919 11396
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 13611 10364 13919 10373
rect 13611 10362 13617 10364
rect 13673 10362 13697 10364
rect 13753 10362 13777 10364
rect 13833 10362 13857 10364
rect 13913 10362 13919 10364
rect 13673 10310 13675 10362
rect 13855 10310 13857 10362
rect 13611 10308 13617 10310
rect 13673 10308 13697 10310
rect 13753 10308 13777 10310
rect 13833 10308 13857 10310
rect 13913 10308 13919 10310
rect 13611 10299 13919 10308
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10520 4146 10548 4558
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10612 3534 10640 4082
rect 10888 3602 10916 4082
rect 11256 4078 11284 4966
rect 11808 4554 11836 5170
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4826 12020 4966
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12452 4622 12480 5238
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 13372 4214 13400 9862
rect 13611 9276 13919 9285
rect 13611 9274 13617 9276
rect 13673 9274 13697 9276
rect 13753 9274 13777 9276
rect 13833 9274 13857 9276
rect 13913 9274 13919 9276
rect 13673 9222 13675 9274
rect 13855 9222 13857 9274
rect 13611 9220 13617 9222
rect 13673 9220 13697 9222
rect 13753 9220 13777 9222
rect 13833 9220 13857 9222
rect 13913 9220 13919 9222
rect 13611 9211 13919 9220
rect 13611 8188 13919 8197
rect 13611 8186 13617 8188
rect 13673 8186 13697 8188
rect 13753 8186 13777 8188
rect 13833 8186 13857 8188
rect 13913 8186 13919 8188
rect 13673 8134 13675 8186
rect 13855 8134 13857 8186
rect 13611 8132 13617 8134
rect 13673 8132 13697 8134
rect 13753 8132 13777 8134
rect 13833 8132 13857 8134
rect 13913 8132 13919 8134
rect 13611 8123 13919 8132
rect 13611 7100 13919 7109
rect 13611 7098 13617 7100
rect 13673 7098 13697 7100
rect 13753 7098 13777 7100
rect 13833 7098 13857 7100
rect 13913 7098 13919 7100
rect 13673 7046 13675 7098
rect 13855 7046 13857 7098
rect 13611 7044 13617 7046
rect 13673 7044 13697 7046
rect 13753 7044 13777 7046
rect 13833 7044 13857 7046
rect 13913 7044 13919 7046
rect 13611 7035 13919 7044
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6390 13676 6598
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13611 6012 13919 6021
rect 13611 6010 13617 6012
rect 13673 6010 13697 6012
rect 13753 6010 13777 6012
rect 13833 6010 13857 6012
rect 13913 6010 13919 6012
rect 13673 5958 13675 6010
rect 13855 5958 13857 6010
rect 13611 5956 13617 5958
rect 13673 5956 13697 5958
rect 13753 5956 13777 5958
rect 13833 5956 13857 5958
rect 13913 5956 13919 5958
rect 13611 5947 13919 5956
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13611 4924 13919 4933
rect 13611 4922 13617 4924
rect 13673 4922 13697 4924
rect 13753 4922 13777 4924
rect 13833 4922 13857 4924
rect 13913 4922 13919 4924
rect 13673 4870 13675 4922
rect 13855 4870 13857 4922
rect 13611 4868 13617 4870
rect 13673 4868 13697 4870
rect 13753 4868 13777 4870
rect 13833 4868 13857 4870
rect 13913 4868 13919 4870
rect 13611 4859 13919 4868
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10888 3058 10916 3538
rect 13004 3534 13032 3878
rect 13611 3836 13919 3845
rect 13611 3834 13617 3836
rect 13673 3834 13697 3836
rect 13753 3834 13777 3836
rect 13833 3834 13857 3836
rect 13913 3834 13919 3836
rect 13673 3782 13675 3834
rect 13855 3782 13857 3834
rect 13611 3780 13617 3782
rect 13673 3780 13697 3782
rect 13753 3780 13777 3782
rect 13833 3780 13857 3782
rect 13913 3780 13919 3782
rect 13611 3771 13919 3780
rect 14016 3738 14044 4082
rect 14200 4078 14228 4626
rect 14292 4622 14320 4966
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12360 3194 12388 3470
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 13611 2748 13919 2757
rect 13611 2746 13617 2748
rect 13673 2746 13697 2748
rect 13753 2746 13777 2748
rect 13833 2746 13857 2748
rect 13913 2746 13919 2748
rect 13673 2694 13675 2746
rect 13855 2694 13857 2746
rect 13611 2692 13617 2694
rect 13673 2692 13697 2694
rect 13753 2692 13777 2694
rect 13833 2692 13857 2694
rect 13913 2692 13919 2694
rect 13611 2683 13919 2692
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 14016 2446 14044 3674
rect 14200 2990 14228 4014
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 2990 14320 3334
rect 14384 3194 14412 10406
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15120 7206 15148 8910
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6866 15148 7142
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15212 5234 15240 7414
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 6798 15700 7142
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4146 14964 4966
rect 15856 4622 15884 11222
rect 16776 11150 16804 11766
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8498 16344 8910
rect 16592 8906 16620 9862
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16684 8294 16712 11018
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15948 7546 15976 7754
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 16684 7478 16712 8230
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4214 15608 4422
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14752 3194 14780 3402
rect 15672 3194 15700 3470
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14384 2514 14412 3130
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 15488 2446 15516 2926
rect 15856 2774 15884 4558
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 3942 16344 4422
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 15856 2746 15976 2774
rect 15948 2650 15976 2746
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16316 2446 16344 3878
rect 16684 3602 16712 3878
rect 16868 3738 16896 12406
rect 17052 12406 17172 12434
rect 17236 16204 17356 16232
rect 17236 12434 17264 16204
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17420 15638 17448 16050
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17328 14482 17356 15370
rect 17512 15178 17540 16594
rect 17604 16454 17632 17478
rect 17831 17436 18139 17445
rect 17831 17434 17837 17436
rect 17893 17434 17917 17436
rect 17973 17434 17997 17436
rect 18053 17434 18077 17436
rect 18133 17434 18139 17436
rect 17893 17382 17895 17434
rect 18075 17382 18077 17434
rect 17831 17380 17837 17382
rect 17893 17380 17917 17382
rect 17973 17380 17997 17382
rect 18053 17380 18077 17382
rect 18133 17380 18139 17382
rect 17831 17371 18139 17380
rect 18248 17270 18276 18022
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17420 15150 17540 15178
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17420 12481 17448 15150
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17406 12472 17462 12481
rect 17236 12406 17356 12434
rect 17406 12407 17462 12416
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16960 11150 16988 12106
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 17052 8498 17080 12406
rect 17328 10062 17356 12406
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17052 7342 17080 8434
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16960 3194 16988 3402
rect 17144 3194 17172 9658
rect 17236 9178 17264 9930
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17328 8922 17356 9998
rect 17420 9586 17448 12407
rect 17512 12238 17540 13194
rect 17604 12986 17632 16390
rect 17831 16348 18139 16357
rect 17831 16346 17837 16348
rect 17893 16346 17917 16348
rect 17973 16346 17997 16348
rect 18053 16346 18077 16348
rect 18133 16346 18139 16348
rect 17893 16294 17895 16346
rect 18075 16294 18077 16346
rect 17831 16292 17837 16294
rect 17893 16292 17917 16294
rect 17973 16292 17997 16294
rect 18053 16292 18077 16294
rect 18133 16292 18139 16294
rect 17831 16283 18139 16292
rect 18248 16182 18276 17206
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17696 15434 17724 16050
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17696 14414 17724 15370
rect 17831 15260 18139 15269
rect 17831 15258 17837 15260
rect 17893 15258 17917 15260
rect 17973 15258 17997 15260
rect 18053 15258 18077 15260
rect 18133 15258 18139 15260
rect 17893 15206 17895 15258
rect 18075 15206 18077 15258
rect 17831 15204 17837 15206
rect 17893 15204 17917 15206
rect 17973 15204 17997 15206
rect 18053 15204 18077 15206
rect 18133 15204 18139 15206
rect 17831 15195 18139 15204
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18156 14414 18184 14894
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 17696 13938 17724 14350
rect 17831 14172 18139 14181
rect 17831 14170 17837 14172
rect 17893 14170 17917 14172
rect 17973 14170 17997 14172
rect 18053 14170 18077 14172
rect 18133 14170 18139 14172
rect 17893 14118 17895 14170
rect 18075 14118 18077 14170
rect 17831 14116 17837 14118
rect 17893 14116 17917 14118
rect 17973 14116 17997 14118
rect 18053 14116 18077 14118
rect 18133 14116 18139 14118
rect 17831 14107 18139 14116
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 18248 13190 18276 14962
rect 18340 13462 18368 15438
rect 18432 15162 18460 21966
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18524 18358 18552 18566
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18328 13456 18380 13462
rect 18328 13398 18380 13404
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 17831 13084 18139 13093
rect 17831 13082 17837 13084
rect 17893 13082 17917 13084
rect 17973 13082 17997 13084
rect 18053 13082 18077 13084
rect 18133 13082 18139 13084
rect 17893 13030 17895 13082
rect 18075 13030 18077 13082
rect 17831 13028 17837 13030
rect 17893 13028 17917 13030
rect 17973 13028 17997 13030
rect 18053 13028 18077 13030
rect 18133 13028 18139 13030
rect 17831 13019 18139 13028
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12306 18092 12786
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 11150 17540 12174
rect 17831 11996 18139 12005
rect 17831 11994 17837 11996
rect 17893 11994 17917 11996
rect 17973 11994 17997 11996
rect 18053 11994 18077 11996
rect 18133 11994 18139 11996
rect 17893 11942 17895 11994
rect 18075 11942 18077 11994
rect 17831 11940 17837 11942
rect 17893 11940 17917 11942
rect 17973 11940 17997 11942
rect 18053 11940 18077 11942
rect 18133 11940 18139 11942
rect 17831 11931 18139 11940
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17831 10908 18139 10917
rect 17831 10906 17837 10908
rect 17893 10906 17917 10908
rect 17973 10906 17997 10908
rect 18053 10906 18077 10908
rect 18133 10906 18139 10908
rect 17893 10854 17895 10906
rect 18075 10854 18077 10906
rect 17831 10852 17837 10854
rect 17893 10852 17917 10854
rect 17973 10852 17997 10854
rect 18053 10852 18077 10854
rect 18133 10852 18139 10854
rect 17831 10843 18139 10852
rect 18248 10742 18276 13126
rect 18340 12918 18368 13262
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18432 12850 18460 14350
rect 18800 13938 18828 20470
rect 18984 20466 19012 26454
rect 19352 26450 19380 28086
rect 19996 28014 20024 28494
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19892 27532 19944 27538
rect 19892 27474 19944 27480
rect 19524 27396 19576 27402
rect 19524 27338 19576 27344
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19352 24750 19380 26386
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19352 22574 19380 23802
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19444 22030 19472 23054
rect 19536 22094 19564 27338
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19812 27062 19840 27270
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19628 23254 19656 25842
rect 19812 25498 19840 26998
rect 19904 26246 19932 27474
rect 20548 26790 20576 28358
rect 20916 28150 20944 28494
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 21008 26994 21036 27338
rect 21192 26994 21220 27406
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20904 26784 20956 26790
rect 20904 26726 20956 26732
rect 19892 26240 19944 26246
rect 19892 26182 19944 26188
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19720 23594 19748 24074
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19616 23248 19668 23254
rect 19616 23190 19668 23196
rect 19720 23118 19748 23530
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19536 22066 19748 22094
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19352 20618 19380 21898
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19076 20602 19380 20618
rect 19064 20596 19380 20602
rect 19116 20590 19380 20596
rect 19064 20538 19116 20544
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19156 20460 19208 20466
rect 19340 20460 19392 20466
rect 19156 20402 19208 20408
rect 19260 20420 19340 20448
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19076 19378 19104 20198
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19168 19174 19196 20402
rect 19260 20058 19288 20420
rect 19340 20402 19392 20408
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19352 19922 19380 19994
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19444 19530 19472 21490
rect 19536 20058 19564 21966
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 21486 19656 21830
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19720 20874 19748 22066
rect 19812 21554 19840 22374
rect 19904 21962 19932 26182
rect 20916 25294 20944 26726
rect 21192 26518 21220 26930
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 21180 26240 21232 26246
rect 21180 26182 21232 26188
rect 21192 25906 21220 26182
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21192 25362 21220 25842
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 20904 25288 20956 25294
rect 21284 25242 21312 28970
rect 21928 28121 21956 31078
rect 22052 31036 22360 31045
rect 22052 31034 22058 31036
rect 22114 31034 22138 31036
rect 22194 31034 22218 31036
rect 22274 31034 22298 31036
rect 22354 31034 22360 31036
rect 22114 30982 22116 31034
rect 22296 30982 22298 31034
rect 22052 30980 22058 30982
rect 22114 30980 22138 30982
rect 22194 30980 22218 30982
rect 22274 30980 22298 30982
rect 22354 30980 22360 30982
rect 22052 30971 22360 30980
rect 22052 29948 22360 29957
rect 22052 29946 22058 29948
rect 22114 29946 22138 29948
rect 22194 29946 22218 29948
rect 22274 29946 22298 29948
rect 22354 29946 22360 29948
rect 22114 29894 22116 29946
rect 22296 29894 22298 29946
rect 22052 29892 22058 29894
rect 22114 29892 22138 29894
rect 22194 29892 22218 29894
rect 22274 29892 22298 29894
rect 22354 29892 22360 29894
rect 22052 29883 22360 29892
rect 22756 29322 22784 31282
rect 23032 30938 23060 31282
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 23216 30734 23244 31962
rect 23400 31754 23428 32302
rect 23664 31816 23716 31822
rect 23664 31758 23716 31764
rect 23388 31748 23440 31754
rect 23388 31690 23440 31696
rect 23400 30870 23428 31690
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23492 31346 23520 31622
rect 23480 31340 23532 31346
rect 23480 31282 23532 31288
rect 23676 31278 23704 31758
rect 24504 31346 24532 32370
rect 24596 31754 24624 32370
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 25056 31890 25084 32166
rect 25044 31884 25096 31890
rect 25044 31826 25096 31832
rect 25136 31884 25188 31890
rect 25136 31826 25188 31832
rect 24596 31726 24808 31754
rect 24780 31686 24808 31726
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 23664 31272 23716 31278
rect 23664 31214 23716 31220
rect 23388 30864 23440 30870
rect 23388 30806 23440 30812
rect 23676 30802 23704 31214
rect 23664 30796 23716 30802
rect 23664 30738 23716 30744
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23216 29782 23244 30670
rect 23204 29776 23256 29782
rect 23204 29718 23256 29724
rect 24504 29560 24532 31282
rect 24676 30252 24728 30258
rect 24676 30194 24728 30200
rect 24584 29572 24636 29578
rect 24504 29532 24584 29560
rect 24584 29514 24636 29520
rect 22756 29294 22876 29322
rect 22848 29170 22876 29294
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22836 29164 22888 29170
rect 22836 29106 22888 29112
rect 23388 29164 23440 29170
rect 23388 29106 23440 29112
rect 22052 28860 22360 28869
rect 22052 28858 22058 28860
rect 22114 28858 22138 28860
rect 22194 28858 22218 28860
rect 22274 28858 22298 28860
rect 22354 28858 22360 28860
rect 22114 28806 22116 28858
rect 22296 28806 22298 28858
rect 22052 28804 22058 28806
rect 22114 28804 22138 28806
rect 22194 28804 22218 28806
rect 22274 28804 22298 28806
rect 22354 28804 22360 28806
rect 22052 28795 22360 28804
rect 22388 28218 22416 29106
rect 22468 29028 22520 29034
rect 22468 28970 22520 28976
rect 22480 28218 22508 28970
rect 22756 28422 22784 29106
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22376 28212 22428 28218
rect 22376 28154 22428 28160
rect 22468 28212 22520 28218
rect 22468 28154 22520 28160
rect 21914 28112 21970 28121
rect 21914 28047 21970 28056
rect 22284 28076 22336 28082
rect 21928 27334 21956 28047
rect 22284 28018 22336 28024
rect 22296 27962 22324 28018
rect 22296 27934 22416 27962
rect 22052 27772 22360 27781
rect 22052 27770 22058 27772
rect 22114 27770 22138 27772
rect 22194 27770 22218 27772
rect 22274 27770 22298 27772
rect 22354 27770 22360 27772
rect 22114 27718 22116 27770
rect 22296 27718 22298 27770
rect 22052 27716 22058 27718
rect 22114 27716 22138 27718
rect 22194 27716 22218 27718
rect 22274 27716 22298 27718
rect 22354 27716 22360 27718
rect 22052 27707 22360 27716
rect 22388 27674 22416 27934
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 22376 27328 22428 27334
rect 22376 27270 22428 27276
rect 21928 25974 21956 27270
rect 22052 26684 22360 26693
rect 22052 26682 22058 26684
rect 22114 26682 22138 26684
rect 22194 26682 22218 26684
rect 22274 26682 22298 26684
rect 22354 26682 22360 26684
rect 22114 26630 22116 26682
rect 22296 26630 22298 26682
rect 22052 26628 22058 26630
rect 22114 26628 22138 26630
rect 22194 26628 22218 26630
rect 22274 26628 22298 26630
rect 22354 26628 22360 26630
rect 22052 26619 22360 26628
rect 21916 25968 21968 25974
rect 21916 25910 21968 25916
rect 22388 25906 22416 27270
rect 22756 26518 22784 28358
rect 22848 28014 22876 28494
rect 22836 28008 22888 28014
rect 22836 27950 22888 27956
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22052 25596 22360 25605
rect 22052 25594 22058 25596
rect 22114 25594 22138 25596
rect 22194 25594 22218 25596
rect 22274 25594 22298 25596
rect 22354 25594 22360 25596
rect 22114 25542 22116 25594
rect 22296 25542 22298 25594
rect 22052 25540 22058 25542
rect 22114 25540 22138 25542
rect 22194 25540 22218 25542
rect 22274 25540 22298 25542
rect 22354 25540 22360 25542
rect 22052 25531 22360 25540
rect 20904 25230 20956 25236
rect 21088 25220 21140 25226
rect 21088 25162 21140 25168
rect 21192 25214 21312 25242
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 23730 20484 24550
rect 20640 23866 20668 24822
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 21008 24410 21036 24754
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 21100 24274 21128 25162
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20916 23882 20944 24210
rect 20628 23860 20680 23866
rect 20916 23854 21036 23882
rect 20628 23802 20680 23808
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 19996 22642 20024 23190
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19996 22234 20024 22578
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19892 21956 19944 21962
rect 19892 21898 19944 21904
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 19892 21344 19944 21350
rect 19892 21286 19944 21292
rect 19798 21040 19854 21049
rect 19904 21010 19932 21286
rect 19996 21010 20024 22170
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 19798 20975 19854 20984
rect 19892 21004 19944 21010
rect 19812 20942 19840 20975
rect 19892 20946 19944 20952
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19904 20890 19932 20946
rect 19708 20868 19760 20874
rect 19904 20862 20024 20890
rect 19708 20810 19760 20816
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19352 19502 19472 19530
rect 19536 19514 19564 19790
rect 19628 19786 19656 20538
rect 19720 20466 19748 20810
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19812 20398 19840 20538
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19524 19508 19576 19514
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19352 18970 19380 19502
rect 19524 19450 19576 19456
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19444 18766 19472 19382
rect 19628 18970 19656 19722
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 17066 19288 17614
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19260 16250 19288 16458
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19352 15094 19380 18634
rect 19444 17338 19472 18702
rect 19720 18698 19748 20198
rect 19812 19514 19840 20334
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19800 19508 19852 19514
rect 19800 19450 19852 19456
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19524 17060 19576 17066
rect 19524 17002 19576 17008
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19444 15892 19472 16730
rect 19536 16590 19564 17002
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 16250 19564 16526
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19628 16046 19656 18566
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19444 15864 19564 15892
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19352 14346 19380 15030
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19444 14006 19472 14554
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18340 12374 18368 12718
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18432 11218 18460 11630
rect 18524 11626 18552 13194
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12170 18736 12786
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 17831 9820 18139 9829
rect 17831 9818 17837 9820
rect 17893 9818 17917 9820
rect 17973 9818 17997 9820
rect 18053 9818 18077 9820
rect 18133 9818 18139 9820
rect 17893 9766 17895 9818
rect 18075 9766 18077 9818
rect 17831 9764 17837 9766
rect 17893 9764 17917 9766
rect 17973 9764 17997 9766
rect 18053 9764 18077 9766
rect 18133 9764 18139 9766
rect 17831 9755 18139 9764
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17236 8894 17356 8922
rect 17420 8906 17448 9318
rect 17408 8900 17460 8906
rect 17236 8838 17264 8894
rect 17408 8842 17460 8848
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 6798 17264 8774
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17328 7546 17356 8502
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17420 5234 17448 7482
rect 17512 6730 17540 9590
rect 18800 9586 18828 12174
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17696 8634 17724 9454
rect 17788 8838 17816 9522
rect 17880 8906 17908 9522
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17831 8732 18139 8741
rect 17831 8730 17837 8732
rect 17893 8730 17917 8732
rect 17973 8730 17997 8732
rect 18053 8730 18077 8732
rect 18133 8730 18139 8732
rect 17893 8678 17895 8730
rect 18075 8678 18077 8730
rect 17831 8676 17837 8678
rect 17893 8676 17917 8678
rect 17973 8676 17997 8678
rect 18053 8676 18077 8678
rect 18133 8676 18139 8678
rect 17831 8667 18139 8676
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7478 17632 7686
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17696 7410 17724 8570
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 8090 18276 8434
rect 18340 8430 18368 9386
rect 18524 9382 18552 9522
rect 19260 9518 19288 10066
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19352 9382 19380 9522
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 18524 8566 18552 9318
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 17831 7644 18139 7653
rect 17831 7642 17837 7644
rect 17893 7642 17917 7644
rect 17973 7642 17997 7644
rect 18053 7642 18077 7644
rect 18133 7642 18139 7644
rect 17893 7590 17895 7642
rect 18075 7590 18077 7642
rect 17831 7588 17837 7590
rect 17893 7588 17917 7590
rect 17973 7588 17997 7590
rect 18053 7588 18077 7590
rect 18133 7588 18139 7590
rect 17831 7579 18139 7588
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17880 6934 17908 7346
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17880 6798 17908 6870
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17831 6556 18139 6565
rect 17831 6554 17837 6556
rect 17893 6554 17917 6556
rect 17973 6554 17997 6556
rect 18053 6554 18077 6556
rect 18133 6554 18139 6556
rect 17893 6502 17895 6554
rect 18075 6502 18077 6554
rect 17831 6500 17837 6502
rect 17893 6500 17917 6502
rect 17973 6500 17997 6502
rect 18053 6500 18077 6502
rect 18133 6500 18139 6502
rect 17831 6491 18139 6500
rect 17831 5468 18139 5477
rect 17831 5466 17837 5468
rect 17893 5466 17917 5468
rect 17973 5466 17997 5468
rect 18053 5466 18077 5468
rect 18133 5466 18139 5468
rect 17893 5414 17895 5466
rect 18075 5414 18077 5466
rect 17831 5412 17837 5414
rect 17893 5412 17917 5414
rect 17973 5412 17997 5414
rect 18053 5412 18077 5414
rect 18133 5412 18139 5414
rect 17831 5403 18139 5412
rect 18248 5302 18276 8026
rect 18340 6662 18368 8366
rect 18524 8294 18552 8502
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 19444 7206 19472 13942
rect 19536 12434 19564 15864
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19628 14278 19656 14826
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19720 14414 19748 14758
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19628 12918 19656 14214
rect 19720 13938 19748 14350
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19812 13326 19840 14214
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19812 12442 19840 12786
rect 19800 12436 19852 12442
rect 19536 12406 19656 12434
rect 19628 12238 19656 12406
rect 19800 12378 19852 12384
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19524 11280 19576 11286
rect 19904 11234 19932 19654
rect 19996 15570 20024 20862
rect 20088 20058 20116 22034
rect 20456 21622 20484 23666
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20272 20466 20484 20482
rect 20272 20460 20496 20466
rect 20272 20454 20444 20460
rect 20272 20330 20300 20454
rect 20444 20402 20496 20408
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 20088 18630 20116 19722
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 11694 20024 12582
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19524 11222 19576 11228
rect 19536 9654 19564 11222
rect 19812 11206 19932 11234
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19812 9450 19840 11206
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 9450 19932 11086
rect 19996 10742 20024 11630
rect 20088 11150 20116 15846
rect 20180 14074 20208 19790
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20364 15026 20392 18158
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 16590 20484 16934
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20548 16250 20576 22578
rect 20732 22030 20760 23734
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23118 20852 23598
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 19922 20668 20402
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20180 12102 20208 14010
rect 20260 12436 20312 12442
rect 20364 12434 20392 14962
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14006 20484 14758
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20548 13394 20576 16050
rect 20824 15502 20852 19722
rect 20916 18766 20944 23666
rect 21008 22642 21036 23854
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21192 21010 21220 25214
rect 22572 25158 22600 26250
rect 23400 25838 23428 29106
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23584 28150 23612 28494
rect 23572 28144 23624 28150
rect 23572 28086 23624 28092
rect 24596 27606 24624 29514
rect 24688 28558 24716 30194
rect 24780 29646 24808 31622
rect 25148 31482 25176 31826
rect 26608 31816 26660 31822
rect 26608 31758 26660 31764
rect 26272 31580 26580 31589
rect 26272 31578 26278 31580
rect 26334 31578 26358 31580
rect 26414 31578 26438 31580
rect 26494 31578 26518 31580
rect 26574 31578 26580 31580
rect 26334 31526 26336 31578
rect 26516 31526 26518 31578
rect 26272 31524 26278 31526
rect 26334 31524 26358 31526
rect 26414 31524 26438 31526
rect 26494 31524 26518 31526
rect 26574 31524 26580 31526
rect 26272 31515 26580 31524
rect 26620 31482 26648 31758
rect 27724 31754 27752 32370
rect 26700 31748 26752 31754
rect 26700 31690 26752 31696
rect 27712 31748 27764 31754
rect 27712 31690 27764 31696
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25228 31476 25280 31482
rect 25228 31418 25280 31424
rect 25780 31476 25832 31482
rect 25780 31418 25832 31424
rect 26608 31476 26660 31482
rect 26608 31418 26660 31424
rect 25240 31346 25268 31418
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25044 31272 25096 31278
rect 25332 31226 25360 31282
rect 25044 31214 25096 31220
rect 25056 30734 25084 31214
rect 25240 31198 25360 31226
rect 25240 30802 25268 31198
rect 25228 30796 25280 30802
rect 25228 30738 25280 30744
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 25056 30190 25084 30670
rect 25240 30258 25268 30738
rect 25608 30734 25636 31282
rect 25792 31278 25820 31418
rect 26712 31346 26740 31690
rect 26700 31340 26752 31346
rect 26700 31282 26752 31288
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25596 30728 25648 30734
rect 25596 30670 25648 30676
rect 25608 30274 25636 30670
rect 25608 30258 25728 30274
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 25228 30252 25280 30258
rect 25608 30252 25740 30258
rect 25608 30246 25688 30252
rect 25228 30194 25280 30200
rect 25688 30194 25740 30200
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 25056 29850 25084 30126
rect 25148 29850 25176 30194
rect 25044 29844 25096 29850
rect 25044 29786 25096 29792
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24676 27668 24728 27674
rect 24676 27610 24728 27616
rect 24584 27600 24636 27606
rect 24584 27542 24636 27548
rect 24584 26308 24636 26314
rect 24584 26250 24636 26256
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 24596 25294 24624 26250
rect 24688 25906 24716 27610
rect 24780 26994 24808 29582
rect 24858 28112 24914 28121
rect 25148 28098 25176 29786
rect 25240 29238 25268 30194
rect 25792 29458 25820 31214
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26068 30734 26096 31078
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 26068 30394 26096 30670
rect 26272 30492 26580 30501
rect 26272 30490 26278 30492
rect 26334 30490 26358 30492
rect 26414 30490 26438 30492
rect 26494 30490 26518 30492
rect 26574 30490 26580 30492
rect 26334 30438 26336 30490
rect 26516 30438 26518 30490
rect 26272 30436 26278 30438
rect 26334 30436 26358 30438
rect 26414 30436 26438 30438
rect 26494 30436 26518 30438
rect 26574 30436 26580 30438
rect 26272 30427 26580 30436
rect 26056 30388 26108 30394
rect 26056 30330 26108 30336
rect 25700 29430 25820 29458
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 24858 28047 24860 28056
rect 24912 28047 24914 28056
rect 25056 28070 25176 28098
rect 25700 28082 25728 29430
rect 26272 29404 26580 29413
rect 26272 29402 26278 29404
rect 26334 29402 26358 29404
rect 26414 29402 26438 29404
rect 26494 29402 26518 29404
rect 26574 29402 26580 29404
rect 26334 29350 26336 29402
rect 26516 29350 26518 29402
rect 26272 29348 26278 29350
rect 26334 29348 26358 29350
rect 26414 29348 26438 29350
rect 26494 29348 26518 29350
rect 26574 29348 26580 29350
rect 26272 29339 26580 29348
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25688 28076 25740 28082
rect 24860 28018 24912 28024
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24872 26382 24900 28018
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 25056 26042 25084 28070
rect 25688 28018 25740 28024
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25148 26994 25176 27950
rect 25700 27554 25728 28018
rect 25792 28014 25820 29106
rect 26712 28626 26740 31282
rect 26976 30660 27028 30666
rect 26976 30602 27028 30608
rect 27620 30660 27672 30666
rect 27620 30602 27672 30608
rect 26988 30258 27016 30602
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 26988 29646 27016 30194
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27160 29708 27212 29714
rect 27160 29650 27212 29656
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26700 28620 26752 28626
rect 26700 28562 26752 28568
rect 26272 28316 26580 28325
rect 26272 28314 26278 28316
rect 26334 28314 26358 28316
rect 26414 28314 26438 28316
rect 26494 28314 26518 28316
rect 26574 28314 26580 28316
rect 26334 28262 26336 28314
rect 26516 28262 26518 28314
rect 26272 28260 26278 28262
rect 26334 28260 26358 28262
rect 26414 28260 26438 28262
rect 26494 28260 26518 28262
rect 26574 28260 26580 28262
rect 26272 28251 26580 28260
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 25516 27526 25728 27554
rect 25516 27130 25544 27526
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25596 27396 25648 27402
rect 25596 27338 25648 27344
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 25504 27124 25556 27130
rect 25504 27066 25556 27072
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25148 26586 25176 26930
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 24676 25900 24728 25906
rect 25056 25888 25084 25978
rect 25056 25860 25176 25888
rect 24676 25842 24728 25848
rect 24688 25294 24716 25842
rect 25044 25764 25096 25770
rect 25044 25706 25096 25712
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24676 25288 24728 25294
rect 24676 25230 24728 25236
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22100 24880 22152 24886
rect 22100 24822 22152 24828
rect 21548 24812 21600 24818
rect 21548 24754 21600 24760
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21284 24206 21312 24618
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21284 21146 21312 24142
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21100 19854 21128 20402
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21376 19990 21404 20266
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 16114 20944 17478
rect 21008 17202 21036 19110
rect 21560 17814 21588 24754
rect 22112 24732 22140 24822
rect 22192 24744 22244 24750
rect 22112 24704 22192 24732
rect 22192 24686 22244 24692
rect 22052 24508 22360 24517
rect 22052 24506 22058 24508
rect 22114 24506 22138 24508
rect 22194 24506 22218 24508
rect 22274 24506 22298 24508
rect 22354 24506 22360 24508
rect 22114 24454 22116 24506
rect 22296 24454 22298 24506
rect 22052 24452 22058 24454
rect 22114 24452 22138 24454
rect 22194 24452 22218 24454
rect 22274 24452 22298 24454
rect 22354 24452 22360 24454
rect 22052 24443 22360 24452
rect 21916 23792 21968 23798
rect 21916 23734 21968 23740
rect 21928 23322 21956 23734
rect 22052 23420 22360 23429
rect 22052 23418 22058 23420
rect 22114 23418 22138 23420
rect 22194 23418 22218 23420
rect 22274 23418 22298 23420
rect 22354 23418 22360 23420
rect 22114 23366 22116 23418
rect 22296 23366 22298 23418
rect 22052 23364 22058 23366
rect 22114 23364 22138 23366
rect 22194 23364 22218 23366
rect 22274 23364 22298 23366
rect 22354 23364 22360 23366
rect 22052 23355 22360 23364
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21744 19786 21772 20198
rect 21732 19780 21784 19786
rect 21732 19722 21784 19728
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21560 17610 21588 17750
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21008 16794 21036 17138
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21192 16454 21220 17206
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16182 21220 16390
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20364 12406 20484 12434
rect 20260 12378 20312 12384
rect 20272 12170 20300 12378
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11150 20208 12038
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 20364 9654 20392 12174
rect 20456 11014 20484 12406
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20548 11354 20576 12174
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20456 9926 20484 10950
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19536 7546 19564 8910
rect 19904 8430 19932 8910
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19720 6798 19748 8298
rect 20364 7002 20392 9590
rect 20548 9382 20576 11018
rect 20640 10062 20668 14010
rect 20732 12170 20760 14486
rect 20824 13870 20852 14962
rect 20916 14822 20944 14962
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20812 12436 20864 12442
rect 20916 12434 20944 14758
rect 21008 14414 21036 15302
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21100 12782 21128 16050
rect 21836 15162 21864 22578
rect 22052 22332 22360 22341
rect 22052 22330 22058 22332
rect 22114 22330 22138 22332
rect 22194 22330 22218 22332
rect 22274 22330 22298 22332
rect 22354 22330 22360 22332
rect 22114 22278 22116 22330
rect 22296 22278 22298 22330
rect 22052 22276 22058 22278
rect 22114 22276 22138 22278
rect 22194 22276 22218 22278
rect 22274 22276 22298 22278
rect 22354 22276 22360 22278
rect 22052 22267 22360 22276
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21554 22324 21830
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22052 21244 22360 21253
rect 22052 21242 22058 21244
rect 22114 21242 22138 21244
rect 22194 21242 22218 21244
rect 22274 21242 22298 21244
rect 22354 21242 22360 21244
rect 22114 21190 22116 21242
rect 22296 21190 22298 21242
rect 22052 21188 22058 21190
rect 22114 21188 22138 21190
rect 22194 21188 22218 21190
rect 22274 21188 22298 21190
rect 22354 21188 22360 21190
rect 22052 21179 22360 21188
rect 22388 20534 22416 21422
rect 22572 20942 22600 25094
rect 23492 24342 23520 25230
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23584 24138 23612 24890
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23572 24132 23624 24138
rect 23572 24074 23624 24080
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22376 20528 22428 20534
rect 22376 20470 22428 20476
rect 22572 20398 22600 20742
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22052 20156 22360 20165
rect 22052 20154 22058 20156
rect 22114 20154 22138 20156
rect 22194 20154 22218 20156
rect 22274 20154 22298 20156
rect 22354 20154 22360 20156
rect 22114 20102 22116 20154
rect 22296 20102 22298 20154
rect 22052 20100 22058 20102
rect 22114 20100 22138 20102
rect 22194 20100 22218 20102
rect 22274 20100 22298 20102
rect 22354 20100 22360 20102
rect 22052 20091 22360 20100
rect 22052 19068 22360 19077
rect 22052 19066 22058 19068
rect 22114 19066 22138 19068
rect 22194 19066 22218 19068
rect 22274 19066 22298 19068
rect 22354 19066 22360 19068
rect 22114 19014 22116 19066
rect 22296 19014 22298 19066
rect 22052 19012 22058 19014
rect 22114 19012 22138 19014
rect 22194 19012 22218 19014
rect 22274 19012 22298 19014
rect 22354 19012 22360 19014
rect 22052 19003 22360 19012
rect 22052 17980 22360 17989
rect 22052 17978 22058 17980
rect 22114 17978 22138 17980
rect 22194 17978 22218 17980
rect 22274 17978 22298 17980
rect 22354 17978 22360 17980
rect 22114 17926 22116 17978
rect 22296 17926 22298 17978
rect 22052 17924 22058 17926
rect 22114 17924 22138 17926
rect 22194 17924 22218 17926
rect 22274 17924 22298 17926
rect 22354 17924 22360 17926
rect 22052 17915 22360 17924
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22052 16892 22360 16901
rect 22052 16890 22058 16892
rect 22114 16890 22138 16892
rect 22194 16890 22218 16892
rect 22274 16890 22298 16892
rect 22354 16890 22360 16892
rect 22114 16838 22116 16890
rect 22296 16838 22298 16890
rect 22052 16836 22058 16838
rect 22114 16836 22138 16838
rect 22194 16836 22218 16838
rect 22274 16836 22298 16838
rect 22354 16836 22360 16838
rect 22052 16827 22360 16836
rect 22468 16516 22520 16522
rect 22468 16458 22520 16464
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15638 21956 16050
rect 22052 15804 22360 15813
rect 22052 15802 22058 15804
rect 22114 15802 22138 15804
rect 22194 15802 22218 15804
rect 22274 15802 22298 15804
rect 22354 15802 22360 15804
rect 22114 15750 22116 15802
rect 22296 15750 22298 15802
rect 22052 15748 22058 15750
rect 22114 15748 22138 15750
rect 22194 15748 22218 15750
rect 22274 15748 22298 15750
rect 22354 15748 22360 15750
rect 22052 15739 22360 15748
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20864 12406 20944 12434
rect 20812 12378 20864 12384
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20640 9586 20668 9862
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20456 8974 20484 9318
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20456 8498 20484 8774
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 7478 20484 7686
rect 20548 7546 20576 8434
rect 20732 7886 20760 12106
rect 20824 11234 20852 12378
rect 21100 12306 21128 12582
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21192 11880 21220 14214
rect 21270 12472 21326 12481
rect 21928 12442 21956 15030
rect 22296 14822 22324 15098
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22052 14716 22360 14725
rect 22052 14714 22058 14716
rect 22114 14714 22138 14716
rect 22194 14714 22218 14716
rect 22274 14714 22298 14716
rect 22354 14714 22360 14716
rect 22114 14662 22116 14714
rect 22296 14662 22298 14714
rect 22052 14660 22058 14662
rect 22114 14660 22138 14662
rect 22194 14660 22218 14662
rect 22274 14660 22298 14662
rect 22354 14660 22360 14662
rect 22052 14651 22360 14660
rect 22388 14618 22416 15370
rect 22480 15026 22508 16458
rect 22572 15570 22600 17070
rect 22664 16250 22692 22102
rect 22756 20602 22784 23054
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 23032 22234 23060 22374
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23584 22094 23612 24074
rect 23676 23730 23704 24822
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23768 24342 23796 24754
rect 23756 24336 23808 24342
rect 23756 24278 23808 24284
rect 24688 24070 24716 25230
rect 25056 24682 25084 25706
rect 25148 25226 25176 25860
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25148 24954 25176 25162
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25240 24818 25268 27066
rect 25608 26994 25636 27338
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 26444 25556 26450
rect 25504 26386 25556 26392
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25332 24818 25360 26318
rect 25516 25974 25544 26386
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 25504 25968 25556 25974
rect 25504 25910 25556 25916
rect 25608 25498 25636 26318
rect 25700 26042 25728 27406
rect 25792 27334 25820 27950
rect 25872 27940 25924 27946
rect 25872 27882 25924 27888
rect 25884 27538 25912 27882
rect 25872 27532 25924 27538
rect 25872 27474 25924 27480
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25884 26994 25912 27474
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27062 26188 27406
rect 26252 27402 26280 27950
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26272 27228 26580 27237
rect 26272 27226 26278 27228
rect 26334 27226 26358 27228
rect 26414 27226 26438 27228
rect 26494 27226 26518 27228
rect 26574 27226 26580 27228
rect 26334 27174 26336 27226
rect 26516 27174 26518 27226
rect 26272 27172 26278 27174
rect 26334 27172 26358 27174
rect 26414 27172 26438 27174
rect 26494 27172 26518 27174
rect 26574 27172 26580 27174
rect 26272 27163 26580 27172
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 25688 26036 25740 26042
rect 25688 25978 25740 25984
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25044 24676 25096 24682
rect 25044 24618 25096 24624
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24688 23730 24716 24006
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24964 23186 24992 23462
rect 24952 23180 25004 23186
rect 24952 23122 25004 23128
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24952 22976 25004 22982
rect 25056 22964 25084 24618
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25228 24404 25280 24410
rect 25228 24346 25280 24352
rect 25240 24206 25268 24346
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25136 24132 25188 24138
rect 25136 24074 25188 24080
rect 25004 22936 25084 22964
rect 24952 22918 25004 22924
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24584 22432 24636 22438
rect 24584 22374 24636 22380
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23492 22066 23612 22094
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22112 13977 22140 14282
rect 22098 13968 22154 13977
rect 22204 13938 22232 14282
rect 22480 13938 22508 14826
rect 22098 13903 22154 13912
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22204 13818 22232 13874
rect 22204 13790 22416 13818
rect 22052 13628 22360 13637
rect 22052 13626 22058 13628
rect 22114 13626 22138 13628
rect 22194 13626 22218 13628
rect 22274 13626 22298 13628
rect 22354 13626 22360 13628
rect 22114 13574 22116 13626
rect 22296 13574 22298 13626
rect 22052 13572 22058 13574
rect 22114 13572 22138 13574
rect 22194 13572 22218 13574
rect 22274 13572 22298 13574
rect 22354 13572 22360 13574
rect 22052 13563 22360 13572
rect 22388 13394 22416 13790
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22296 12730 22324 12786
rect 22296 12702 22416 12730
rect 22052 12540 22360 12549
rect 22052 12538 22058 12540
rect 22114 12538 22138 12540
rect 22194 12538 22218 12540
rect 22274 12538 22298 12540
rect 22354 12538 22360 12540
rect 22114 12486 22116 12538
rect 22296 12486 22298 12538
rect 22052 12484 22058 12486
rect 22114 12484 22138 12486
rect 22194 12484 22218 12486
rect 22274 12484 22298 12486
rect 22354 12484 22360 12486
rect 22052 12475 22360 12484
rect 21270 12407 21326 12416
rect 21916 12436 21968 12442
rect 21284 12170 21312 12407
rect 21916 12378 21968 12384
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 21008 11852 21220 11880
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 11354 20944 11698
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20824 11206 20944 11234
rect 20916 11082 20944 11206
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20824 9586 20852 9862
rect 20916 9586 20944 11018
rect 21008 10690 21036 11852
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21100 11286 21128 11698
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 21180 11144 21232 11150
rect 21284 11132 21312 12106
rect 21364 11620 21416 11626
rect 21364 11562 21416 11568
rect 21376 11150 21404 11562
rect 22112 11558 22140 12106
rect 22204 11898 22232 12106
rect 22388 11898 22416 12702
rect 22480 12238 22508 13874
rect 22940 12986 22968 21966
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23124 21622 23152 21898
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23216 19922 23244 21422
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23216 19378 23244 19858
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23400 19310 23428 20810
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23492 18766 23520 22066
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23584 21146 23612 21422
rect 23860 21350 23888 22170
rect 24596 22030 24624 22374
rect 24780 22234 24808 22510
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23952 20942 23980 21286
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23124 17134 23152 18158
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22572 12594 22600 12786
rect 22572 12566 22692 12594
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22480 11830 22508 12174
rect 22664 12102 22692 12566
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22756 11880 22784 12378
rect 22940 12170 22968 12786
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23032 12442 23060 12718
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23124 12374 23152 16050
rect 23216 14890 23244 17274
rect 23584 17270 23612 18566
rect 23860 18222 23888 18702
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23572 17264 23624 17270
rect 23572 17206 23624 17212
rect 23860 17202 23888 18158
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 24412 16998 24440 18566
rect 24596 18290 24624 18566
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24780 17814 24808 18702
rect 24872 18290 24900 22918
rect 24964 22166 24992 22918
rect 24952 22160 25004 22166
rect 24952 22102 25004 22108
rect 24952 21888 25004 21894
rect 24952 21830 25004 21836
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24964 21146 24992 21830
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 24964 21010 24992 21082
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18426 24992 18566
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24780 16998 24808 17614
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 23400 15434 23428 16934
rect 24412 16046 24440 16934
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24596 15910 24624 16526
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23388 15156 23440 15162
rect 23492 15144 23520 15438
rect 23440 15116 23520 15144
rect 23388 15098 23440 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 14550 23336 14758
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23400 14346 23428 14962
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 24044 14006 24072 14758
rect 24596 14482 24624 15846
rect 24780 15570 24808 16934
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24872 14414 24900 17478
rect 25056 17202 25084 21830
rect 25148 20942 25176 24074
rect 25240 23798 25268 24142
rect 25320 24064 25372 24070
rect 25320 24006 25372 24012
rect 25228 23792 25280 23798
rect 25228 23734 25280 23740
rect 25332 23186 25360 24006
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 25228 22976 25280 22982
rect 25228 22918 25280 22924
rect 25240 22710 25268 22918
rect 25228 22704 25280 22710
rect 25228 22646 25280 22652
rect 25240 22098 25268 22646
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25976 22030 26004 24550
rect 26160 22574 26188 26862
rect 26620 26602 26648 27814
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 26528 26574 26648 26602
rect 26528 26518 26556 26574
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26528 26382 26556 26454
rect 26516 26376 26568 26382
rect 26608 26376 26660 26382
rect 26516 26318 26568 26324
rect 26606 26344 26608 26353
rect 26660 26344 26662 26353
rect 26606 26279 26662 26288
rect 26608 26240 26660 26246
rect 26608 26182 26660 26188
rect 26272 26140 26580 26149
rect 26272 26138 26278 26140
rect 26334 26138 26358 26140
rect 26414 26138 26438 26140
rect 26494 26138 26518 26140
rect 26574 26138 26580 26140
rect 26334 26086 26336 26138
rect 26516 26086 26518 26138
rect 26272 26084 26278 26086
rect 26334 26084 26358 26086
rect 26414 26084 26438 26086
rect 26494 26084 26518 26086
rect 26574 26084 26580 26086
rect 26272 26075 26580 26084
rect 26516 25900 26568 25906
rect 26620 25888 26648 26182
rect 26568 25860 26648 25888
rect 26516 25842 26568 25848
rect 26528 25226 26556 25842
rect 26712 25838 26740 27270
rect 26792 26512 26844 26518
rect 26792 26454 26844 26460
rect 26700 25832 26752 25838
rect 26700 25774 26752 25780
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 26516 25220 26568 25226
rect 26516 25162 26568 25168
rect 26272 25052 26580 25061
rect 26272 25050 26278 25052
rect 26334 25050 26358 25052
rect 26414 25050 26438 25052
rect 26494 25050 26518 25052
rect 26574 25050 26580 25052
rect 26334 24998 26336 25050
rect 26516 24998 26518 25050
rect 26272 24996 26278 24998
rect 26334 24996 26358 24998
rect 26414 24996 26438 24998
rect 26494 24996 26518 24998
rect 26574 24996 26580 24998
rect 26272 24987 26580 24996
rect 26620 24614 26648 25298
rect 26608 24608 26660 24614
rect 26608 24550 26660 24556
rect 26712 24206 26740 25774
rect 26804 25498 26832 26454
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26272 23964 26580 23973
rect 26272 23962 26278 23964
rect 26334 23962 26358 23964
rect 26414 23962 26438 23964
rect 26494 23962 26518 23964
rect 26574 23962 26580 23964
rect 26334 23910 26336 23962
rect 26516 23910 26518 23962
rect 26272 23908 26278 23910
rect 26334 23908 26358 23910
rect 26414 23908 26438 23910
rect 26494 23908 26518 23910
rect 26574 23908 26580 23910
rect 26272 23899 26580 23908
rect 26272 22876 26580 22885
rect 26272 22874 26278 22876
rect 26334 22874 26358 22876
rect 26414 22874 26438 22876
rect 26494 22874 26518 22876
rect 26574 22874 26580 22876
rect 26334 22822 26336 22874
rect 26516 22822 26518 22874
rect 26272 22820 26278 22822
rect 26334 22820 26358 22822
rect 26414 22820 26438 22822
rect 26494 22820 26518 22822
rect 26574 22820 26580 22822
rect 26272 22811 26580 22820
rect 26988 22574 27016 29582
rect 27172 29170 27200 29650
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 27344 29164 27396 29170
rect 27344 29106 27396 29112
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 27080 27334 27108 28018
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 27080 26586 27108 27270
rect 27264 26994 27292 28358
rect 27356 28150 27384 29106
rect 27344 28144 27396 28150
rect 27344 28086 27396 28092
rect 27448 26994 27476 29990
rect 27540 29646 27568 30194
rect 27632 29646 27660 30602
rect 28092 30326 28120 32370
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 33140 32224 33192 32230
rect 33140 32166 33192 32172
rect 29092 31272 29144 31278
rect 29092 31214 29144 31220
rect 28540 31136 28592 31142
rect 28540 31078 28592 31084
rect 28552 30326 28580 31078
rect 29104 30802 29132 31214
rect 29092 30796 29144 30802
rect 29092 30738 29144 30744
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 28724 30660 28776 30666
rect 28724 30602 28776 30608
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 28540 30320 28592 30326
rect 28540 30262 28592 30268
rect 28736 30258 28764 30602
rect 28724 30252 28776 30258
rect 28724 30194 28776 30200
rect 28632 30184 28684 30190
rect 28632 30126 28684 30132
rect 28080 30116 28132 30122
rect 28080 30058 28132 30064
rect 27528 29640 27580 29646
rect 27528 29582 27580 29588
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27632 29306 27660 29582
rect 27712 29572 27764 29578
rect 27712 29514 27764 29520
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27528 29028 27580 29034
rect 27724 28994 27752 29514
rect 28092 29170 28120 30058
rect 28644 30054 28672 30126
rect 28632 30048 28684 30054
rect 28632 29990 28684 29996
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28368 29306 28396 29582
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 28644 29102 28672 29990
rect 28920 29782 28948 30670
rect 29104 30394 29132 30738
rect 29092 30388 29144 30394
rect 29092 30330 29144 30336
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29184 30252 29236 30258
rect 29184 30194 29236 30200
rect 28908 29776 28960 29782
rect 28908 29718 28960 29724
rect 29012 29714 29040 30194
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 29196 29646 29224 30194
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 29184 29640 29236 29646
rect 29184 29582 29236 29588
rect 28172 29096 28224 29102
rect 28172 29038 28224 29044
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 27528 28970 27580 28976
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27068 26580 27120 26586
rect 27068 26522 27120 26528
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 27080 25158 27108 25774
rect 27172 25770 27200 26318
rect 27264 26042 27292 26930
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 27160 25764 27212 25770
rect 27160 25706 27212 25712
rect 27448 25378 27476 26930
rect 27540 26246 27568 28970
rect 27632 28966 27752 28994
rect 27632 28626 27660 28966
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27632 26926 27660 28562
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27724 27470 27752 28018
rect 27908 27606 27936 28494
rect 27896 27600 27948 27606
rect 27896 27542 27948 27548
rect 28184 27470 28212 29038
rect 28920 28966 28948 29582
rect 29196 29306 29224 29582
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 28908 28960 28960 28966
rect 28908 28902 28960 28908
rect 28920 28762 28948 28902
rect 28908 28756 28960 28762
rect 28908 28698 28960 28704
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 27618 26344 27674 26353
rect 27618 26279 27674 26288
rect 27528 26240 27580 26246
rect 27528 26182 27580 26188
rect 27540 25838 27568 26182
rect 27632 25906 27660 26279
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27356 25350 27476 25378
rect 27356 25294 27384 25350
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 27080 24886 27108 25094
rect 27068 24880 27120 24886
rect 27068 24822 27120 24828
rect 27160 24880 27212 24886
rect 27160 24822 27212 24828
rect 27172 23662 27200 24822
rect 27540 24410 27568 25774
rect 27632 25498 27660 25842
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 28184 24750 28212 27406
rect 28736 27334 28764 28494
rect 29000 28076 29052 28082
rect 29000 28018 29052 28024
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28632 26512 28684 26518
rect 28632 26454 28684 26460
rect 28644 25974 28672 26454
rect 28632 25968 28684 25974
rect 28632 25910 28684 25916
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 28644 23798 28672 25910
rect 28724 24812 28776 24818
rect 28724 24754 28776 24760
rect 28632 23792 28684 23798
rect 28632 23734 28684 23740
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 28736 23254 28764 24754
rect 29012 24342 29040 28018
rect 30012 27872 30064 27878
rect 30012 27814 30064 27820
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29932 26926 29960 27406
rect 30024 26994 30052 27814
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 29920 26920 29972 26926
rect 29920 26862 29972 26868
rect 29092 26308 29144 26314
rect 29092 26250 29144 26256
rect 29104 24818 29132 26250
rect 29932 26042 29960 26862
rect 29920 26036 29972 26042
rect 29920 25978 29972 25984
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 30116 24750 30144 25230
rect 30104 24744 30156 24750
rect 30104 24686 30156 24692
rect 29000 24336 29052 24342
rect 29000 24278 29052 24284
rect 30116 23866 30144 24686
rect 30104 23860 30156 23866
rect 30104 23802 30156 23808
rect 28724 23248 28776 23254
rect 28724 23190 28776 23196
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26976 22432 27028 22438
rect 26976 22374 27028 22380
rect 26988 22098 27016 22374
rect 26148 22094 26200 22098
rect 26148 22092 26372 22094
rect 26200 22066 26372 22092
rect 26148 22034 26200 22040
rect 26344 22030 26372 22066
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26272 21788 26580 21797
rect 26272 21786 26278 21788
rect 26334 21786 26358 21788
rect 26414 21786 26438 21788
rect 26494 21786 26518 21788
rect 26574 21786 26580 21788
rect 26334 21734 26336 21786
rect 26516 21734 26518 21786
rect 26272 21732 26278 21734
rect 26334 21732 26358 21734
rect 26414 21732 26438 21734
rect 26494 21732 26518 21734
rect 26574 21732 26580 21734
rect 26272 21723 26580 21732
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25148 18766 25176 20878
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25240 19446 25268 20742
rect 26272 20700 26580 20709
rect 26272 20698 26278 20700
rect 26334 20698 26358 20700
rect 26414 20698 26438 20700
rect 26494 20698 26518 20700
rect 26574 20698 26580 20700
rect 26334 20646 26336 20698
rect 26516 20646 26518 20698
rect 26272 20644 26278 20646
rect 26334 20644 26358 20646
rect 26414 20644 26438 20646
rect 26494 20644 26518 20646
rect 26574 20644 26580 20646
rect 26272 20635 26580 20644
rect 25872 20392 25924 20398
rect 25872 20334 25924 20340
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25884 18970 25912 20334
rect 26272 19612 26580 19621
rect 26272 19610 26278 19612
rect 26334 19610 26358 19612
rect 26414 19610 26438 19612
rect 26494 19610 26518 19612
rect 26574 19610 26580 19612
rect 26334 19558 26336 19610
rect 26516 19558 26518 19610
rect 26272 19556 26278 19558
rect 26334 19556 26358 19558
rect 26414 19556 26438 19558
rect 26494 19556 26518 19558
rect 26574 19556 26580 19558
rect 26272 19547 26580 19556
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25964 18760 26016 18766
rect 26240 18760 26292 18766
rect 26016 18720 26096 18748
rect 25964 18702 26016 18708
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25700 18426 25728 18634
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 25148 15706 25176 16050
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25148 15162 25176 15370
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24780 14006 24808 14214
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 23296 12708 23348 12714
rect 23296 12650 23348 12656
rect 23112 12368 23164 12374
rect 23112 12310 23164 12316
rect 23308 12238 23336 12650
rect 23388 12436 23440 12442
rect 24596 12434 24624 13874
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 24596 12406 24716 12434
rect 23388 12378 23440 12384
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22836 11892 22888 11898
rect 22756 11852 22836 11880
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22052 11452 22360 11461
rect 22052 11450 22058 11452
rect 22114 11450 22138 11452
rect 22194 11450 22218 11452
rect 22274 11450 22298 11452
rect 22354 11450 22360 11452
rect 22114 11398 22116 11450
rect 22296 11398 22298 11450
rect 22052 11396 22058 11398
rect 22114 11396 22138 11398
rect 22194 11396 22218 11398
rect 22274 11396 22298 11398
rect 22354 11396 22360 11398
rect 22052 11387 22360 11396
rect 21232 11104 21312 11132
rect 21364 11144 21416 11150
rect 21180 11086 21232 11092
rect 21364 11086 21416 11092
rect 21008 10662 21128 10690
rect 21100 10062 21128 10662
rect 22052 10364 22360 10373
rect 22052 10362 22058 10364
rect 22114 10362 22138 10364
rect 22194 10362 22218 10364
rect 22274 10362 22298 10364
rect 22354 10362 22360 10364
rect 22114 10310 22116 10362
rect 22296 10310 22298 10362
rect 22052 10308 22058 10310
rect 22114 10308 22138 10310
rect 22194 10308 22218 10310
rect 22274 10308 22298 10310
rect 22354 10308 22360 10310
rect 22052 10299 22360 10308
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20824 9178 20852 9522
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20916 8634 20944 9522
rect 21008 9042 21036 9590
rect 21100 9450 21128 9998
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20824 7546 20852 7754
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20916 7478 20944 8570
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21008 7546 21036 8502
rect 21100 8498 21128 9386
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21192 8362 21220 9386
rect 22052 9276 22360 9285
rect 22052 9274 22058 9276
rect 22114 9274 22138 9276
rect 22194 9274 22218 9276
rect 22274 9274 22298 9276
rect 22354 9274 22360 9276
rect 22114 9222 22116 9274
rect 22296 9222 22298 9274
rect 22052 9220 22058 9222
rect 22114 9220 22138 9222
rect 22194 9220 22218 9222
rect 22274 9220 22298 9222
rect 22354 9220 22360 9222
rect 22052 9211 22360 9220
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 19536 6254 19564 6734
rect 20732 6390 20760 7142
rect 21008 6458 21036 7482
rect 21284 6866 21312 8366
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21744 7274 21772 8230
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21836 6798 21864 8774
rect 22052 8188 22360 8197
rect 22052 8186 22058 8188
rect 22114 8186 22138 8188
rect 22194 8186 22218 8188
rect 22274 8186 22298 8188
rect 22354 8186 22360 8188
rect 22114 8134 22116 8186
rect 22296 8134 22298 8186
rect 22052 8132 22058 8134
rect 22114 8132 22138 8134
rect 22194 8132 22218 8134
rect 22274 8132 22298 8134
rect 22354 8132 22360 8134
rect 22052 8123 22360 8132
rect 22388 7410 22416 11494
rect 22572 8634 22600 11698
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22052 7100 22360 7109
rect 22052 7098 22058 7100
rect 22114 7098 22138 7100
rect 22194 7098 22218 7100
rect 22274 7098 22298 7100
rect 22354 7098 22360 7100
rect 22114 7046 22116 7098
rect 22296 7046 22298 7098
rect 22052 7044 22058 7046
rect 22114 7044 22138 7046
rect 22194 7044 22218 7046
rect 22274 7044 22298 7046
rect 22354 7044 22360 7046
rect 22052 7035 22360 7044
rect 22664 6866 22692 11698
rect 22756 8566 22784 11852
rect 22836 11834 22888 11840
rect 22940 11744 22968 12106
rect 23020 11756 23072 11762
rect 22940 11716 23020 11744
rect 23020 11698 23072 11704
rect 23400 11558 23428 12378
rect 24688 12306 24716 12406
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24596 11830 24624 12038
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 23848 11688 23900 11694
rect 24688 11642 24716 12242
rect 24780 12102 24808 12854
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24872 12238 24900 12378
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11898 24808 12038
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 23848 11630 23900 11636
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23860 10470 23888 11630
rect 24596 11614 24716 11642
rect 24596 11150 24624 11614
rect 25056 11286 25084 13874
rect 25148 13802 25176 14962
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 10130 23888 10406
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22848 8974 22876 9114
rect 22836 8968 22888 8974
rect 22836 8910 22888 8916
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17420 4622 17448 5170
rect 18432 4622 18460 6122
rect 19536 5370 19564 6190
rect 22664 6186 22692 6802
rect 22848 6662 22876 8910
rect 23676 8906 23704 9454
rect 24596 8974 24624 11086
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10062 24900 11018
rect 25332 10266 25360 18022
rect 25516 10810 25544 18226
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25700 17338 25728 17614
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25792 17270 25820 17478
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25608 14278 25636 17138
rect 25792 14618 25820 17206
rect 26068 17202 26096 18720
rect 26240 18702 26292 18708
rect 26252 18630 26280 18702
rect 27080 18630 27108 21966
rect 27172 21690 27200 22578
rect 27540 21962 27568 23054
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27528 21956 27580 21962
rect 27528 21898 27580 21904
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27632 21486 27660 22986
rect 28000 22642 28028 23054
rect 28276 22710 28304 23054
rect 28540 23044 28592 23050
rect 28540 22986 28592 22992
rect 28264 22704 28316 22710
rect 28264 22646 28316 22652
rect 28552 22642 28580 22986
rect 29736 22976 29788 22982
rect 29736 22918 29788 22924
rect 27988 22636 28040 22642
rect 28540 22636 28592 22642
rect 28040 22596 28212 22624
rect 27988 22578 28040 22584
rect 27988 22500 28040 22506
rect 27988 22442 28040 22448
rect 28000 21554 28028 22442
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27908 20398 27936 21286
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27264 18766 27292 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27356 18834 27384 19110
rect 27712 18896 27764 18902
rect 27712 18838 27764 18844
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26272 18524 26580 18533
rect 26272 18522 26278 18524
rect 26334 18522 26358 18524
rect 26414 18522 26438 18524
rect 26494 18522 26518 18524
rect 26574 18522 26580 18524
rect 26334 18470 26336 18522
rect 26516 18470 26518 18522
rect 26272 18468 26278 18470
rect 26334 18468 26358 18470
rect 26414 18468 26438 18470
rect 26494 18468 26518 18470
rect 26574 18468 26580 18470
rect 26272 18459 26580 18468
rect 27264 18222 27292 18702
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27724 17678 27752 18838
rect 27908 18766 27936 19314
rect 27896 18760 27948 18766
rect 27896 18702 27948 18708
rect 27908 17746 27936 18702
rect 28000 17882 28028 20402
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 26272 17436 26580 17445
rect 26272 17434 26278 17436
rect 26334 17434 26358 17436
rect 26414 17434 26438 17436
rect 26494 17434 26518 17436
rect 26574 17434 26580 17436
rect 26334 17382 26336 17434
rect 26516 17382 26518 17434
rect 26272 17380 26278 17382
rect 26334 17380 26358 17382
rect 26414 17380 26438 17382
rect 26494 17380 26518 17382
rect 26574 17380 26580 17382
rect 26272 17371 26580 17380
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26068 16658 26096 17138
rect 26620 17134 26648 17546
rect 26608 17128 26660 17134
rect 26608 17070 26660 17076
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25976 16182 26004 16390
rect 26068 16250 26096 16458
rect 26056 16244 26108 16250
rect 26056 16186 26108 16192
rect 25964 16176 26016 16182
rect 25964 16118 26016 16124
rect 26160 16130 26188 16730
rect 26272 16348 26580 16357
rect 26272 16346 26278 16348
rect 26334 16346 26358 16348
rect 26414 16346 26438 16348
rect 26494 16346 26518 16348
rect 26574 16346 26580 16348
rect 26334 16294 26336 16346
rect 26516 16294 26518 16346
rect 26272 16292 26278 16294
rect 26334 16292 26358 16294
rect 26414 16292 26438 16294
rect 26494 16292 26518 16294
rect 26574 16292 26580 16294
rect 26272 16283 26580 16292
rect 26160 16114 26280 16130
rect 26620 16114 26648 17070
rect 26700 16516 26752 16522
rect 26700 16458 26752 16464
rect 26160 16108 26292 16114
rect 26160 16102 26240 16108
rect 26240 16050 26292 16056
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25780 14612 25832 14618
rect 25780 14554 25832 14560
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 26068 13326 26096 15642
rect 26272 15260 26580 15269
rect 26272 15258 26278 15260
rect 26334 15258 26358 15260
rect 26414 15258 26438 15260
rect 26494 15258 26518 15260
rect 26574 15258 26580 15260
rect 26334 15206 26336 15258
rect 26516 15206 26518 15258
rect 26272 15204 26278 15206
rect 26334 15204 26358 15206
rect 26414 15204 26438 15206
rect 26494 15204 26518 15206
rect 26574 15204 26580 15206
rect 26272 15195 26580 15204
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26436 14414 26464 14894
rect 26620 14618 26648 16050
rect 26712 15094 26740 16458
rect 27724 16232 27752 17614
rect 27816 17338 27844 17614
rect 27804 17332 27856 17338
rect 27804 17274 27856 17280
rect 27724 16204 27844 16232
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 26700 15088 26752 15094
rect 26700 15030 26752 15036
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26272 14172 26580 14181
rect 26272 14170 26278 14172
rect 26334 14170 26358 14172
rect 26414 14170 26438 14172
rect 26494 14170 26518 14172
rect 26574 14170 26580 14172
rect 26334 14118 26336 14170
rect 26516 14118 26518 14170
rect 26272 14116 26278 14118
rect 26334 14116 26358 14118
rect 26414 14116 26438 14118
rect 26494 14116 26518 14118
rect 26574 14116 26580 14118
rect 26272 14107 26580 14116
rect 26620 13870 26648 14554
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26988 13530 27016 14350
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 26272 13084 26580 13093
rect 26272 13082 26278 13084
rect 26334 13082 26358 13084
rect 26414 13082 26438 13084
rect 26494 13082 26518 13084
rect 26574 13082 26580 13084
rect 26334 13030 26336 13082
rect 26516 13030 26518 13082
rect 26272 13028 26278 13030
rect 26334 13028 26358 13030
rect 26414 13028 26438 13030
rect 26494 13028 26518 13030
rect 26574 13028 26580 13030
rect 26272 13019 26580 13028
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 26272 11996 26580 12005
rect 26272 11994 26278 11996
rect 26334 11994 26358 11996
rect 26414 11994 26438 11996
rect 26494 11994 26518 11996
rect 26574 11994 26580 11996
rect 26334 11942 26336 11994
rect 26516 11942 26518 11994
rect 26272 11940 26278 11942
rect 26334 11940 26358 11942
rect 26414 11940 26438 11942
rect 26494 11940 26518 11942
rect 26574 11940 26580 11942
rect 26272 11931 26580 11940
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25780 11280 25832 11286
rect 25780 11222 25832 11228
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 25700 9654 25728 10610
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23676 8634 23704 8842
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24044 7886 24072 8298
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7478 23428 7686
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22652 6180 22704 6186
rect 22652 6122 22704 6128
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19996 4622 20024 6054
rect 22052 6012 22360 6021
rect 22052 6010 22058 6012
rect 22114 6010 22138 6012
rect 22194 6010 22218 6012
rect 22274 6010 22298 6012
rect 22354 6010 22360 6012
rect 22114 5958 22116 6010
rect 22296 5958 22298 6010
rect 22052 5956 22058 5958
rect 22114 5956 22138 5958
rect 22194 5956 22218 5958
rect 22274 5956 22298 5958
rect 22354 5956 22360 5958
rect 22052 5947 22360 5956
rect 23400 5302 23428 7414
rect 24596 7342 24624 8910
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8566 25084 8774
rect 25700 8634 25728 9590
rect 25792 8838 25820 11222
rect 25976 10674 26004 11698
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 26068 11150 26096 11494
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26160 10674 26188 11154
rect 26272 10908 26580 10917
rect 26272 10906 26278 10908
rect 26334 10906 26358 10908
rect 26414 10906 26438 10908
rect 26494 10906 26518 10908
rect 26574 10906 26580 10908
rect 26334 10854 26336 10906
rect 26516 10854 26518 10906
rect 26272 10852 26278 10854
rect 26334 10852 26358 10854
rect 26414 10852 26438 10854
rect 26494 10852 26518 10854
rect 26574 10852 26580 10854
rect 26272 10843 26580 10852
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 25792 8498 25820 8774
rect 25884 8634 25912 10610
rect 25976 10470 26004 10610
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 26160 10266 26188 10610
rect 26252 10266 26280 10610
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 26272 9820 26580 9829
rect 26272 9818 26278 9820
rect 26334 9818 26358 9820
rect 26414 9818 26438 9820
rect 26494 9818 26518 9820
rect 26574 9818 26580 9820
rect 26334 9766 26336 9818
rect 26516 9766 26518 9818
rect 26272 9764 26278 9766
rect 26334 9764 26358 9766
rect 26414 9764 26438 9766
rect 26494 9764 26518 9766
rect 26574 9764 26580 9766
rect 26272 9755 26580 9764
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 23768 6798 23796 7278
rect 24044 6798 24072 7278
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 24964 6730 24992 8434
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 25056 7478 25084 8366
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 25056 6730 25084 7414
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23584 6390 23612 6598
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24688 5710 24716 6054
rect 25608 5710 25636 7142
rect 25884 6662 25912 8570
rect 25976 7546 26004 9522
rect 27264 9450 27292 12786
rect 27356 12434 27384 13806
rect 27540 12918 27568 14214
rect 27528 12912 27580 12918
rect 27528 12854 27580 12860
rect 27632 12782 27660 14214
rect 27724 13938 27752 16050
rect 27816 15502 27844 16204
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 28092 15450 28120 20198
rect 28184 19446 28212 22596
rect 28540 22578 28592 22584
rect 29748 22574 29776 22918
rect 29736 22568 29788 22574
rect 29736 22510 29788 22516
rect 30102 22536 30158 22545
rect 30102 22471 30104 22480
rect 30156 22471 30158 22480
rect 30104 22442 30156 22448
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28460 21962 28488 22170
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 28460 21622 28488 21898
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 29748 21554 29776 21830
rect 30104 21684 30156 21690
rect 30208 21672 30236 32166
rect 30493 32124 30801 32133
rect 30493 32122 30499 32124
rect 30555 32122 30579 32124
rect 30635 32122 30659 32124
rect 30715 32122 30739 32124
rect 30795 32122 30801 32124
rect 30555 32070 30557 32122
rect 30737 32070 30739 32122
rect 30493 32068 30499 32070
rect 30555 32068 30579 32070
rect 30635 32068 30659 32070
rect 30715 32068 30739 32070
rect 30795 32068 30801 32070
rect 30493 32059 30801 32068
rect 30493 31036 30801 31045
rect 30493 31034 30499 31036
rect 30555 31034 30579 31036
rect 30635 31034 30659 31036
rect 30715 31034 30739 31036
rect 30795 31034 30801 31036
rect 30555 30982 30557 31034
rect 30737 30982 30739 31034
rect 30493 30980 30499 30982
rect 30555 30980 30579 30982
rect 30635 30980 30659 30982
rect 30715 30980 30739 30982
rect 30795 30980 30801 30982
rect 30493 30971 30801 30980
rect 30493 29948 30801 29957
rect 30493 29946 30499 29948
rect 30555 29946 30579 29948
rect 30635 29946 30659 29948
rect 30715 29946 30739 29948
rect 30795 29946 30801 29948
rect 30555 29894 30557 29946
rect 30737 29894 30739 29946
rect 30493 29892 30499 29894
rect 30555 29892 30579 29894
rect 30635 29892 30659 29894
rect 30715 29892 30739 29894
rect 30795 29892 30801 29894
rect 30493 29883 30801 29892
rect 30493 28860 30801 28869
rect 30493 28858 30499 28860
rect 30555 28858 30579 28860
rect 30635 28858 30659 28860
rect 30715 28858 30739 28860
rect 30795 28858 30801 28860
rect 30555 28806 30557 28858
rect 30737 28806 30739 28858
rect 30493 28804 30499 28806
rect 30555 28804 30579 28806
rect 30635 28804 30659 28806
rect 30715 28804 30739 28806
rect 30795 28804 30801 28806
rect 30493 28795 30801 28804
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 30493 27772 30801 27781
rect 30493 27770 30499 27772
rect 30555 27770 30579 27772
rect 30635 27770 30659 27772
rect 30715 27770 30739 27772
rect 30795 27770 30801 27772
rect 30555 27718 30557 27770
rect 30737 27718 30739 27770
rect 30493 27716 30499 27718
rect 30555 27716 30579 27718
rect 30635 27716 30659 27718
rect 30715 27716 30739 27718
rect 30795 27716 30801 27718
rect 30493 27707 30801 27716
rect 31128 27130 31156 28086
rect 32680 28076 32732 28082
rect 32680 28018 32732 28024
rect 32220 27396 32272 27402
rect 32220 27338 32272 27344
rect 31208 27328 31260 27334
rect 31208 27270 31260 27276
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 30493 26684 30801 26693
rect 30493 26682 30499 26684
rect 30555 26682 30579 26684
rect 30635 26682 30659 26684
rect 30715 26682 30739 26684
rect 30795 26682 30801 26684
rect 30555 26630 30557 26682
rect 30737 26630 30739 26682
rect 30493 26628 30499 26630
rect 30555 26628 30579 26630
rect 30635 26628 30659 26630
rect 30715 26628 30739 26630
rect 30795 26628 30801 26630
rect 30493 26619 30801 26628
rect 31220 26314 31248 27270
rect 32232 26586 32260 27338
rect 32220 26580 32272 26586
rect 32220 26522 32272 26528
rect 32692 26382 32720 28018
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 32680 26376 32732 26382
rect 32680 26318 32732 26324
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 31484 25968 31536 25974
rect 31484 25910 31536 25916
rect 30493 25596 30801 25605
rect 30493 25594 30499 25596
rect 30555 25594 30579 25596
rect 30635 25594 30659 25596
rect 30715 25594 30739 25596
rect 30795 25594 30801 25596
rect 30555 25542 30557 25594
rect 30737 25542 30739 25594
rect 30493 25540 30499 25542
rect 30555 25540 30579 25542
rect 30635 25540 30659 25542
rect 30715 25540 30739 25542
rect 30795 25540 30801 25542
rect 30493 25531 30801 25540
rect 31496 25294 31524 25910
rect 31944 25900 31996 25906
rect 31944 25842 31996 25848
rect 31484 25288 31536 25294
rect 31484 25230 31536 25236
rect 30380 25220 30432 25226
rect 30380 25162 30432 25168
rect 30392 24410 30420 25162
rect 31392 25152 31444 25158
rect 31392 25094 31444 25100
rect 30493 24508 30801 24517
rect 30493 24506 30499 24508
rect 30555 24506 30579 24508
rect 30635 24506 30659 24508
rect 30715 24506 30739 24508
rect 30795 24506 30801 24508
rect 30555 24454 30557 24506
rect 30737 24454 30739 24506
rect 30493 24452 30499 24454
rect 30555 24452 30579 24454
rect 30635 24452 30659 24454
rect 30715 24452 30739 24454
rect 30795 24452 30801 24454
rect 30493 24443 30801 24452
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 30493 23420 30801 23429
rect 30493 23418 30499 23420
rect 30555 23418 30579 23420
rect 30635 23418 30659 23420
rect 30715 23418 30739 23420
rect 30795 23418 30801 23420
rect 30555 23366 30557 23418
rect 30737 23366 30739 23418
rect 30493 23364 30499 23366
rect 30555 23364 30579 23366
rect 30635 23364 30659 23366
rect 30715 23364 30739 23366
rect 30795 23364 30801 23366
rect 30493 23355 30801 23364
rect 30380 22432 30432 22438
rect 30380 22374 30432 22380
rect 30392 22166 30420 22374
rect 30493 22332 30801 22341
rect 30493 22330 30499 22332
rect 30555 22330 30579 22332
rect 30635 22330 30659 22332
rect 30715 22330 30739 22332
rect 30795 22330 30801 22332
rect 30555 22278 30557 22330
rect 30737 22278 30739 22330
rect 30493 22276 30499 22278
rect 30555 22276 30579 22278
rect 30635 22276 30659 22278
rect 30715 22276 30739 22278
rect 30795 22276 30801 22278
rect 30493 22267 30801 22276
rect 30380 22160 30432 22166
rect 30380 22102 30432 22108
rect 30288 21956 30340 21962
rect 30288 21898 30340 21904
rect 30300 21690 30328 21898
rect 30156 21644 30236 21672
rect 30288 21684 30340 21690
rect 30104 21626 30156 21632
rect 30288 21626 30340 21632
rect 30392 21554 30420 22102
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 30380 21548 30432 21554
rect 30380 21490 30432 21496
rect 30104 21412 30156 21418
rect 30104 21354 30156 21360
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28460 21049 28488 21286
rect 28446 21040 28502 21049
rect 28446 20975 28502 20984
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28552 18766 28580 19246
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 28368 18290 28396 18566
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28552 18154 28580 18702
rect 28540 18148 28592 18154
rect 28540 18090 28592 18096
rect 28644 18034 28672 18702
rect 29012 18222 29040 19314
rect 29092 18420 29144 18426
rect 29092 18362 29144 18368
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 28552 18006 28672 18034
rect 28552 17678 28580 18006
rect 29012 17882 29040 18158
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28552 17202 28580 17614
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17338 28856 17478
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28920 17202 28948 17614
rect 29104 17338 29132 18362
rect 29196 18290 29224 19450
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29288 18766 29316 19246
rect 29276 18760 29328 18766
rect 29276 18702 29328 18708
rect 29380 18698 29408 19314
rect 30116 18766 30144 21354
rect 30493 21244 30801 21253
rect 30493 21242 30499 21244
rect 30555 21242 30579 21244
rect 30635 21242 30659 21244
rect 30715 21242 30739 21244
rect 30795 21242 30801 21244
rect 30555 21190 30557 21242
rect 30737 21190 30739 21242
rect 30493 21188 30499 21190
rect 30555 21188 30579 21190
rect 30635 21188 30659 21190
rect 30715 21188 30739 21190
rect 30795 21188 30801 21190
rect 30493 21179 30801 21188
rect 30944 21146 30972 24142
rect 31404 24070 31432 25094
rect 31496 24954 31524 25230
rect 31484 24948 31536 24954
rect 31484 24890 31536 24896
rect 31392 24064 31444 24070
rect 31392 24006 31444 24012
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 31036 22642 31064 23122
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31116 22568 31168 22574
rect 31300 22568 31352 22574
rect 31116 22510 31168 22516
rect 31298 22536 31300 22545
rect 31352 22536 31354 22545
rect 31024 22024 31076 22030
rect 31024 21966 31076 21972
rect 31036 21622 31064 21966
rect 31024 21616 31076 21622
rect 31024 21558 31076 21564
rect 31128 21554 31156 22510
rect 31298 22471 31354 22480
rect 31404 22030 31432 22578
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31404 21622 31432 21966
rect 31392 21616 31444 21622
rect 31392 21558 31444 21564
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 31128 21010 31156 21490
rect 31116 21004 31168 21010
rect 31116 20946 31168 20952
rect 31588 20602 31616 21966
rect 31772 21690 31800 23054
rect 31864 22778 31892 23258
rect 31852 22772 31904 22778
rect 31852 22714 31904 22720
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31956 21146 31984 25842
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 32324 24818 32352 25638
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32416 24274 32444 26318
rect 32692 26234 32720 26318
rect 32692 26206 32812 26234
rect 32784 25906 32812 26206
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32404 24268 32456 24274
rect 32404 24210 32456 24216
rect 32784 24206 32812 25842
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 33152 23322 33180 32166
rect 34713 31580 35021 31589
rect 34713 31578 34719 31580
rect 34775 31578 34799 31580
rect 34855 31578 34879 31580
rect 34935 31578 34959 31580
rect 35015 31578 35021 31580
rect 34775 31526 34777 31578
rect 34957 31526 34959 31578
rect 34713 31524 34719 31526
rect 34775 31524 34799 31526
rect 34855 31524 34879 31526
rect 34935 31524 34959 31526
rect 35015 31524 35021 31526
rect 34713 31515 35021 31524
rect 34713 30492 35021 30501
rect 34713 30490 34719 30492
rect 34775 30490 34799 30492
rect 34855 30490 34879 30492
rect 34935 30490 34959 30492
rect 35015 30490 35021 30492
rect 34775 30438 34777 30490
rect 34957 30438 34959 30490
rect 34713 30436 34719 30438
rect 34775 30436 34799 30438
rect 34855 30436 34879 30438
rect 34935 30436 34959 30438
rect 35015 30436 35021 30438
rect 34713 30427 35021 30436
rect 34713 29404 35021 29413
rect 34713 29402 34719 29404
rect 34775 29402 34799 29404
rect 34855 29402 34879 29404
rect 34935 29402 34959 29404
rect 35015 29402 35021 29404
rect 34775 29350 34777 29402
rect 34957 29350 34959 29402
rect 34713 29348 34719 29350
rect 34775 29348 34799 29350
rect 34855 29348 34879 29350
rect 34935 29348 34959 29350
rect 35015 29348 35021 29350
rect 34713 29339 35021 29348
rect 34713 28316 35021 28325
rect 34713 28314 34719 28316
rect 34775 28314 34799 28316
rect 34855 28314 34879 28316
rect 34935 28314 34959 28316
rect 35015 28314 35021 28316
rect 34775 28262 34777 28314
rect 34957 28262 34959 28314
rect 34713 28260 34719 28262
rect 34775 28260 34799 28262
rect 34855 28260 34879 28262
rect 34935 28260 34959 28262
rect 35015 28260 35021 28262
rect 34713 28251 35021 28260
rect 34713 27228 35021 27237
rect 34713 27226 34719 27228
rect 34775 27226 34799 27228
rect 34855 27226 34879 27228
rect 34935 27226 34959 27228
rect 35015 27226 35021 27228
rect 34775 27174 34777 27226
rect 34957 27174 34959 27226
rect 34713 27172 34719 27174
rect 34775 27172 34799 27174
rect 34855 27172 34879 27174
rect 34935 27172 34959 27174
rect 35015 27172 35021 27174
rect 34713 27163 35021 27172
rect 34713 26140 35021 26149
rect 34713 26138 34719 26140
rect 34775 26138 34799 26140
rect 34855 26138 34879 26140
rect 34935 26138 34959 26140
rect 35015 26138 35021 26140
rect 34775 26086 34777 26138
rect 34957 26086 34959 26138
rect 34713 26084 34719 26086
rect 34775 26084 34799 26086
rect 34855 26084 34879 26086
rect 34935 26084 34959 26086
rect 35015 26084 35021 26086
rect 34713 26075 35021 26084
rect 34713 25052 35021 25061
rect 34713 25050 34719 25052
rect 34775 25050 34799 25052
rect 34855 25050 34879 25052
rect 34935 25050 34959 25052
rect 35015 25050 35021 25052
rect 34775 24998 34777 25050
rect 34957 24998 34959 25050
rect 34713 24996 34719 24998
rect 34775 24996 34799 24998
rect 34855 24996 34879 24998
rect 34935 24996 34959 24998
rect 35015 24996 35021 24998
rect 34713 24987 35021 24996
rect 34713 23964 35021 23973
rect 34713 23962 34719 23964
rect 34775 23962 34799 23964
rect 34855 23962 34879 23964
rect 34935 23962 34959 23964
rect 35015 23962 35021 23964
rect 34775 23910 34777 23962
rect 34957 23910 34959 23962
rect 34713 23908 34719 23910
rect 34775 23908 34799 23910
rect 34855 23908 34879 23910
rect 34935 23908 34959 23910
rect 35015 23908 35021 23910
rect 34713 23899 35021 23908
rect 33140 23316 33192 23322
rect 33140 23258 33192 23264
rect 32680 23180 32732 23186
rect 32680 23122 32732 23128
rect 33140 23180 33192 23186
rect 33140 23122 33192 23128
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32048 22778 32076 23054
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32416 22574 32444 23054
rect 32692 22642 32720 23122
rect 33152 22710 33180 23122
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32404 22568 32456 22574
rect 32404 22510 32456 22516
rect 32416 22030 32444 22510
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 32220 21412 32272 21418
rect 32220 21354 32272 21360
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 32232 20942 32260 21354
rect 32416 21146 32444 21966
rect 32600 21554 32628 21966
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32496 20936 32548 20942
rect 32496 20878 32548 20884
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 31944 20392 31996 20398
rect 31944 20334 31996 20340
rect 30493 20156 30801 20165
rect 30493 20154 30499 20156
rect 30555 20154 30579 20156
rect 30635 20154 30659 20156
rect 30715 20154 30739 20156
rect 30795 20154 30801 20156
rect 30555 20102 30557 20154
rect 30737 20102 30739 20154
rect 30493 20100 30499 20102
rect 30555 20100 30579 20102
rect 30635 20100 30659 20102
rect 30715 20100 30739 20102
rect 30795 20100 30801 20102
rect 30493 20091 30801 20100
rect 31956 19854 31984 20334
rect 32232 19854 32260 20878
rect 32404 20460 32456 20466
rect 32404 20402 32456 20408
rect 32312 20324 32364 20330
rect 32312 20266 32364 20272
rect 32324 19990 32352 20266
rect 32312 19984 32364 19990
rect 32312 19926 32364 19932
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 31956 19446 31984 19790
rect 32232 19514 32260 19790
rect 32416 19718 32444 20402
rect 32508 19922 32536 20878
rect 32600 20602 32628 21490
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32496 19916 32548 19922
rect 32496 19858 32548 19864
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32220 19508 32272 19514
rect 32220 19450 32272 19456
rect 31944 19440 31996 19446
rect 31944 19382 31996 19388
rect 32416 19378 32444 19654
rect 32508 19530 32536 19858
rect 32508 19514 32628 19530
rect 32508 19508 32640 19514
rect 32508 19502 32588 19508
rect 32588 19450 32640 19456
rect 31392 19372 31444 19378
rect 31392 19314 31444 19320
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 30493 19068 30801 19077
rect 30493 19066 30499 19068
rect 30555 19066 30579 19068
rect 30635 19066 30659 19068
rect 30715 19066 30739 19068
rect 30795 19066 30801 19068
rect 30555 19014 30557 19066
rect 30737 19014 30739 19066
rect 30493 19012 30499 19014
rect 30555 19012 30579 19014
rect 30635 19012 30659 19014
rect 30715 19012 30739 19014
rect 30795 19012 30801 19014
rect 30493 19003 30801 19012
rect 29828 18760 29880 18766
rect 29748 18720 29828 18748
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29748 18290 29776 18720
rect 29828 18702 29880 18708
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 28540 17196 28592 17202
rect 28540 17138 28592 17144
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29012 16114 29040 16594
rect 29104 16522 29132 17274
rect 29748 16658 29776 18226
rect 30116 18222 30144 18702
rect 31404 18358 31432 19314
rect 32416 18834 32444 19314
rect 32404 18828 32456 18834
rect 32404 18770 32456 18776
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 31392 18352 31444 18358
rect 31392 18294 31444 18300
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30493 17980 30801 17989
rect 30493 17978 30499 17980
rect 30555 17978 30579 17980
rect 30635 17978 30659 17980
rect 30715 17978 30739 17980
rect 30795 17978 30801 17980
rect 30555 17926 30557 17978
rect 30737 17926 30739 17978
rect 30493 17924 30499 17926
rect 30555 17924 30579 17926
rect 30635 17924 30659 17926
rect 30715 17924 30739 17926
rect 30795 17924 30801 17926
rect 30493 17915 30801 17924
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 30944 17338 30972 17614
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 29092 16516 29144 16522
rect 29092 16458 29144 16464
rect 29104 16250 29132 16458
rect 30300 16454 30328 17070
rect 30493 16892 30801 16901
rect 30493 16890 30499 16892
rect 30555 16890 30579 16892
rect 30635 16890 30659 16892
rect 30715 16890 30739 16892
rect 30795 16890 30801 16892
rect 30555 16838 30557 16890
rect 30737 16838 30739 16890
rect 30493 16836 30499 16838
rect 30555 16836 30579 16838
rect 30635 16836 30659 16838
rect 30715 16836 30739 16838
rect 30795 16836 30801 16838
rect 30493 16827 30801 16836
rect 31128 16794 31156 17546
rect 31404 17202 31432 18294
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31312 16794 31340 16934
rect 31116 16788 31168 16794
rect 31116 16730 31168 16736
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30288 16448 30340 16454
rect 31312 16402 31340 16730
rect 31404 16658 31432 17138
rect 31588 16726 31616 17138
rect 31576 16720 31628 16726
rect 31576 16662 31628 16668
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 30288 16390 30340 16396
rect 29092 16244 29144 16250
rect 29092 16186 29144 16192
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15570 28212 15846
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28448 15496 28500 15502
rect 27816 13977 27844 15438
rect 28092 15422 28212 15450
rect 28448 15438 28500 15444
rect 27802 13968 27858 13977
rect 27712 13932 27764 13938
rect 27802 13903 27804 13912
rect 27712 13874 27764 13880
rect 27856 13903 27858 13912
rect 27804 13874 27856 13880
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27356 12406 27476 12434
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 27356 10742 27384 10950
rect 27344 10736 27396 10742
rect 27344 10678 27396 10684
rect 27252 9444 27304 9450
rect 27252 9386 27304 9392
rect 27448 9178 27476 12406
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 27724 10690 27752 11018
rect 27632 10674 27752 10690
rect 27632 10668 27764 10674
rect 27632 10662 27712 10668
rect 27632 10198 27660 10662
rect 27712 10610 27764 10616
rect 27712 10532 27764 10538
rect 27712 10474 27764 10480
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 27724 9722 27752 10474
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27816 9586 27844 12174
rect 28000 11354 28028 12786
rect 28080 12708 28132 12714
rect 28080 12650 28132 12656
rect 28092 11762 28120 12650
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27988 11348 28040 11354
rect 27988 11290 28040 11296
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 26272 8732 26580 8741
rect 26272 8730 26278 8732
rect 26334 8730 26358 8732
rect 26414 8730 26438 8732
rect 26494 8730 26518 8732
rect 26574 8730 26580 8732
rect 26334 8678 26336 8730
rect 26516 8678 26518 8730
rect 26272 8676 26278 8678
rect 26334 8676 26358 8678
rect 26414 8676 26438 8678
rect 26494 8676 26518 8678
rect 26574 8676 26580 8678
rect 26272 8667 26580 8676
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 25976 5914 26004 7482
rect 26068 7410 26096 8434
rect 26272 7644 26580 7653
rect 26272 7642 26278 7644
rect 26334 7642 26358 7644
rect 26414 7642 26438 7644
rect 26494 7642 26518 7644
rect 26574 7642 26580 7644
rect 26334 7590 26336 7642
rect 26516 7590 26518 7642
rect 26272 7588 26278 7590
rect 26334 7588 26358 7590
rect 26414 7588 26438 7590
rect 26494 7588 26518 7590
rect 26574 7588 26580 7590
rect 26272 7579 26580 7588
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 27908 6662 27936 10610
rect 28092 8294 28120 11698
rect 28184 10810 28212 15422
rect 28460 12986 28488 15438
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28264 12912 28316 12918
rect 28264 12854 28316 12860
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 28092 8090 28120 8230
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 26272 6556 26580 6565
rect 26272 6554 26278 6556
rect 26334 6554 26358 6556
rect 26414 6554 26438 6556
rect 26494 6554 26518 6556
rect 26574 6554 26580 6556
rect 26334 6502 26336 6554
rect 26516 6502 26518 6554
rect 26272 6500 26278 6502
rect 26334 6500 26358 6502
rect 26414 6500 26438 6502
rect 26494 6500 26518 6502
rect 26574 6500 26580 6502
rect 26272 6491 26580 6500
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 24688 5370 24716 5646
rect 27908 5642 27936 6598
rect 27896 5636 27948 5642
rect 27896 5578 27948 5584
rect 26272 5468 26580 5477
rect 26272 5466 26278 5468
rect 26334 5466 26358 5468
rect 26414 5466 26438 5468
rect 26494 5466 26518 5468
rect 26574 5466 26580 5468
rect 26334 5414 26336 5466
rect 26516 5414 26518 5466
rect 26272 5412 26278 5414
rect 26334 5412 26358 5414
rect 26414 5412 26438 5414
rect 26494 5412 26518 5414
rect 26574 5412 26580 5414
rect 26272 5403 26580 5412
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25044 5092 25096 5098
rect 25044 5034 25096 5040
rect 22052 4924 22360 4933
rect 22052 4922 22058 4924
rect 22114 4922 22138 4924
rect 22194 4922 22218 4924
rect 22274 4922 22298 4924
rect 22354 4922 22360 4924
rect 22114 4870 22116 4922
rect 22296 4870 22298 4922
rect 22052 4868 22058 4870
rect 22114 4868 22138 4870
rect 22194 4868 22218 4870
rect 22274 4868 22298 4870
rect 22354 4868 22360 4870
rect 22052 4859 22360 4868
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 17420 4146 17448 4558
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 17512 4146 17540 4422
rect 17831 4380 18139 4389
rect 17831 4378 17837 4380
rect 17893 4378 17917 4380
rect 17973 4378 17997 4380
rect 18053 4378 18077 4380
rect 18133 4378 18139 4380
rect 17893 4326 17895 4378
rect 18075 4326 18077 4378
rect 17831 4324 17837 4326
rect 17893 4324 17917 4326
rect 17973 4324 17997 4326
rect 18053 4324 18077 4326
rect 18133 4324 18139 4326
rect 17831 4315 18139 4324
rect 18248 4162 18276 4422
rect 17972 4146 18276 4162
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17960 4140 18276 4146
rect 18012 4134 18276 4140
rect 17960 4082 18012 4088
rect 19076 3942 19104 4422
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 17831 3292 18139 3301
rect 17831 3290 17837 3292
rect 17893 3290 17917 3292
rect 17973 3290 17997 3292
rect 18053 3290 18077 3292
rect 18133 3290 18139 3292
rect 17893 3238 17895 3290
rect 18075 3238 18077 3290
rect 17831 3236 17837 3238
rect 17893 3236 17917 3238
rect 17973 3236 17997 3238
rect 18053 3236 18077 3238
rect 18133 3236 18139 3238
rect 17831 3227 18139 3236
rect 18248 3194 18276 3334
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18248 2514 18276 3130
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 19076 2446 19104 3878
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 3194 19472 3470
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19720 3058 19748 4082
rect 19812 3466 19840 4422
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 20456 2990 20484 4626
rect 20732 3058 20760 4694
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 20824 3738 20852 4422
rect 20916 4146 20944 4558
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 21560 4146 21588 4422
rect 22112 4146 22140 4422
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20824 2446 20852 3674
rect 21100 3126 21128 3878
rect 21192 3194 21220 4082
rect 22296 4026 22324 4082
rect 22296 3998 22416 4026
rect 22052 3836 22360 3845
rect 22052 3834 22058 3836
rect 22114 3834 22138 3836
rect 22194 3834 22218 3836
rect 22274 3834 22298 3836
rect 22354 3834 22360 3836
rect 22114 3782 22116 3834
rect 22296 3782 22298 3834
rect 22052 3780 22058 3782
rect 22114 3780 22138 3782
rect 22194 3780 22218 3782
rect 22274 3780 22298 3782
rect 22354 3780 22360 3782
rect 22052 3771 22360 3780
rect 22388 3738 22416 3998
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22480 3534 22508 4218
rect 24596 4146 24624 4422
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21088 3120 21140 3126
rect 21088 3062 21140 3068
rect 21100 2446 21128 3062
rect 22756 3058 22784 3538
rect 23400 3534 23428 3878
rect 24688 3754 24716 4694
rect 25056 4690 25084 5034
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24596 3738 24716 3754
rect 24584 3732 24716 3738
rect 24636 3726 24716 3732
rect 24584 3674 24636 3680
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22052 2748 22360 2757
rect 22052 2746 22058 2748
rect 22114 2746 22138 2748
rect 22194 2746 22218 2748
rect 22274 2746 22298 2748
rect 22354 2746 22360 2748
rect 22114 2694 22116 2746
rect 22296 2694 22298 2746
rect 22052 2692 22058 2694
rect 22114 2692 22138 2694
rect 22194 2692 22218 2694
rect 22274 2692 22298 2694
rect 22354 2692 22360 2694
rect 22052 2683 22360 2692
rect 23400 2446 23428 3470
rect 24688 2774 24716 3726
rect 25700 3534 25728 4966
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25792 3466 25820 5170
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 25884 4214 25912 4558
rect 26148 4548 26200 4554
rect 26148 4490 26200 4496
rect 26160 4282 26188 4490
rect 26272 4380 26580 4389
rect 26272 4378 26278 4380
rect 26334 4378 26358 4380
rect 26414 4378 26438 4380
rect 26494 4378 26518 4380
rect 26574 4378 26580 4380
rect 26334 4326 26336 4378
rect 26516 4326 26518 4378
rect 26272 4324 26278 4326
rect 26334 4324 26358 4326
rect 26414 4324 26438 4326
rect 26494 4324 26518 4326
rect 26574 4324 26580 4326
rect 26272 4315 26580 4324
rect 26148 4276 26200 4282
rect 26148 4218 26200 4224
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25884 3534 25912 4150
rect 26620 4146 26648 5102
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25056 2774 25084 2926
rect 25792 2854 25820 3402
rect 26160 2990 26188 3538
rect 26620 3534 26648 3878
rect 26804 3670 26832 4422
rect 28092 4214 28120 7754
rect 28276 6730 28304 12854
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 28368 11830 28396 12582
rect 28552 12238 28580 12922
rect 28644 12238 28672 13806
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 28632 12232 28684 12238
rect 28632 12174 28684 12180
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 28368 10674 28396 11290
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28368 7818 28396 10610
rect 28460 10606 28488 12106
rect 28552 11626 28580 12174
rect 28736 11898 28764 13942
rect 28828 12374 28856 14350
rect 29012 14346 29040 16050
rect 30116 16046 30144 16390
rect 30300 16114 30328 16390
rect 30944 16374 31340 16402
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 30104 16040 30156 16046
rect 30104 15982 30156 15988
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29472 15570 29500 15846
rect 30493 15804 30801 15813
rect 30493 15802 30499 15804
rect 30555 15802 30579 15804
rect 30635 15802 30659 15804
rect 30715 15802 30739 15804
rect 30795 15802 30801 15804
rect 30555 15750 30557 15802
rect 30737 15750 30739 15802
rect 30493 15748 30499 15750
rect 30555 15748 30579 15750
rect 30635 15748 30659 15750
rect 30715 15748 30739 15750
rect 30795 15748 30801 15750
rect 30493 15739 30801 15748
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29920 15020 29972 15026
rect 29920 14962 29972 14968
rect 29644 14884 29696 14890
rect 29644 14826 29696 14832
rect 29000 14340 29052 14346
rect 29000 14282 29052 14288
rect 29012 14074 29040 14282
rect 29000 14068 29052 14074
rect 29000 14010 29052 14016
rect 28908 14000 28960 14006
rect 28906 13968 28908 13977
rect 28960 13968 28962 13977
rect 29656 13938 29684 14826
rect 29932 14074 29960 14962
rect 30493 14716 30801 14725
rect 30493 14714 30499 14716
rect 30555 14714 30579 14716
rect 30635 14714 30659 14716
rect 30715 14714 30739 14716
rect 30795 14714 30801 14716
rect 30555 14662 30557 14714
rect 30737 14662 30739 14714
rect 30493 14660 30499 14662
rect 30555 14660 30579 14662
rect 30635 14660 30659 14662
rect 30715 14660 30739 14662
rect 30795 14660 30801 14662
rect 30493 14651 30801 14660
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 30116 14074 30144 14350
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 28906 13903 28962 13912
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 29656 13734 29684 13874
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 29644 13728 29696 13734
rect 29644 13670 29696 13676
rect 28920 12714 28948 13670
rect 29656 12850 29684 13670
rect 30288 12912 30340 12918
rect 30392 12866 30420 13874
rect 30493 13628 30801 13637
rect 30493 13626 30499 13628
rect 30555 13626 30579 13628
rect 30635 13626 30659 13628
rect 30715 13626 30739 13628
rect 30795 13626 30801 13628
rect 30555 13574 30557 13626
rect 30737 13574 30739 13626
rect 30493 13572 30499 13574
rect 30555 13572 30579 13574
rect 30635 13572 30659 13574
rect 30715 13572 30739 13574
rect 30795 13572 30801 13574
rect 30493 13563 30801 13572
rect 30340 12860 30420 12866
rect 30288 12854 30420 12860
rect 29644 12844 29696 12850
rect 30300 12838 30420 12854
rect 29644 12786 29696 12792
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 28908 12708 28960 12714
rect 28908 12650 28960 12656
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 30208 11762 30236 12718
rect 30392 11830 30420 12838
rect 30493 12540 30801 12549
rect 30493 12538 30499 12540
rect 30555 12538 30579 12540
rect 30635 12538 30659 12540
rect 30715 12538 30739 12540
rect 30795 12538 30801 12540
rect 30555 12486 30557 12538
rect 30737 12486 30739 12538
rect 30493 12484 30499 12486
rect 30555 12484 30579 12486
rect 30635 12484 30659 12486
rect 30715 12484 30739 12486
rect 30795 12484 30801 12486
rect 30493 12475 30801 12484
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28724 11552 28776 11558
rect 28724 11494 28776 11500
rect 28736 10810 28764 11494
rect 30208 11150 30236 11698
rect 29368 11144 29420 11150
rect 29368 11086 29420 11092
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28448 10600 28500 10606
rect 28448 10542 28500 10548
rect 28736 10130 28764 10746
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 28920 10130 28948 10610
rect 28724 10124 28776 10130
rect 28724 10066 28776 10072
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 29012 9874 29040 9930
rect 28920 9846 29040 9874
rect 28920 9586 28948 9846
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 29380 9518 29408 11086
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29748 10062 29776 10950
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 29932 10062 29960 10610
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 29920 10056 29972 10062
rect 29920 9998 29972 10004
rect 30208 9586 30236 11086
rect 30288 10056 30340 10062
rect 30288 9998 30340 10004
rect 30196 9580 30248 9586
rect 30196 9522 30248 9528
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28828 8974 28856 9318
rect 28816 8968 28868 8974
rect 29092 8968 29144 8974
rect 28816 8910 28868 8916
rect 28920 8916 29092 8922
rect 28920 8910 29144 8916
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28264 6724 28316 6730
rect 28264 6666 28316 6672
rect 28276 6458 28304 6666
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28828 6186 28856 8910
rect 28920 8894 29132 8910
rect 28920 8838 28948 8894
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28920 6798 28948 8570
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 28816 6180 28868 6186
rect 28816 6122 28868 6128
rect 29012 5846 29040 8774
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29104 7546 29132 8502
rect 29092 7540 29144 7546
rect 29092 7482 29144 7488
rect 29104 6798 29132 7482
rect 29092 6792 29144 6798
rect 29092 6734 29144 6740
rect 29196 6390 29224 8774
rect 29380 7478 29408 9454
rect 30208 8974 30236 9522
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29748 8498 29776 8774
rect 30208 8498 30236 8910
rect 30300 8906 30328 9998
rect 30392 9110 30420 11766
rect 30493 11452 30801 11461
rect 30493 11450 30499 11452
rect 30555 11450 30579 11452
rect 30635 11450 30659 11452
rect 30715 11450 30739 11452
rect 30795 11450 30801 11452
rect 30555 11398 30557 11450
rect 30737 11398 30739 11450
rect 30493 11396 30499 11398
rect 30555 11396 30579 11398
rect 30635 11396 30659 11398
rect 30715 11396 30739 11398
rect 30795 11396 30801 11398
rect 30493 11387 30801 11396
rect 30852 10742 30880 11834
rect 30944 11218 30972 16374
rect 31404 16182 31432 16594
rect 32048 16590 32076 18702
rect 32416 18290 32444 18770
rect 32496 18420 32548 18426
rect 32496 18362 32548 18368
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32312 18216 32364 18222
rect 32312 18158 32364 18164
rect 32324 17746 32352 18158
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32220 17332 32272 17338
rect 32220 17274 32272 17280
rect 32232 16794 32260 17274
rect 32416 17202 32444 18226
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32036 16584 32088 16590
rect 32036 16526 32088 16532
rect 31392 16176 31444 16182
rect 31392 16118 31444 16124
rect 32312 16040 32364 16046
rect 32312 15982 32364 15988
rect 32220 15972 32272 15978
rect 32220 15914 32272 15920
rect 31760 15700 31812 15706
rect 31760 15642 31812 15648
rect 31772 14482 31800 15642
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 31944 14272 31996 14278
rect 31944 14214 31996 14220
rect 31956 14074 31984 14214
rect 31944 14068 31996 14074
rect 31944 14010 31996 14016
rect 32036 14068 32088 14074
rect 32036 14010 32088 14016
rect 32048 13870 32076 14010
rect 32036 13864 32088 13870
rect 32036 13806 32088 13812
rect 32140 12986 32168 14350
rect 32128 12980 32180 12986
rect 32128 12922 32180 12928
rect 31024 12708 31076 12714
rect 31024 12650 31076 12656
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 30840 10736 30892 10742
rect 30840 10678 30892 10684
rect 31036 10470 31064 12650
rect 32128 12368 32180 12374
rect 32128 12310 32180 12316
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 11898 31248 12038
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31220 11354 31248 11834
rect 32140 11762 32168 12310
rect 32232 11898 32260 15914
rect 32324 15706 32352 15982
rect 32312 15700 32364 15706
rect 32312 15642 32364 15648
rect 32312 14476 32364 14482
rect 32312 14418 32364 14424
rect 32324 13870 32352 14418
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32324 13530 32352 13806
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32508 12850 32536 18362
rect 32600 16658 32628 19450
rect 32692 19242 32720 22578
rect 33152 22098 33180 22646
rect 33336 22574 33364 23054
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33520 22710 33548 22918
rect 34713 22876 35021 22885
rect 34713 22874 34719 22876
rect 34775 22874 34799 22876
rect 34855 22874 34879 22876
rect 34935 22874 34959 22876
rect 35015 22874 35021 22876
rect 34775 22822 34777 22874
rect 34957 22822 34959 22874
rect 34713 22820 34719 22822
rect 34775 22820 34799 22822
rect 34855 22820 34879 22822
rect 34935 22820 34959 22822
rect 35015 22820 35021 22822
rect 34713 22811 35021 22820
rect 33508 22704 33560 22710
rect 33508 22646 33560 22652
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33140 22092 33192 22098
rect 33140 22034 33192 22040
rect 33336 22030 33364 22510
rect 33704 22234 33732 22578
rect 33692 22228 33744 22234
rect 33692 22170 33744 22176
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32956 20936 33008 20942
rect 32956 20878 33008 20884
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 32772 20868 32824 20874
rect 32772 20810 32824 20816
rect 32784 20466 32812 20810
rect 32772 20460 32824 20466
rect 32772 20402 32824 20408
rect 32680 19236 32732 19242
rect 32680 19178 32732 19184
rect 32784 18902 32812 20402
rect 32968 20330 32996 20878
rect 33060 20466 33088 20878
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 32956 20324 33008 20330
rect 32956 20266 33008 20272
rect 33060 19514 33088 20402
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 33336 18970 33364 21966
rect 34713 21788 35021 21797
rect 34713 21786 34719 21788
rect 34775 21786 34799 21788
rect 34855 21786 34879 21788
rect 34935 21786 34959 21788
rect 35015 21786 35021 21788
rect 34775 21734 34777 21786
rect 34957 21734 34959 21786
rect 34713 21732 34719 21734
rect 34775 21732 34799 21734
rect 34855 21732 34879 21734
rect 34935 21732 34959 21734
rect 35015 21732 35021 21734
rect 34713 21723 35021 21732
rect 34713 20700 35021 20709
rect 34713 20698 34719 20700
rect 34775 20698 34799 20700
rect 34855 20698 34879 20700
rect 34935 20698 34959 20700
rect 35015 20698 35021 20700
rect 34775 20646 34777 20698
rect 34957 20646 34959 20698
rect 34713 20644 34719 20646
rect 34775 20644 34799 20646
rect 34855 20644 34879 20646
rect 34935 20644 34959 20646
rect 35015 20644 35021 20646
rect 34713 20635 35021 20644
rect 34713 19612 35021 19621
rect 34713 19610 34719 19612
rect 34775 19610 34799 19612
rect 34855 19610 34879 19612
rect 34935 19610 34959 19612
rect 35015 19610 35021 19612
rect 34775 19558 34777 19610
rect 34957 19558 34959 19610
rect 34713 19556 34719 19558
rect 34775 19556 34799 19558
rect 34855 19556 34879 19558
rect 34935 19556 34959 19558
rect 35015 19556 35021 19558
rect 34713 19547 35021 19556
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 32772 18896 32824 18902
rect 32692 18844 32772 18850
rect 32692 18838 32824 18844
rect 32692 18822 32812 18838
rect 32692 18426 32720 18822
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32680 18420 32732 18426
rect 32680 18362 32732 18368
rect 32784 17678 32812 18702
rect 34713 18524 35021 18533
rect 34713 18522 34719 18524
rect 34775 18522 34799 18524
rect 34855 18522 34879 18524
rect 34935 18522 34959 18524
rect 35015 18522 35021 18524
rect 34775 18470 34777 18522
rect 34957 18470 34959 18522
rect 34713 18468 34719 18470
rect 34775 18468 34799 18470
rect 34855 18468 34879 18470
rect 34935 18468 34959 18470
rect 35015 18468 35021 18470
rect 34713 18459 35021 18468
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 32772 17672 32824 17678
rect 32772 17614 32824 17620
rect 32876 17338 32904 18158
rect 34348 17921 34376 18158
rect 34334 17912 34390 17921
rect 34334 17847 34390 17856
rect 33232 17536 33284 17542
rect 33232 17478 33284 17484
rect 33244 17338 33272 17478
rect 34713 17436 35021 17445
rect 34713 17434 34719 17436
rect 34775 17434 34799 17436
rect 34855 17434 34879 17436
rect 34935 17434 34959 17436
rect 35015 17434 35021 17436
rect 34775 17382 34777 17434
rect 34957 17382 34959 17434
rect 34713 17380 34719 17382
rect 34775 17380 34799 17382
rect 34855 17380 34879 17382
rect 34935 17380 34959 17382
rect 35015 17380 35021 17382
rect 34713 17371 35021 17380
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33232 17332 33284 17338
rect 33232 17274 33284 17280
rect 32772 17196 32824 17202
rect 32772 17138 32824 17144
rect 32784 16998 32812 17138
rect 32772 16992 32824 16998
rect 32772 16934 32824 16940
rect 32588 16652 32640 16658
rect 32588 16594 32640 16600
rect 32600 16250 32628 16594
rect 32588 16244 32640 16250
rect 32588 16186 32640 16192
rect 32784 14278 32812 16934
rect 33692 16720 33744 16726
rect 33692 16662 33744 16668
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 33060 15366 33088 16186
rect 33232 16176 33284 16182
rect 33232 16118 33284 16124
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 33244 14618 33272 16118
rect 33704 15502 33732 16662
rect 34713 16348 35021 16357
rect 34713 16346 34719 16348
rect 34775 16346 34799 16348
rect 34855 16346 34879 16348
rect 34935 16346 34959 16348
rect 35015 16346 35021 16348
rect 34775 16294 34777 16346
rect 34957 16294 34959 16346
rect 34713 16292 34719 16294
rect 34775 16292 34799 16294
rect 34855 16292 34879 16294
rect 34935 16292 34959 16294
rect 35015 16292 35021 16294
rect 34713 16283 35021 16292
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33888 15706 33916 16050
rect 33876 15700 33928 15706
rect 33876 15642 33928 15648
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33232 14612 33284 14618
rect 33232 14554 33284 14560
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32784 13870 32812 14214
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 33244 12986 33272 14554
rect 33428 13734 33456 15438
rect 33600 15428 33652 15434
rect 33600 15370 33652 15376
rect 33612 15162 33640 15370
rect 34713 15260 35021 15269
rect 34713 15258 34719 15260
rect 34775 15258 34799 15260
rect 34855 15258 34879 15260
rect 34935 15258 34959 15260
rect 35015 15258 35021 15260
rect 34775 15206 34777 15258
rect 34957 15206 34959 15258
rect 34713 15204 34719 15206
rect 34775 15204 34799 15206
rect 34855 15204 34879 15206
rect 34935 15204 34959 15206
rect 35015 15204 35021 15206
rect 34713 15195 35021 15204
rect 33600 15156 33652 15162
rect 33600 15098 33652 15104
rect 33416 13728 33468 13734
rect 33416 13670 33468 13676
rect 33232 12980 33284 12986
rect 33232 12922 33284 12928
rect 33428 12850 33456 13670
rect 33612 13326 33640 15098
rect 34713 14172 35021 14181
rect 34713 14170 34719 14172
rect 34775 14170 34799 14172
rect 34855 14170 34879 14172
rect 34935 14170 34959 14172
rect 35015 14170 35021 14172
rect 34775 14118 34777 14170
rect 34957 14118 34959 14170
rect 34713 14116 34719 14118
rect 34775 14116 34799 14118
rect 34855 14116 34879 14118
rect 34935 14116 34959 14118
rect 35015 14116 35021 14118
rect 34713 14107 35021 14116
rect 33692 14068 33744 14074
rect 33692 14010 33744 14016
rect 33600 13320 33652 13326
rect 33600 13262 33652 13268
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 33416 12844 33468 12850
rect 33416 12786 33468 12792
rect 32220 11892 32272 11898
rect 32220 11834 32272 11840
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 31576 11552 31628 11558
rect 31576 11494 31628 11500
rect 31208 11348 31260 11354
rect 31208 11290 31260 11296
rect 31588 11082 31616 11494
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 30493 10364 30801 10373
rect 30493 10362 30499 10364
rect 30555 10362 30579 10364
rect 30635 10362 30659 10364
rect 30715 10362 30739 10364
rect 30795 10362 30801 10364
rect 30555 10310 30557 10362
rect 30737 10310 30739 10362
rect 30493 10308 30499 10310
rect 30555 10308 30579 10310
rect 30635 10308 30659 10310
rect 30715 10308 30739 10310
rect 30795 10308 30801 10310
rect 30493 10299 30801 10308
rect 31392 9648 31444 9654
rect 31392 9590 31444 9596
rect 30493 9276 30801 9285
rect 30493 9274 30499 9276
rect 30555 9274 30579 9276
rect 30635 9274 30659 9276
rect 30715 9274 30739 9276
rect 30795 9274 30801 9276
rect 30555 9222 30557 9274
rect 30737 9222 30739 9274
rect 30493 9220 30499 9222
rect 30555 9220 30579 9222
rect 30635 9220 30659 9222
rect 30715 9220 30739 9222
rect 30795 9220 30801 9222
rect 30493 9211 30801 9220
rect 30380 9104 30432 9110
rect 30380 9046 30432 9052
rect 30288 8900 30340 8906
rect 30288 8842 30340 8848
rect 30300 8634 30328 8842
rect 31404 8634 31432 9590
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31772 8566 31800 9318
rect 31760 8560 31812 8566
rect 31760 8502 31812 8508
rect 32140 8498 32168 11698
rect 33416 11688 33468 11694
rect 33416 11630 33468 11636
rect 32312 11552 32364 11558
rect 32312 11494 32364 11500
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32232 10606 32260 11086
rect 32324 10742 32352 11494
rect 32312 10736 32364 10742
rect 32312 10678 32364 10684
rect 32220 10600 32272 10606
rect 32220 10542 32272 10548
rect 32232 10266 32260 10542
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32220 10260 32272 10266
rect 32220 10202 32272 10208
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 32232 9178 32260 9862
rect 32324 9654 32352 10406
rect 33428 10062 33456 11630
rect 33612 10810 33640 11834
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33704 10062 33732 14010
rect 34713 13084 35021 13093
rect 34713 13082 34719 13084
rect 34775 13082 34799 13084
rect 34855 13082 34879 13084
rect 34935 13082 34959 13084
rect 35015 13082 35021 13084
rect 34775 13030 34777 13082
rect 34957 13030 34959 13082
rect 34713 13028 34719 13030
rect 34775 13028 34799 13030
rect 34855 13028 34879 13030
rect 34935 13028 34959 13030
rect 35015 13028 35021 13030
rect 34713 13019 35021 13028
rect 34713 11996 35021 12005
rect 34713 11994 34719 11996
rect 34775 11994 34799 11996
rect 34855 11994 34879 11996
rect 34935 11994 34959 11996
rect 35015 11994 35021 11996
rect 34775 11942 34777 11994
rect 34957 11942 34959 11994
rect 34713 11940 34719 11942
rect 34775 11940 34799 11942
rect 34855 11940 34879 11942
rect 34935 11940 34959 11942
rect 35015 11940 35021 11942
rect 34713 11931 35021 11940
rect 34713 10908 35021 10917
rect 34713 10906 34719 10908
rect 34775 10906 34799 10908
rect 34855 10906 34879 10908
rect 34935 10906 34959 10908
rect 35015 10906 35021 10908
rect 34775 10854 34777 10906
rect 34957 10854 34959 10906
rect 34713 10852 34719 10854
rect 34775 10852 34799 10854
rect 34855 10852 34879 10854
rect 34935 10852 34959 10854
rect 35015 10852 35021 10854
rect 34713 10843 35021 10852
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33692 10056 33744 10062
rect 33692 9998 33744 10004
rect 33692 9920 33744 9926
rect 33692 9862 33744 9868
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 32312 9648 32364 9654
rect 32312 9590 32364 9596
rect 33704 9382 33732 9862
rect 33692 9376 33744 9382
rect 33692 9318 33744 9324
rect 32220 9172 32272 9178
rect 32220 9114 32272 9120
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32324 8498 32352 8910
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 30493 8188 30801 8197
rect 30493 8186 30499 8188
rect 30555 8186 30579 8188
rect 30635 8186 30659 8188
rect 30715 8186 30739 8188
rect 30795 8186 30801 8188
rect 30555 8134 30557 8186
rect 30737 8134 30739 8186
rect 30493 8132 30499 8134
rect 30555 8132 30579 8134
rect 30635 8132 30659 8134
rect 30715 8132 30739 8134
rect 30795 8132 30801 8134
rect 30493 8123 30801 8132
rect 30380 7744 30432 7750
rect 30380 7686 30432 7692
rect 29368 7472 29420 7478
rect 29368 7414 29420 7420
rect 29276 6724 29328 6730
rect 29276 6666 29328 6672
rect 29184 6384 29236 6390
rect 29184 6326 29236 6332
rect 29288 5914 29316 6666
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 29380 5710 29408 7414
rect 30392 7410 30420 7686
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29840 6254 29868 6734
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 27068 4140 27120 4146
rect 27068 4082 27120 4088
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 26792 3664 26844 3670
rect 26792 3606 26844 3612
rect 27080 3618 27108 4082
rect 27816 3738 27844 4082
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 27620 3664 27672 3670
rect 26608 3528 26660 3534
rect 26608 3470 26660 3476
rect 26272 3292 26580 3301
rect 26272 3290 26278 3292
rect 26334 3290 26358 3292
rect 26414 3290 26438 3292
rect 26494 3290 26518 3292
rect 26574 3290 26580 3292
rect 26334 3238 26336 3290
rect 26516 3238 26518 3290
rect 26272 3236 26278 3238
rect 26334 3236 26358 3238
rect 26414 3236 26438 3238
rect 26494 3236 26518 3238
rect 26574 3236 26580 3238
rect 26272 3227 26580 3236
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26620 2854 26648 3470
rect 26804 3058 26832 3606
rect 27080 3602 27200 3618
rect 27620 3606 27672 3612
rect 27080 3596 27212 3602
rect 27080 3590 27160 3596
rect 27160 3538 27212 3544
rect 27632 3058 27660 3606
rect 28368 3534 28396 3878
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 26792 3052 26844 3058
rect 26792 2994 26844 3000
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 24688 2746 25084 2774
rect 25056 2446 25084 2746
rect 26252 2446 26280 2790
rect 27632 2446 27660 2994
rect 28368 2446 28396 3470
rect 29840 3194 29868 6190
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 30392 3126 30420 7346
rect 30493 7100 30801 7109
rect 30493 7098 30499 7100
rect 30555 7098 30579 7100
rect 30635 7098 30659 7100
rect 30715 7098 30739 7100
rect 30795 7098 30801 7100
rect 30555 7046 30557 7098
rect 30737 7046 30739 7098
rect 30493 7044 30499 7046
rect 30555 7044 30579 7046
rect 30635 7044 30659 7046
rect 30715 7044 30739 7046
rect 30795 7044 30801 7046
rect 30493 7035 30801 7044
rect 30852 6458 30880 8434
rect 32324 8090 32352 8434
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 33704 7886 33732 9318
rect 33888 8906 33916 9862
rect 34713 9820 35021 9829
rect 34713 9818 34719 9820
rect 34775 9818 34799 9820
rect 34855 9818 34879 9820
rect 34935 9818 34959 9820
rect 35015 9818 35021 9820
rect 34775 9766 34777 9818
rect 34957 9766 34959 9818
rect 34713 9764 34719 9766
rect 34775 9764 34799 9766
rect 34855 9764 34879 9766
rect 34935 9764 34959 9766
rect 35015 9764 35021 9766
rect 34713 9755 35021 9764
rect 33876 8900 33928 8906
rect 33876 8842 33928 8848
rect 34713 8732 35021 8741
rect 34713 8730 34719 8732
rect 34775 8730 34799 8732
rect 34855 8730 34879 8732
rect 34935 8730 34959 8732
rect 35015 8730 35021 8732
rect 34775 8678 34777 8730
rect 34957 8678 34959 8730
rect 34713 8676 34719 8678
rect 34775 8676 34799 8678
rect 34855 8676 34879 8678
rect 34935 8676 34959 8678
rect 35015 8676 35021 8678
rect 34713 8667 35021 8676
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 34713 7644 35021 7653
rect 34713 7642 34719 7644
rect 34775 7642 34799 7644
rect 34855 7642 34879 7644
rect 34935 7642 34959 7644
rect 35015 7642 35021 7644
rect 34775 7590 34777 7642
rect 34957 7590 34959 7642
rect 34713 7588 34719 7590
rect 34775 7588 34799 7590
rect 34855 7588 34879 7590
rect 34935 7588 34959 7590
rect 35015 7588 35021 7590
rect 34713 7579 35021 7588
rect 34713 6556 35021 6565
rect 34713 6554 34719 6556
rect 34775 6554 34799 6556
rect 34855 6554 34879 6556
rect 34935 6554 34959 6556
rect 35015 6554 35021 6556
rect 34775 6502 34777 6554
rect 34957 6502 34959 6554
rect 34713 6500 34719 6502
rect 34775 6500 34799 6502
rect 34855 6500 34879 6502
rect 34935 6500 34959 6502
rect 35015 6500 35021 6502
rect 34713 6491 35021 6500
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30493 6012 30801 6021
rect 30493 6010 30499 6012
rect 30555 6010 30579 6012
rect 30635 6010 30659 6012
rect 30715 6010 30739 6012
rect 30795 6010 30801 6012
rect 30555 5958 30557 6010
rect 30737 5958 30739 6010
rect 30493 5956 30499 5958
rect 30555 5956 30579 5958
rect 30635 5956 30659 5958
rect 30715 5956 30739 5958
rect 30795 5956 30801 5958
rect 30493 5947 30801 5956
rect 34713 5468 35021 5477
rect 34713 5466 34719 5468
rect 34775 5466 34799 5468
rect 34855 5466 34879 5468
rect 34935 5466 34959 5468
rect 35015 5466 35021 5468
rect 34775 5414 34777 5466
rect 34957 5414 34959 5466
rect 34713 5412 34719 5414
rect 34775 5412 34799 5414
rect 34855 5412 34879 5414
rect 34935 5412 34959 5414
rect 35015 5412 35021 5414
rect 34713 5403 35021 5412
rect 30493 4924 30801 4933
rect 30493 4922 30499 4924
rect 30555 4922 30579 4924
rect 30635 4922 30659 4924
rect 30715 4922 30739 4924
rect 30795 4922 30801 4924
rect 30555 4870 30557 4922
rect 30737 4870 30739 4922
rect 30493 4868 30499 4870
rect 30555 4868 30579 4870
rect 30635 4868 30659 4870
rect 30715 4868 30739 4870
rect 30795 4868 30801 4870
rect 30493 4859 30801 4868
rect 34713 4380 35021 4389
rect 34713 4378 34719 4380
rect 34775 4378 34799 4380
rect 34855 4378 34879 4380
rect 34935 4378 34959 4380
rect 35015 4378 35021 4380
rect 34775 4326 34777 4378
rect 34957 4326 34959 4378
rect 34713 4324 34719 4326
rect 34775 4324 34799 4326
rect 34855 4324 34879 4326
rect 34935 4324 34959 4326
rect 35015 4324 35021 4326
rect 34713 4315 35021 4324
rect 30493 3836 30801 3845
rect 30493 3834 30499 3836
rect 30555 3834 30579 3836
rect 30635 3834 30659 3836
rect 30715 3834 30739 3836
rect 30795 3834 30801 3836
rect 30555 3782 30557 3834
rect 30737 3782 30739 3834
rect 30493 3780 30499 3782
rect 30555 3780 30579 3782
rect 30635 3780 30659 3782
rect 30715 3780 30739 3782
rect 30795 3780 30801 3782
rect 30493 3771 30801 3780
rect 34713 3292 35021 3301
rect 34713 3290 34719 3292
rect 34775 3290 34799 3292
rect 34855 3290 34879 3292
rect 34935 3290 34959 3292
rect 35015 3290 35021 3292
rect 34775 3238 34777 3290
rect 34957 3238 34959 3290
rect 34713 3236 34719 3238
rect 34775 3236 34799 3238
rect 34855 3236 34879 3238
rect 34935 3236 34959 3238
rect 35015 3236 35021 3238
rect 34713 3227 35021 3236
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 30493 2748 30801 2757
rect 30493 2746 30499 2748
rect 30555 2746 30579 2748
rect 30635 2746 30659 2748
rect 30715 2746 30739 2748
rect 30795 2746 30801 2748
rect 30555 2694 30557 2746
rect 30737 2694 30739 2746
rect 30493 2692 30499 2694
rect 30555 2692 30579 2694
rect 30635 2692 30659 2694
rect 30715 2692 30739 2694
rect 30795 2692 30801 2694
rect 30493 2683 30801 2692
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7760 1306 7788 2382
rect 7668 1278 7788 1306
rect 7668 800 7696 1278
rect 8956 800 8984 2382
rect 9390 2204 9698 2213
rect 9390 2202 9396 2204
rect 9452 2202 9476 2204
rect 9532 2202 9556 2204
rect 9612 2202 9636 2204
rect 9692 2202 9698 2204
rect 9452 2150 9454 2202
rect 9634 2150 9636 2202
rect 9390 2148 9396 2150
rect 9452 2148 9476 2150
rect 9532 2148 9556 2150
rect 9612 2148 9636 2150
rect 9692 2148 9698 2150
rect 9390 2139 9698 2148
rect 10244 800 10272 2382
rect 11532 800 11560 2382
rect 12820 800 12848 2382
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 19248 2372 19300 2378
rect 19248 2314 19300 2320
rect 20536 2372 20588 2378
rect 20536 2314 20588 2320
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 24400 2372 24452 2378
rect 24400 2314 24452 2320
rect 25688 2372 25740 2378
rect 25688 2314 25740 2320
rect 26976 2372 27028 2378
rect 26976 2314 27028 2320
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 14108 800 14136 2314
rect 15396 800 15424 2314
rect 16684 800 16712 2314
rect 17831 2204 18139 2213
rect 17831 2202 17837 2204
rect 17893 2202 17917 2204
rect 17973 2202 17997 2204
rect 18053 2202 18077 2204
rect 18133 2202 18139 2204
rect 17893 2150 17895 2202
rect 18075 2150 18077 2202
rect 17831 2148 17837 2150
rect 17893 2148 17917 2150
rect 17973 2148 17997 2150
rect 18053 2148 18077 2150
rect 18133 2148 18139 2150
rect 17831 2139 18139 2148
rect 17972 870 18092 898
rect 17972 800 18000 870
rect 1214 0 1270 800
rect 2502 0 2558 800
rect 3790 0 3846 800
rect 5078 0 5134 800
rect 6366 0 6422 800
rect 7654 0 7710 800
rect 8942 0 8998 800
rect 10230 0 10286 800
rect 11518 0 11574 800
rect 12806 0 12862 800
rect 14094 0 14150 800
rect 15382 0 15438 800
rect 16670 0 16726 800
rect 17958 0 18014 800
rect 18064 762 18092 870
rect 18248 762 18276 2314
rect 19260 800 19288 2314
rect 20548 800 20576 2314
rect 21836 800 21864 2314
rect 23124 800 23152 2314
rect 24412 800 24440 2314
rect 25700 800 25728 2314
rect 26272 2204 26580 2213
rect 26272 2202 26278 2204
rect 26334 2202 26358 2204
rect 26414 2202 26438 2204
rect 26494 2202 26518 2204
rect 26574 2202 26580 2204
rect 26334 2150 26336 2202
rect 26516 2150 26518 2202
rect 26272 2148 26278 2150
rect 26334 2148 26358 2150
rect 26414 2148 26438 2150
rect 26494 2148 26518 2150
rect 26574 2148 26580 2150
rect 26272 2139 26580 2148
rect 26988 800 27016 2314
rect 28276 800 28304 2314
rect 29564 800 29592 2382
rect 30852 800 30880 2382
rect 32140 800 32168 2382
rect 33428 800 33456 2382
rect 34612 2304 34664 2310
rect 34612 2246 34664 2252
rect 34624 1170 34652 2246
rect 34713 2204 35021 2213
rect 34713 2202 34719 2204
rect 34775 2202 34799 2204
rect 34855 2202 34879 2204
rect 34935 2202 34959 2204
rect 35015 2202 35021 2204
rect 34775 2150 34777 2202
rect 34957 2150 34959 2202
rect 34713 2148 34719 2150
rect 34775 2148 34799 2150
rect 34855 2148 34879 2150
rect 34935 2148 34959 2150
rect 35015 2148 35021 2150
rect 34713 2139 35021 2148
rect 34624 1142 34744 1170
rect 34716 800 34744 1142
rect 18064 734 18276 762
rect 19246 0 19302 800
rect 20534 0 20590 800
rect 21822 0 21878 800
rect 23110 0 23166 800
rect 24398 0 24454 800
rect 25686 0 25742 800
rect 26974 0 27030 800
rect 28262 0 28318 800
rect 29550 0 29606 800
rect 30838 0 30894 800
rect 32126 0 32182 800
rect 33414 0 33470 800
rect 34702 0 34758 800
<< via2 >>
rect 9396 33754 9452 33756
rect 9476 33754 9532 33756
rect 9556 33754 9612 33756
rect 9636 33754 9692 33756
rect 9396 33702 9442 33754
rect 9442 33702 9452 33754
rect 9476 33702 9506 33754
rect 9506 33702 9518 33754
rect 9518 33702 9532 33754
rect 9556 33702 9570 33754
rect 9570 33702 9582 33754
rect 9582 33702 9612 33754
rect 9636 33702 9646 33754
rect 9646 33702 9692 33754
rect 9396 33700 9452 33702
rect 9476 33700 9532 33702
rect 9556 33700 9612 33702
rect 9636 33700 9692 33702
rect 17837 33754 17893 33756
rect 17917 33754 17973 33756
rect 17997 33754 18053 33756
rect 18077 33754 18133 33756
rect 17837 33702 17883 33754
rect 17883 33702 17893 33754
rect 17917 33702 17947 33754
rect 17947 33702 17959 33754
rect 17959 33702 17973 33754
rect 17997 33702 18011 33754
rect 18011 33702 18023 33754
rect 18023 33702 18053 33754
rect 18077 33702 18087 33754
rect 18087 33702 18133 33754
rect 17837 33700 17893 33702
rect 17917 33700 17973 33702
rect 17997 33700 18053 33702
rect 18077 33700 18133 33702
rect 26278 33754 26334 33756
rect 26358 33754 26414 33756
rect 26438 33754 26494 33756
rect 26518 33754 26574 33756
rect 26278 33702 26324 33754
rect 26324 33702 26334 33754
rect 26358 33702 26388 33754
rect 26388 33702 26400 33754
rect 26400 33702 26414 33754
rect 26438 33702 26452 33754
rect 26452 33702 26464 33754
rect 26464 33702 26494 33754
rect 26518 33702 26528 33754
rect 26528 33702 26574 33754
rect 26278 33700 26334 33702
rect 26358 33700 26414 33702
rect 26438 33700 26494 33702
rect 26518 33700 26574 33702
rect 34719 33754 34775 33756
rect 34799 33754 34855 33756
rect 34879 33754 34935 33756
rect 34959 33754 35015 33756
rect 34719 33702 34765 33754
rect 34765 33702 34775 33754
rect 34799 33702 34829 33754
rect 34829 33702 34841 33754
rect 34841 33702 34855 33754
rect 34879 33702 34893 33754
rect 34893 33702 34905 33754
rect 34905 33702 34935 33754
rect 34959 33702 34969 33754
rect 34969 33702 35015 33754
rect 34719 33700 34775 33702
rect 34799 33700 34855 33702
rect 34879 33700 34935 33702
rect 34959 33700 35015 33702
rect 5176 33210 5232 33212
rect 5256 33210 5312 33212
rect 5336 33210 5392 33212
rect 5416 33210 5472 33212
rect 5176 33158 5222 33210
rect 5222 33158 5232 33210
rect 5256 33158 5286 33210
rect 5286 33158 5298 33210
rect 5298 33158 5312 33210
rect 5336 33158 5350 33210
rect 5350 33158 5362 33210
rect 5362 33158 5392 33210
rect 5416 33158 5426 33210
rect 5426 33158 5472 33210
rect 5176 33156 5232 33158
rect 5256 33156 5312 33158
rect 5336 33156 5392 33158
rect 5416 33156 5472 33158
rect 5176 32122 5232 32124
rect 5256 32122 5312 32124
rect 5336 32122 5392 32124
rect 5416 32122 5472 32124
rect 5176 32070 5222 32122
rect 5222 32070 5232 32122
rect 5256 32070 5286 32122
rect 5286 32070 5298 32122
rect 5298 32070 5312 32122
rect 5336 32070 5350 32122
rect 5350 32070 5362 32122
rect 5362 32070 5392 32122
rect 5416 32070 5426 32122
rect 5426 32070 5472 32122
rect 5176 32068 5232 32070
rect 5256 32068 5312 32070
rect 5336 32068 5392 32070
rect 5416 32068 5472 32070
rect 3698 19796 3700 19816
rect 3700 19796 3752 19816
rect 3752 19796 3754 19816
rect 3698 19760 3754 19796
rect 4158 19896 4214 19952
rect 9396 32666 9452 32668
rect 9476 32666 9532 32668
rect 9556 32666 9612 32668
rect 9636 32666 9692 32668
rect 9396 32614 9442 32666
rect 9442 32614 9452 32666
rect 9476 32614 9506 32666
rect 9506 32614 9518 32666
rect 9518 32614 9532 32666
rect 9556 32614 9570 32666
rect 9570 32614 9582 32666
rect 9582 32614 9612 32666
rect 9636 32614 9646 32666
rect 9646 32614 9692 32666
rect 9396 32612 9452 32614
rect 9476 32612 9532 32614
rect 9556 32612 9612 32614
rect 9636 32612 9692 32614
rect 5176 31034 5232 31036
rect 5256 31034 5312 31036
rect 5336 31034 5392 31036
rect 5416 31034 5472 31036
rect 5176 30982 5222 31034
rect 5222 30982 5232 31034
rect 5256 30982 5286 31034
rect 5286 30982 5298 31034
rect 5298 30982 5312 31034
rect 5336 30982 5350 31034
rect 5350 30982 5362 31034
rect 5362 30982 5392 31034
rect 5416 30982 5426 31034
rect 5426 30982 5472 31034
rect 5176 30980 5232 30982
rect 5256 30980 5312 30982
rect 5336 30980 5392 30982
rect 5416 30980 5472 30982
rect 5176 29946 5232 29948
rect 5256 29946 5312 29948
rect 5336 29946 5392 29948
rect 5416 29946 5472 29948
rect 5176 29894 5222 29946
rect 5222 29894 5232 29946
rect 5256 29894 5286 29946
rect 5286 29894 5298 29946
rect 5298 29894 5312 29946
rect 5336 29894 5350 29946
rect 5350 29894 5362 29946
rect 5362 29894 5392 29946
rect 5416 29894 5426 29946
rect 5426 29894 5472 29946
rect 5176 29892 5232 29894
rect 5256 29892 5312 29894
rect 5336 29892 5392 29894
rect 5416 29892 5472 29894
rect 5176 28858 5232 28860
rect 5256 28858 5312 28860
rect 5336 28858 5392 28860
rect 5416 28858 5472 28860
rect 5176 28806 5222 28858
rect 5222 28806 5232 28858
rect 5256 28806 5286 28858
rect 5286 28806 5298 28858
rect 5298 28806 5312 28858
rect 5336 28806 5350 28858
rect 5350 28806 5362 28858
rect 5362 28806 5392 28858
rect 5416 28806 5426 28858
rect 5426 28806 5472 28858
rect 5176 28804 5232 28806
rect 5256 28804 5312 28806
rect 5336 28804 5392 28806
rect 5416 28804 5472 28806
rect 9396 31578 9452 31580
rect 9476 31578 9532 31580
rect 9556 31578 9612 31580
rect 9636 31578 9692 31580
rect 9396 31526 9442 31578
rect 9442 31526 9452 31578
rect 9476 31526 9506 31578
rect 9506 31526 9518 31578
rect 9518 31526 9532 31578
rect 9556 31526 9570 31578
rect 9570 31526 9582 31578
rect 9582 31526 9612 31578
rect 9636 31526 9646 31578
rect 9646 31526 9692 31578
rect 9396 31524 9452 31526
rect 9476 31524 9532 31526
rect 9556 31524 9612 31526
rect 9636 31524 9692 31526
rect 13617 33210 13673 33212
rect 13697 33210 13753 33212
rect 13777 33210 13833 33212
rect 13857 33210 13913 33212
rect 13617 33158 13663 33210
rect 13663 33158 13673 33210
rect 13697 33158 13727 33210
rect 13727 33158 13739 33210
rect 13739 33158 13753 33210
rect 13777 33158 13791 33210
rect 13791 33158 13803 33210
rect 13803 33158 13833 33210
rect 13857 33158 13867 33210
rect 13867 33158 13913 33210
rect 13617 33156 13673 33158
rect 13697 33156 13753 33158
rect 13777 33156 13833 33158
rect 13857 33156 13913 33158
rect 9396 30490 9452 30492
rect 9476 30490 9532 30492
rect 9556 30490 9612 30492
rect 9636 30490 9692 30492
rect 9396 30438 9442 30490
rect 9442 30438 9452 30490
rect 9476 30438 9506 30490
rect 9506 30438 9518 30490
rect 9518 30438 9532 30490
rect 9556 30438 9570 30490
rect 9570 30438 9582 30490
rect 9582 30438 9612 30490
rect 9636 30438 9646 30490
rect 9646 30438 9692 30490
rect 9396 30436 9452 30438
rect 9476 30436 9532 30438
rect 9556 30436 9612 30438
rect 9636 30436 9692 30438
rect 9396 29402 9452 29404
rect 9476 29402 9532 29404
rect 9556 29402 9612 29404
rect 9636 29402 9692 29404
rect 9396 29350 9442 29402
rect 9442 29350 9452 29402
rect 9476 29350 9506 29402
rect 9506 29350 9518 29402
rect 9518 29350 9532 29402
rect 9556 29350 9570 29402
rect 9570 29350 9582 29402
rect 9582 29350 9612 29402
rect 9636 29350 9646 29402
rect 9646 29350 9692 29402
rect 9396 29348 9452 29350
rect 9476 29348 9532 29350
rect 9556 29348 9612 29350
rect 9636 29348 9692 29350
rect 9396 28314 9452 28316
rect 9476 28314 9532 28316
rect 9556 28314 9612 28316
rect 9636 28314 9692 28316
rect 9396 28262 9442 28314
rect 9442 28262 9452 28314
rect 9476 28262 9506 28314
rect 9506 28262 9518 28314
rect 9518 28262 9532 28314
rect 9556 28262 9570 28314
rect 9570 28262 9582 28314
rect 9582 28262 9612 28314
rect 9636 28262 9646 28314
rect 9646 28262 9692 28314
rect 9396 28260 9452 28262
rect 9476 28260 9532 28262
rect 9556 28260 9612 28262
rect 9636 28260 9692 28262
rect 5176 27770 5232 27772
rect 5256 27770 5312 27772
rect 5336 27770 5392 27772
rect 5416 27770 5472 27772
rect 5176 27718 5222 27770
rect 5222 27718 5232 27770
rect 5256 27718 5286 27770
rect 5286 27718 5298 27770
rect 5298 27718 5312 27770
rect 5336 27718 5350 27770
rect 5350 27718 5362 27770
rect 5362 27718 5392 27770
rect 5416 27718 5426 27770
rect 5426 27718 5472 27770
rect 5176 27716 5232 27718
rect 5256 27716 5312 27718
rect 5336 27716 5392 27718
rect 5416 27716 5472 27718
rect 5176 26682 5232 26684
rect 5256 26682 5312 26684
rect 5336 26682 5392 26684
rect 5416 26682 5472 26684
rect 5176 26630 5222 26682
rect 5222 26630 5232 26682
rect 5256 26630 5286 26682
rect 5286 26630 5298 26682
rect 5298 26630 5312 26682
rect 5336 26630 5350 26682
rect 5350 26630 5362 26682
rect 5362 26630 5392 26682
rect 5416 26630 5426 26682
rect 5426 26630 5472 26682
rect 5176 26628 5232 26630
rect 5256 26628 5312 26630
rect 5336 26628 5392 26630
rect 5416 26628 5472 26630
rect 9396 27226 9452 27228
rect 9476 27226 9532 27228
rect 9556 27226 9612 27228
rect 9636 27226 9692 27228
rect 9396 27174 9442 27226
rect 9442 27174 9452 27226
rect 9476 27174 9506 27226
rect 9506 27174 9518 27226
rect 9518 27174 9532 27226
rect 9556 27174 9570 27226
rect 9570 27174 9582 27226
rect 9582 27174 9612 27226
rect 9636 27174 9646 27226
rect 9646 27174 9692 27226
rect 9396 27172 9452 27174
rect 9476 27172 9532 27174
rect 9556 27172 9612 27174
rect 9636 27172 9692 27174
rect 9396 26138 9452 26140
rect 9476 26138 9532 26140
rect 9556 26138 9612 26140
rect 9636 26138 9692 26140
rect 9396 26086 9442 26138
rect 9442 26086 9452 26138
rect 9476 26086 9506 26138
rect 9506 26086 9518 26138
rect 9518 26086 9532 26138
rect 9556 26086 9570 26138
rect 9570 26086 9582 26138
rect 9582 26086 9612 26138
rect 9636 26086 9646 26138
rect 9646 26086 9692 26138
rect 9396 26084 9452 26086
rect 9476 26084 9532 26086
rect 9556 26084 9612 26086
rect 9636 26084 9692 26086
rect 5176 25594 5232 25596
rect 5256 25594 5312 25596
rect 5336 25594 5392 25596
rect 5416 25594 5472 25596
rect 5176 25542 5222 25594
rect 5222 25542 5232 25594
rect 5256 25542 5286 25594
rect 5286 25542 5298 25594
rect 5298 25542 5312 25594
rect 5336 25542 5350 25594
rect 5350 25542 5362 25594
rect 5362 25542 5392 25594
rect 5416 25542 5426 25594
rect 5426 25542 5472 25594
rect 5176 25540 5232 25542
rect 5256 25540 5312 25542
rect 5336 25540 5392 25542
rect 5416 25540 5472 25542
rect 5176 24506 5232 24508
rect 5256 24506 5312 24508
rect 5336 24506 5392 24508
rect 5416 24506 5472 24508
rect 5176 24454 5222 24506
rect 5222 24454 5232 24506
rect 5256 24454 5286 24506
rect 5286 24454 5298 24506
rect 5298 24454 5312 24506
rect 5336 24454 5350 24506
rect 5350 24454 5362 24506
rect 5362 24454 5392 24506
rect 5416 24454 5426 24506
rect 5426 24454 5472 24506
rect 5176 24452 5232 24454
rect 5256 24452 5312 24454
rect 5336 24452 5392 24454
rect 5416 24452 5472 24454
rect 9396 25050 9452 25052
rect 9476 25050 9532 25052
rect 9556 25050 9612 25052
rect 9636 25050 9692 25052
rect 9396 24998 9442 25050
rect 9442 24998 9452 25050
rect 9476 24998 9506 25050
rect 9506 24998 9518 25050
rect 9518 24998 9532 25050
rect 9556 24998 9570 25050
rect 9570 24998 9582 25050
rect 9582 24998 9612 25050
rect 9636 24998 9646 25050
rect 9646 24998 9692 25050
rect 9396 24996 9452 24998
rect 9476 24996 9532 24998
rect 9556 24996 9612 24998
rect 9636 24996 9692 24998
rect 5176 23418 5232 23420
rect 5256 23418 5312 23420
rect 5336 23418 5392 23420
rect 5416 23418 5472 23420
rect 5176 23366 5222 23418
rect 5222 23366 5232 23418
rect 5256 23366 5286 23418
rect 5286 23366 5298 23418
rect 5298 23366 5312 23418
rect 5336 23366 5350 23418
rect 5350 23366 5362 23418
rect 5362 23366 5392 23418
rect 5416 23366 5426 23418
rect 5426 23366 5472 23418
rect 5176 23364 5232 23366
rect 5256 23364 5312 23366
rect 5336 23364 5392 23366
rect 5416 23364 5472 23366
rect 5176 22330 5232 22332
rect 5256 22330 5312 22332
rect 5336 22330 5392 22332
rect 5416 22330 5472 22332
rect 5176 22278 5222 22330
rect 5222 22278 5232 22330
rect 5256 22278 5286 22330
rect 5286 22278 5298 22330
rect 5298 22278 5312 22330
rect 5336 22278 5350 22330
rect 5350 22278 5362 22330
rect 5362 22278 5392 22330
rect 5416 22278 5426 22330
rect 5426 22278 5472 22330
rect 5176 22276 5232 22278
rect 5256 22276 5312 22278
rect 5336 22276 5392 22278
rect 5416 22276 5472 22278
rect 5176 21242 5232 21244
rect 5256 21242 5312 21244
rect 5336 21242 5392 21244
rect 5416 21242 5472 21244
rect 5176 21190 5222 21242
rect 5222 21190 5232 21242
rect 5256 21190 5286 21242
rect 5286 21190 5298 21242
rect 5298 21190 5312 21242
rect 5336 21190 5350 21242
rect 5350 21190 5362 21242
rect 5362 21190 5392 21242
rect 5416 21190 5426 21242
rect 5426 21190 5472 21242
rect 5176 21188 5232 21190
rect 5256 21188 5312 21190
rect 5336 21188 5392 21190
rect 5416 21188 5472 21190
rect 5176 20154 5232 20156
rect 5256 20154 5312 20156
rect 5336 20154 5392 20156
rect 5416 20154 5472 20156
rect 5176 20102 5222 20154
rect 5222 20102 5232 20154
rect 5256 20102 5286 20154
rect 5286 20102 5298 20154
rect 5298 20102 5312 20154
rect 5336 20102 5350 20154
rect 5350 20102 5362 20154
rect 5362 20102 5392 20154
rect 5416 20102 5426 20154
rect 5426 20102 5472 20154
rect 5176 20100 5232 20102
rect 5256 20100 5312 20102
rect 5336 20100 5392 20102
rect 5416 20100 5472 20102
rect 5354 19896 5410 19952
rect 4894 19760 4950 19816
rect 5176 19066 5232 19068
rect 5256 19066 5312 19068
rect 5336 19066 5392 19068
rect 5416 19066 5472 19068
rect 5176 19014 5222 19066
rect 5222 19014 5232 19066
rect 5256 19014 5286 19066
rect 5286 19014 5298 19066
rect 5298 19014 5312 19066
rect 5336 19014 5350 19066
rect 5350 19014 5362 19066
rect 5362 19014 5392 19066
rect 5416 19014 5426 19066
rect 5426 19014 5472 19066
rect 5176 19012 5232 19014
rect 5256 19012 5312 19014
rect 5336 19012 5392 19014
rect 5416 19012 5472 19014
rect 5176 17978 5232 17980
rect 5256 17978 5312 17980
rect 5336 17978 5392 17980
rect 5416 17978 5472 17980
rect 5176 17926 5222 17978
rect 5222 17926 5232 17978
rect 5256 17926 5286 17978
rect 5286 17926 5298 17978
rect 5298 17926 5312 17978
rect 5336 17926 5350 17978
rect 5350 17926 5362 17978
rect 5362 17926 5392 17978
rect 5416 17926 5426 17978
rect 5426 17926 5472 17978
rect 5176 17924 5232 17926
rect 5256 17924 5312 17926
rect 5336 17924 5392 17926
rect 5416 17924 5472 17926
rect 9396 23962 9452 23964
rect 9476 23962 9532 23964
rect 9556 23962 9612 23964
rect 9636 23962 9692 23964
rect 9396 23910 9442 23962
rect 9442 23910 9452 23962
rect 9476 23910 9506 23962
rect 9506 23910 9518 23962
rect 9518 23910 9532 23962
rect 9556 23910 9570 23962
rect 9570 23910 9582 23962
rect 9582 23910 9612 23962
rect 9636 23910 9646 23962
rect 9646 23910 9692 23962
rect 9396 23908 9452 23910
rect 9476 23908 9532 23910
rect 9556 23908 9612 23910
rect 9636 23908 9692 23910
rect 9396 22874 9452 22876
rect 9476 22874 9532 22876
rect 9556 22874 9612 22876
rect 9636 22874 9692 22876
rect 9396 22822 9442 22874
rect 9442 22822 9452 22874
rect 9476 22822 9506 22874
rect 9506 22822 9518 22874
rect 9518 22822 9532 22874
rect 9556 22822 9570 22874
rect 9570 22822 9582 22874
rect 9582 22822 9612 22874
rect 9636 22822 9646 22874
rect 9646 22822 9692 22874
rect 9396 22820 9452 22822
rect 9476 22820 9532 22822
rect 9556 22820 9612 22822
rect 9636 22820 9692 22822
rect 5176 16890 5232 16892
rect 5256 16890 5312 16892
rect 5336 16890 5392 16892
rect 5416 16890 5472 16892
rect 5176 16838 5222 16890
rect 5222 16838 5232 16890
rect 5256 16838 5286 16890
rect 5286 16838 5298 16890
rect 5298 16838 5312 16890
rect 5336 16838 5350 16890
rect 5350 16838 5362 16890
rect 5362 16838 5392 16890
rect 5416 16838 5426 16890
rect 5426 16838 5472 16890
rect 5176 16836 5232 16838
rect 5256 16836 5312 16838
rect 5336 16836 5392 16838
rect 5416 16836 5472 16838
rect 5176 15802 5232 15804
rect 5256 15802 5312 15804
rect 5336 15802 5392 15804
rect 5416 15802 5472 15804
rect 5176 15750 5222 15802
rect 5222 15750 5232 15802
rect 5256 15750 5286 15802
rect 5286 15750 5298 15802
rect 5298 15750 5312 15802
rect 5336 15750 5350 15802
rect 5350 15750 5362 15802
rect 5362 15750 5392 15802
rect 5416 15750 5426 15802
rect 5426 15750 5472 15802
rect 5176 15748 5232 15750
rect 5256 15748 5312 15750
rect 5336 15748 5392 15750
rect 5416 15748 5472 15750
rect 5176 14714 5232 14716
rect 5256 14714 5312 14716
rect 5336 14714 5392 14716
rect 5416 14714 5472 14716
rect 5176 14662 5222 14714
rect 5222 14662 5232 14714
rect 5256 14662 5286 14714
rect 5286 14662 5298 14714
rect 5298 14662 5312 14714
rect 5336 14662 5350 14714
rect 5350 14662 5362 14714
rect 5362 14662 5392 14714
rect 5416 14662 5426 14714
rect 5426 14662 5472 14714
rect 5176 14660 5232 14662
rect 5256 14660 5312 14662
rect 5336 14660 5392 14662
rect 5416 14660 5472 14662
rect 5176 13626 5232 13628
rect 5256 13626 5312 13628
rect 5336 13626 5392 13628
rect 5416 13626 5472 13628
rect 5176 13574 5222 13626
rect 5222 13574 5232 13626
rect 5256 13574 5286 13626
rect 5286 13574 5298 13626
rect 5298 13574 5312 13626
rect 5336 13574 5350 13626
rect 5350 13574 5362 13626
rect 5362 13574 5392 13626
rect 5416 13574 5426 13626
rect 5426 13574 5472 13626
rect 5176 13572 5232 13574
rect 5256 13572 5312 13574
rect 5336 13572 5392 13574
rect 5416 13572 5472 13574
rect 5176 12538 5232 12540
rect 5256 12538 5312 12540
rect 5336 12538 5392 12540
rect 5416 12538 5472 12540
rect 5176 12486 5222 12538
rect 5222 12486 5232 12538
rect 5256 12486 5286 12538
rect 5286 12486 5298 12538
rect 5298 12486 5312 12538
rect 5336 12486 5350 12538
rect 5350 12486 5362 12538
rect 5362 12486 5392 12538
rect 5416 12486 5426 12538
rect 5426 12486 5472 12538
rect 5176 12484 5232 12486
rect 5256 12484 5312 12486
rect 5336 12484 5392 12486
rect 5416 12484 5472 12486
rect 9396 21786 9452 21788
rect 9476 21786 9532 21788
rect 9556 21786 9612 21788
rect 9636 21786 9692 21788
rect 9396 21734 9442 21786
rect 9442 21734 9452 21786
rect 9476 21734 9506 21786
rect 9506 21734 9518 21786
rect 9518 21734 9532 21786
rect 9556 21734 9570 21786
rect 9570 21734 9582 21786
rect 9582 21734 9612 21786
rect 9636 21734 9646 21786
rect 9646 21734 9692 21786
rect 9396 21732 9452 21734
rect 9476 21732 9532 21734
rect 9556 21732 9612 21734
rect 9636 21732 9692 21734
rect 9396 20698 9452 20700
rect 9476 20698 9532 20700
rect 9556 20698 9612 20700
rect 9636 20698 9692 20700
rect 9396 20646 9442 20698
rect 9442 20646 9452 20698
rect 9476 20646 9506 20698
rect 9506 20646 9518 20698
rect 9518 20646 9532 20698
rect 9556 20646 9570 20698
rect 9570 20646 9582 20698
rect 9582 20646 9612 20698
rect 9636 20646 9646 20698
rect 9646 20646 9692 20698
rect 9396 20644 9452 20646
rect 9476 20644 9532 20646
rect 9556 20644 9612 20646
rect 9636 20644 9692 20646
rect 9396 19610 9452 19612
rect 9476 19610 9532 19612
rect 9556 19610 9612 19612
rect 9636 19610 9692 19612
rect 9396 19558 9442 19610
rect 9442 19558 9452 19610
rect 9476 19558 9506 19610
rect 9506 19558 9518 19610
rect 9518 19558 9532 19610
rect 9556 19558 9570 19610
rect 9570 19558 9582 19610
rect 9582 19558 9612 19610
rect 9636 19558 9646 19610
rect 9646 19558 9692 19610
rect 9396 19556 9452 19558
rect 9476 19556 9532 19558
rect 9556 19556 9612 19558
rect 9636 19556 9692 19558
rect 9396 18522 9452 18524
rect 9476 18522 9532 18524
rect 9556 18522 9612 18524
rect 9636 18522 9692 18524
rect 9396 18470 9442 18522
rect 9442 18470 9452 18522
rect 9476 18470 9506 18522
rect 9506 18470 9518 18522
rect 9518 18470 9532 18522
rect 9556 18470 9570 18522
rect 9570 18470 9582 18522
rect 9582 18470 9612 18522
rect 9636 18470 9646 18522
rect 9646 18470 9692 18522
rect 9396 18468 9452 18470
rect 9476 18468 9532 18470
rect 9556 18468 9612 18470
rect 9636 18468 9692 18470
rect 9396 17434 9452 17436
rect 9476 17434 9532 17436
rect 9556 17434 9612 17436
rect 9636 17434 9692 17436
rect 9396 17382 9442 17434
rect 9442 17382 9452 17434
rect 9476 17382 9506 17434
rect 9506 17382 9518 17434
rect 9518 17382 9532 17434
rect 9556 17382 9570 17434
rect 9570 17382 9582 17434
rect 9582 17382 9612 17434
rect 9636 17382 9646 17434
rect 9646 17382 9692 17434
rect 9396 17380 9452 17382
rect 9476 17380 9532 17382
rect 9556 17380 9612 17382
rect 9636 17380 9692 17382
rect 9396 16346 9452 16348
rect 9476 16346 9532 16348
rect 9556 16346 9612 16348
rect 9636 16346 9692 16348
rect 9396 16294 9442 16346
rect 9442 16294 9452 16346
rect 9476 16294 9506 16346
rect 9506 16294 9518 16346
rect 9518 16294 9532 16346
rect 9556 16294 9570 16346
rect 9570 16294 9582 16346
rect 9582 16294 9612 16346
rect 9636 16294 9646 16346
rect 9646 16294 9692 16346
rect 9396 16292 9452 16294
rect 9476 16292 9532 16294
rect 9556 16292 9612 16294
rect 9636 16292 9692 16294
rect 9396 15258 9452 15260
rect 9476 15258 9532 15260
rect 9556 15258 9612 15260
rect 9636 15258 9692 15260
rect 9396 15206 9442 15258
rect 9442 15206 9452 15258
rect 9476 15206 9506 15258
rect 9506 15206 9518 15258
rect 9518 15206 9532 15258
rect 9556 15206 9570 15258
rect 9570 15206 9582 15258
rect 9582 15206 9612 15258
rect 9636 15206 9646 15258
rect 9646 15206 9692 15258
rect 9396 15204 9452 15206
rect 9476 15204 9532 15206
rect 9556 15204 9612 15206
rect 9636 15204 9692 15206
rect 5176 11450 5232 11452
rect 5256 11450 5312 11452
rect 5336 11450 5392 11452
rect 5416 11450 5472 11452
rect 5176 11398 5222 11450
rect 5222 11398 5232 11450
rect 5256 11398 5286 11450
rect 5286 11398 5298 11450
rect 5298 11398 5312 11450
rect 5336 11398 5350 11450
rect 5350 11398 5362 11450
rect 5362 11398 5392 11450
rect 5416 11398 5426 11450
rect 5426 11398 5472 11450
rect 5176 11396 5232 11398
rect 5256 11396 5312 11398
rect 5336 11396 5392 11398
rect 5416 11396 5472 11398
rect 5176 10362 5232 10364
rect 5256 10362 5312 10364
rect 5336 10362 5392 10364
rect 5416 10362 5472 10364
rect 5176 10310 5222 10362
rect 5222 10310 5232 10362
rect 5256 10310 5286 10362
rect 5286 10310 5298 10362
rect 5298 10310 5312 10362
rect 5336 10310 5350 10362
rect 5350 10310 5362 10362
rect 5362 10310 5392 10362
rect 5416 10310 5426 10362
rect 5426 10310 5472 10362
rect 5176 10308 5232 10310
rect 5256 10308 5312 10310
rect 5336 10308 5392 10310
rect 5416 10308 5472 10310
rect 5176 9274 5232 9276
rect 5256 9274 5312 9276
rect 5336 9274 5392 9276
rect 5416 9274 5472 9276
rect 5176 9222 5222 9274
rect 5222 9222 5232 9274
rect 5256 9222 5286 9274
rect 5286 9222 5298 9274
rect 5298 9222 5312 9274
rect 5336 9222 5350 9274
rect 5350 9222 5362 9274
rect 5362 9222 5392 9274
rect 5416 9222 5426 9274
rect 5426 9222 5472 9274
rect 5176 9220 5232 9222
rect 5256 9220 5312 9222
rect 5336 9220 5392 9222
rect 5416 9220 5472 9222
rect 5176 8186 5232 8188
rect 5256 8186 5312 8188
rect 5336 8186 5392 8188
rect 5416 8186 5472 8188
rect 5176 8134 5222 8186
rect 5222 8134 5232 8186
rect 5256 8134 5286 8186
rect 5286 8134 5298 8186
rect 5298 8134 5312 8186
rect 5336 8134 5350 8186
rect 5350 8134 5362 8186
rect 5362 8134 5392 8186
rect 5416 8134 5426 8186
rect 5426 8134 5472 8186
rect 5176 8132 5232 8134
rect 5256 8132 5312 8134
rect 5336 8132 5392 8134
rect 5416 8132 5472 8134
rect 5176 7098 5232 7100
rect 5256 7098 5312 7100
rect 5336 7098 5392 7100
rect 5416 7098 5472 7100
rect 5176 7046 5222 7098
rect 5222 7046 5232 7098
rect 5256 7046 5286 7098
rect 5286 7046 5298 7098
rect 5298 7046 5312 7098
rect 5336 7046 5350 7098
rect 5350 7046 5362 7098
rect 5362 7046 5392 7098
rect 5416 7046 5426 7098
rect 5426 7046 5472 7098
rect 5176 7044 5232 7046
rect 5256 7044 5312 7046
rect 5336 7044 5392 7046
rect 5416 7044 5472 7046
rect 5176 6010 5232 6012
rect 5256 6010 5312 6012
rect 5336 6010 5392 6012
rect 5416 6010 5472 6012
rect 5176 5958 5222 6010
rect 5222 5958 5232 6010
rect 5256 5958 5286 6010
rect 5286 5958 5298 6010
rect 5298 5958 5312 6010
rect 5336 5958 5350 6010
rect 5350 5958 5362 6010
rect 5362 5958 5392 6010
rect 5416 5958 5426 6010
rect 5426 5958 5472 6010
rect 5176 5956 5232 5958
rect 5256 5956 5312 5958
rect 5336 5956 5392 5958
rect 5416 5956 5472 5958
rect 5176 4922 5232 4924
rect 5256 4922 5312 4924
rect 5336 4922 5392 4924
rect 5416 4922 5472 4924
rect 5176 4870 5222 4922
rect 5222 4870 5232 4922
rect 5256 4870 5286 4922
rect 5286 4870 5298 4922
rect 5298 4870 5312 4922
rect 5336 4870 5350 4922
rect 5350 4870 5362 4922
rect 5362 4870 5392 4922
rect 5416 4870 5426 4922
rect 5426 4870 5472 4922
rect 5176 4868 5232 4870
rect 5256 4868 5312 4870
rect 5336 4868 5392 4870
rect 5416 4868 5472 4870
rect 5176 3834 5232 3836
rect 5256 3834 5312 3836
rect 5336 3834 5392 3836
rect 5416 3834 5472 3836
rect 5176 3782 5222 3834
rect 5222 3782 5232 3834
rect 5256 3782 5286 3834
rect 5286 3782 5298 3834
rect 5298 3782 5312 3834
rect 5336 3782 5350 3834
rect 5350 3782 5362 3834
rect 5362 3782 5392 3834
rect 5416 3782 5426 3834
rect 5426 3782 5472 3834
rect 5176 3780 5232 3782
rect 5256 3780 5312 3782
rect 5336 3780 5392 3782
rect 5416 3780 5472 3782
rect 5176 2746 5232 2748
rect 5256 2746 5312 2748
rect 5336 2746 5392 2748
rect 5416 2746 5472 2748
rect 5176 2694 5222 2746
rect 5222 2694 5232 2746
rect 5256 2694 5286 2746
rect 5286 2694 5298 2746
rect 5298 2694 5312 2746
rect 5336 2694 5350 2746
rect 5350 2694 5362 2746
rect 5362 2694 5392 2746
rect 5416 2694 5426 2746
rect 5426 2694 5472 2746
rect 5176 2692 5232 2694
rect 5256 2692 5312 2694
rect 5336 2692 5392 2694
rect 5416 2692 5472 2694
rect 9396 14170 9452 14172
rect 9476 14170 9532 14172
rect 9556 14170 9612 14172
rect 9636 14170 9692 14172
rect 9396 14118 9442 14170
rect 9442 14118 9452 14170
rect 9476 14118 9506 14170
rect 9506 14118 9518 14170
rect 9518 14118 9532 14170
rect 9556 14118 9570 14170
rect 9570 14118 9582 14170
rect 9582 14118 9612 14170
rect 9636 14118 9646 14170
rect 9646 14118 9692 14170
rect 9396 14116 9452 14118
rect 9476 14116 9532 14118
rect 9556 14116 9612 14118
rect 9636 14116 9692 14118
rect 9396 13082 9452 13084
rect 9476 13082 9532 13084
rect 9556 13082 9612 13084
rect 9636 13082 9692 13084
rect 9396 13030 9442 13082
rect 9442 13030 9452 13082
rect 9476 13030 9506 13082
rect 9506 13030 9518 13082
rect 9518 13030 9532 13082
rect 9556 13030 9570 13082
rect 9570 13030 9582 13082
rect 9582 13030 9612 13082
rect 9636 13030 9646 13082
rect 9646 13030 9692 13082
rect 9396 13028 9452 13030
rect 9476 13028 9532 13030
rect 9556 13028 9612 13030
rect 9636 13028 9692 13030
rect 9396 11994 9452 11996
rect 9476 11994 9532 11996
rect 9556 11994 9612 11996
rect 9636 11994 9692 11996
rect 9396 11942 9442 11994
rect 9442 11942 9452 11994
rect 9476 11942 9506 11994
rect 9506 11942 9518 11994
rect 9518 11942 9532 11994
rect 9556 11942 9570 11994
rect 9570 11942 9582 11994
rect 9582 11942 9612 11994
rect 9636 11942 9646 11994
rect 9646 11942 9692 11994
rect 9396 11940 9452 11942
rect 9476 11940 9532 11942
rect 9556 11940 9612 11942
rect 9636 11940 9692 11942
rect 9396 10906 9452 10908
rect 9476 10906 9532 10908
rect 9556 10906 9612 10908
rect 9636 10906 9692 10908
rect 9396 10854 9442 10906
rect 9442 10854 9452 10906
rect 9476 10854 9506 10906
rect 9506 10854 9518 10906
rect 9518 10854 9532 10906
rect 9556 10854 9570 10906
rect 9570 10854 9582 10906
rect 9582 10854 9612 10906
rect 9636 10854 9646 10906
rect 9646 10854 9692 10906
rect 9396 10852 9452 10854
rect 9476 10852 9532 10854
rect 9556 10852 9612 10854
rect 9636 10852 9692 10854
rect 13617 32122 13673 32124
rect 13697 32122 13753 32124
rect 13777 32122 13833 32124
rect 13857 32122 13913 32124
rect 13617 32070 13663 32122
rect 13663 32070 13673 32122
rect 13697 32070 13727 32122
rect 13727 32070 13739 32122
rect 13739 32070 13753 32122
rect 13777 32070 13791 32122
rect 13791 32070 13803 32122
rect 13803 32070 13833 32122
rect 13857 32070 13867 32122
rect 13867 32070 13913 32122
rect 13617 32068 13673 32070
rect 13697 32068 13753 32070
rect 13777 32068 13833 32070
rect 13857 32068 13913 32070
rect 13617 31034 13673 31036
rect 13697 31034 13753 31036
rect 13777 31034 13833 31036
rect 13857 31034 13913 31036
rect 13617 30982 13663 31034
rect 13663 30982 13673 31034
rect 13697 30982 13727 31034
rect 13727 30982 13739 31034
rect 13739 30982 13753 31034
rect 13777 30982 13791 31034
rect 13791 30982 13803 31034
rect 13803 30982 13833 31034
rect 13857 30982 13867 31034
rect 13867 30982 13913 31034
rect 13617 30980 13673 30982
rect 13697 30980 13753 30982
rect 13777 30980 13833 30982
rect 13857 30980 13913 30982
rect 13617 29946 13673 29948
rect 13697 29946 13753 29948
rect 13777 29946 13833 29948
rect 13857 29946 13913 29948
rect 13617 29894 13663 29946
rect 13663 29894 13673 29946
rect 13697 29894 13727 29946
rect 13727 29894 13739 29946
rect 13739 29894 13753 29946
rect 13777 29894 13791 29946
rect 13791 29894 13803 29946
rect 13803 29894 13833 29946
rect 13857 29894 13867 29946
rect 13867 29894 13913 29946
rect 13617 29892 13673 29894
rect 13697 29892 13753 29894
rect 13777 29892 13833 29894
rect 13857 29892 13913 29894
rect 13617 28858 13673 28860
rect 13697 28858 13753 28860
rect 13777 28858 13833 28860
rect 13857 28858 13913 28860
rect 13617 28806 13663 28858
rect 13663 28806 13673 28858
rect 13697 28806 13727 28858
rect 13727 28806 13739 28858
rect 13739 28806 13753 28858
rect 13777 28806 13791 28858
rect 13791 28806 13803 28858
rect 13803 28806 13833 28858
rect 13857 28806 13867 28858
rect 13867 28806 13913 28858
rect 13617 28804 13673 28806
rect 13697 28804 13753 28806
rect 13777 28804 13833 28806
rect 13857 28804 13913 28806
rect 13617 27770 13673 27772
rect 13697 27770 13753 27772
rect 13777 27770 13833 27772
rect 13857 27770 13913 27772
rect 13617 27718 13663 27770
rect 13663 27718 13673 27770
rect 13697 27718 13727 27770
rect 13727 27718 13739 27770
rect 13739 27718 13753 27770
rect 13777 27718 13791 27770
rect 13791 27718 13803 27770
rect 13803 27718 13833 27770
rect 13857 27718 13867 27770
rect 13867 27718 13913 27770
rect 13617 27716 13673 27718
rect 13697 27716 13753 27718
rect 13777 27716 13833 27718
rect 13857 27716 13913 27718
rect 13617 26682 13673 26684
rect 13697 26682 13753 26684
rect 13777 26682 13833 26684
rect 13857 26682 13913 26684
rect 13617 26630 13663 26682
rect 13663 26630 13673 26682
rect 13697 26630 13727 26682
rect 13727 26630 13739 26682
rect 13739 26630 13753 26682
rect 13777 26630 13791 26682
rect 13791 26630 13803 26682
rect 13803 26630 13833 26682
rect 13857 26630 13867 26682
rect 13867 26630 13913 26682
rect 13617 26628 13673 26630
rect 13697 26628 13753 26630
rect 13777 26628 13833 26630
rect 13857 26628 13913 26630
rect 13617 25594 13673 25596
rect 13697 25594 13753 25596
rect 13777 25594 13833 25596
rect 13857 25594 13913 25596
rect 13617 25542 13663 25594
rect 13663 25542 13673 25594
rect 13697 25542 13727 25594
rect 13727 25542 13739 25594
rect 13739 25542 13753 25594
rect 13777 25542 13791 25594
rect 13791 25542 13803 25594
rect 13803 25542 13833 25594
rect 13857 25542 13867 25594
rect 13867 25542 13913 25594
rect 13617 25540 13673 25542
rect 13697 25540 13753 25542
rect 13777 25540 13833 25542
rect 13857 25540 13913 25542
rect 13617 24506 13673 24508
rect 13697 24506 13753 24508
rect 13777 24506 13833 24508
rect 13857 24506 13913 24508
rect 13617 24454 13663 24506
rect 13663 24454 13673 24506
rect 13697 24454 13727 24506
rect 13727 24454 13739 24506
rect 13739 24454 13753 24506
rect 13777 24454 13791 24506
rect 13791 24454 13803 24506
rect 13803 24454 13833 24506
rect 13857 24454 13867 24506
rect 13867 24454 13913 24506
rect 13617 24452 13673 24454
rect 13697 24452 13753 24454
rect 13777 24452 13833 24454
rect 13857 24452 13913 24454
rect 9396 9818 9452 9820
rect 9476 9818 9532 9820
rect 9556 9818 9612 9820
rect 9636 9818 9692 9820
rect 9396 9766 9442 9818
rect 9442 9766 9452 9818
rect 9476 9766 9506 9818
rect 9506 9766 9518 9818
rect 9518 9766 9532 9818
rect 9556 9766 9570 9818
rect 9570 9766 9582 9818
rect 9582 9766 9612 9818
rect 9636 9766 9646 9818
rect 9646 9766 9692 9818
rect 9396 9764 9452 9766
rect 9476 9764 9532 9766
rect 9556 9764 9612 9766
rect 9636 9764 9692 9766
rect 9396 8730 9452 8732
rect 9476 8730 9532 8732
rect 9556 8730 9612 8732
rect 9636 8730 9692 8732
rect 9396 8678 9442 8730
rect 9442 8678 9452 8730
rect 9476 8678 9506 8730
rect 9506 8678 9518 8730
rect 9518 8678 9532 8730
rect 9556 8678 9570 8730
rect 9570 8678 9582 8730
rect 9582 8678 9612 8730
rect 9636 8678 9646 8730
rect 9646 8678 9692 8730
rect 9396 8676 9452 8678
rect 9476 8676 9532 8678
rect 9556 8676 9612 8678
rect 9636 8676 9692 8678
rect 9396 7642 9452 7644
rect 9476 7642 9532 7644
rect 9556 7642 9612 7644
rect 9636 7642 9692 7644
rect 9396 7590 9442 7642
rect 9442 7590 9452 7642
rect 9476 7590 9506 7642
rect 9506 7590 9518 7642
rect 9518 7590 9532 7642
rect 9556 7590 9570 7642
rect 9570 7590 9582 7642
rect 9582 7590 9612 7642
rect 9636 7590 9646 7642
rect 9646 7590 9692 7642
rect 9396 7588 9452 7590
rect 9476 7588 9532 7590
rect 9556 7588 9612 7590
rect 9636 7588 9692 7590
rect 9396 6554 9452 6556
rect 9476 6554 9532 6556
rect 9556 6554 9612 6556
rect 9636 6554 9692 6556
rect 9396 6502 9442 6554
rect 9442 6502 9452 6554
rect 9476 6502 9506 6554
rect 9506 6502 9518 6554
rect 9518 6502 9532 6554
rect 9556 6502 9570 6554
rect 9570 6502 9582 6554
rect 9582 6502 9612 6554
rect 9636 6502 9646 6554
rect 9646 6502 9692 6554
rect 9396 6500 9452 6502
rect 9476 6500 9532 6502
rect 9556 6500 9612 6502
rect 9636 6500 9692 6502
rect 9396 5466 9452 5468
rect 9476 5466 9532 5468
rect 9556 5466 9612 5468
rect 9636 5466 9692 5468
rect 9396 5414 9442 5466
rect 9442 5414 9452 5466
rect 9476 5414 9506 5466
rect 9506 5414 9518 5466
rect 9518 5414 9532 5466
rect 9556 5414 9570 5466
rect 9570 5414 9582 5466
rect 9582 5414 9612 5466
rect 9636 5414 9646 5466
rect 9646 5414 9692 5466
rect 9396 5412 9452 5414
rect 9476 5412 9532 5414
rect 9556 5412 9612 5414
rect 9636 5412 9692 5414
rect 9396 4378 9452 4380
rect 9476 4378 9532 4380
rect 9556 4378 9612 4380
rect 9636 4378 9692 4380
rect 9396 4326 9442 4378
rect 9442 4326 9452 4378
rect 9476 4326 9506 4378
rect 9506 4326 9518 4378
rect 9518 4326 9532 4378
rect 9556 4326 9570 4378
rect 9570 4326 9582 4378
rect 9582 4326 9612 4378
rect 9636 4326 9646 4378
rect 9646 4326 9692 4378
rect 9396 4324 9452 4326
rect 9476 4324 9532 4326
rect 9556 4324 9612 4326
rect 9636 4324 9692 4326
rect 9396 3290 9452 3292
rect 9476 3290 9532 3292
rect 9556 3290 9612 3292
rect 9636 3290 9692 3292
rect 9396 3238 9442 3290
rect 9442 3238 9452 3290
rect 9476 3238 9506 3290
rect 9506 3238 9518 3290
rect 9518 3238 9532 3290
rect 9556 3238 9570 3290
rect 9570 3238 9582 3290
rect 9582 3238 9612 3290
rect 9636 3238 9646 3290
rect 9646 3238 9692 3290
rect 9396 3236 9452 3238
rect 9476 3236 9532 3238
rect 9556 3236 9612 3238
rect 9636 3236 9692 3238
rect 13617 23418 13673 23420
rect 13697 23418 13753 23420
rect 13777 23418 13833 23420
rect 13857 23418 13913 23420
rect 13617 23366 13663 23418
rect 13663 23366 13673 23418
rect 13697 23366 13727 23418
rect 13727 23366 13739 23418
rect 13739 23366 13753 23418
rect 13777 23366 13791 23418
rect 13791 23366 13803 23418
rect 13803 23366 13833 23418
rect 13857 23366 13867 23418
rect 13867 23366 13913 23418
rect 13617 23364 13673 23366
rect 13697 23364 13753 23366
rect 13777 23364 13833 23366
rect 13857 23364 13913 23366
rect 13617 22330 13673 22332
rect 13697 22330 13753 22332
rect 13777 22330 13833 22332
rect 13857 22330 13913 22332
rect 13617 22278 13663 22330
rect 13663 22278 13673 22330
rect 13697 22278 13727 22330
rect 13727 22278 13739 22330
rect 13739 22278 13753 22330
rect 13777 22278 13791 22330
rect 13791 22278 13803 22330
rect 13803 22278 13833 22330
rect 13857 22278 13867 22330
rect 13867 22278 13913 22330
rect 13617 22276 13673 22278
rect 13697 22276 13753 22278
rect 13777 22276 13833 22278
rect 13857 22276 13913 22278
rect 13617 21242 13673 21244
rect 13697 21242 13753 21244
rect 13777 21242 13833 21244
rect 13857 21242 13913 21244
rect 13617 21190 13663 21242
rect 13663 21190 13673 21242
rect 13697 21190 13727 21242
rect 13727 21190 13739 21242
rect 13739 21190 13753 21242
rect 13777 21190 13791 21242
rect 13791 21190 13803 21242
rect 13803 21190 13833 21242
rect 13857 21190 13867 21242
rect 13867 21190 13913 21242
rect 13617 21188 13673 21190
rect 13697 21188 13753 21190
rect 13777 21188 13833 21190
rect 13857 21188 13913 21190
rect 13617 20154 13673 20156
rect 13697 20154 13753 20156
rect 13777 20154 13833 20156
rect 13857 20154 13913 20156
rect 13617 20102 13663 20154
rect 13663 20102 13673 20154
rect 13697 20102 13727 20154
rect 13727 20102 13739 20154
rect 13739 20102 13753 20154
rect 13777 20102 13791 20154
rect 13791 20102 13803 20154
rect 13803 20102 13833 20154
rect 13857 20102 13867 20154
rect 13867 20102 13913 20154
rect 13617 20100 13673 20102
rect 13697 20100 13753 20102
rect 13777 20100 13833 20102
rect 13857 20100 13913 20102
rect 13617 19066 13673 19068
rect 13697 19066 13753 19068
rect 13777 19066 13833 19068
rect 13857 19066 13913 19068
rect 13617 19014 13663 19066
rect 13663 19014 13673 19066
rect 13697 19014 13727 19066
rect 13727 19014 13739 19066
rect 13739 19014 13753 19066
rect 13777 19014 13791 19066
rect 13791 19014 13803 19066
rect 13803 19014 13833 19066
rect 13857 19014 13867 19066
rect 13867 19014 13913 19066
rect 13617 19012 13673 19014
rect 13697 19012 13753 19014
rect 13777 19012 13833 19014
rect 13857 19012 13913 19014
rect 13617 17978 13673 17980
rect 13697 17978 13753 17980
rect 13777 17978 13833 17980
rect 13857 17978 13913 17980
rect 13617 17926 13663 17978
rect 13663 17926 13673 17978
rect 13697 17926 13727 17978
rect 13727 17926 13739 17978
rect 13739 17926 13753 17978
rect 13777 17926 13791 17978
rect 13791 17926 13803 17978
rect 13803 17926 13833 17978
rect 13857 17926 13867 17978
rect 13867 17926 13913 17978
rect 13617 17924 13673 17926
rect 13697 17924 13753 17926
rect 13777 17924 13833 17926
rect 13857 17924 13913 17926
rect 13617 16890 13673 16892
rect 13697 16890 13753 16892
rect 13777 16890 13833 16892
rect 13857 16890 13913 16892
rect 13617 16838 13663 16890
rect 13663 16838 13673 16890
rect 13697 16838 13727 16890
rect 13727 16838 13739 16890
rect 13739 16838 13753 16890
rect 13777 16838 13791 16890
rect 13791 16838 13803 16890
rect 13803 16838 13833 16890
rect 13857 16838 13867 16890
rect 13867 16838 13913 16890
rect 13617 16836 13673 16838
rect 13697 16836 13753 16838
rect 13777 16836 13833 16838
rect 13857 16836 13913 16838
rect 13617 15802 13673 15804
rect 13697 15802 13753 15804
rect 13777 15802 13833 15804
rect 13857 15802 13913 15804
rect 13617 15750 13663 15802
rect 13663 15750 13673 15802
rect 13697 15750 13727 15802
rect 13727 15750 13739 15802
rect 13739 15750 13753 15802
rect 13777 15750 13791 15802
rect 13791 15750 13803 15802
rect 13803 15750 13833 15802
rect 13857 15750 13867 15802
rect 13867 15750 13913 15802
rect 13617 15748 13673 15750
rect 13697 15748 13753 15750
rect 13777 15748 13833 15750
rect 13857 15748 13913 15750
rect 17837 32666 17893 32668
rect 17917 32666 17973 32668
rect 17997 32666 18053 32668
rect 18077 32666 18133 32668
rect 17837 32614 17883 32666
rect 17883 32614 17893 32666
rect 17917 32614 17947 32666
rect 17947 32614 17959 32666
rect 17959 32614 17973 32666
rect 17997 32614 18011 32666
rect 18011 32614 18023 32666
rect 18023 32614 18053 32666
rect 18077 32614 18087 32666
rect 18087 32614 18133 32666
rect 17837 32612 17893 32614
rect 17917 32612 17973 32614
rect 17997 32612 18053 32614
rect 18077 32612 18133 32614
rect 13617 14714 13673 14716
rect 13697 14714 13753 14716
rect 13777 14714 13833 14716
rect 13857 14714 13913 14716
rect 13617 14662 13663 14714
rect 13663 14662 13673 14714
rect 13697 14662 13727 14714
rect 13727 14662 13739 14714
rect 13739 14662 13753 14714
rect 13777 14662 13791 14714
rect 13791 14662 13803 14714
rect 13803 14662 13833 14714
rect 13857 14662 13867 14714
rect 13867 14662 13913 14714
rect 13617 14660 13673 14662
rect 13697 14660 13753 14662
rect 13777 14660 13833 14662
rect 13857 14660 13913 14662
rect 13617 13626 13673 13628
rect 13697 13626 13753 13628
rect 13777 13626 13833 13628
rect 13857 13626 13913 13628
rect 13617 13574 13663 13626
rect 13663 13574 13673 13626
rect 13697 13574 13727 13626
rect 13727 13574 13739 13626
rect 13739 13574 13753 13626
rect 13777 13574 13791 13626
rect 13791 13574 13803 13626
rect 13803 13574 13833 13626
rect 13857 13574 13867 13626
rect 13867 13574 13913 13626
rect 13617 13572 13673 13574
rect 13697 13572 13753 13574
rect 13777 13572 13833 13574
rect 13857 13572 13913 13574
rect 13617 12538 13673 12540
rect 13697 12538 13753 12540
rect 13777 12538 13833 12540
rect 13857 12538 13913 12540
rect 13617 12486 13663 12538
rect 13663 12486 13673 12538
rect 13697 12486 13727 12538
rect 13727 12486 13739 12538
rect 13739 12486 13753 12538
rect 13777 12486 13791 12538
rect 13791 12486 13803 12538
rect 13803 12486 13833 12538
rect 13857 12486 13867 12538
rect 13867 12486 13913 12538
rect 13617 12484 13673 12486
rect 13697 12484 13753 12486
rect 13777 12484 13833 12486
rect 13857 12484 13913 12486
rect 17837 31578 17893 31580
rect 17917 31578 17973 31580
rect 17997 31578 18053 31580
rect 18077 31578 18133 31580
rect 17837 31526 17883 31578
rect 17883 31526 17893 31578
rect 17917 31526 17947 31578
rect 17947 31526 17959 31578
rect 17959 31526 17973 31578
rect 17997 31526 18011 31578
rect 18011 31526 18023 31578
rect 18023 31526 18053 31578
rect 18077 31526 18087 31578
rect 18087 31526 18133 31578
rect 17837 31524 17893 31526
rect 17917 31524 17973 31526
rect 17997 31524 18053 31526
rect 18077 31524 18133 31526
rect 22058 33210 22114 33212
rect 22138 33210 22194 33212
rect 22218 33210 22274 33212
rect 22298 33210 22354 33212
rect 22058 33158 22104 33210
rect 22104 33158 22114 33210
rect 22138 33158 22168 33210
rect 22168 33158 22180 33210
rect 22180 33158 22194 33210
rect 22218 33158 22232 33210
rect 22232 33158 22244 33210
rect 22244 33158 22274 33210
rect 22298 33158 22308 33210
rect 22308 33158 22354 33210
rect 22058 33156 22114 33158
rect 22138 33156 22194 33158
rect 22218 33156 22274 33158
rect 22298 33156 22354 33158
rect 17837 30490 17893 30492
rect 17917 30490 17973 30492
rect 17997 30490 18053 30492
rect 18077 30490 18133 30492
rect 17837 30438 17883 30490
rect 17883 30438 17893 30490
rect 17917 30438 17947 30490
rect 17947 30438 17959 30490
rect 17959 30438 17973 30490
rect 17997 30438 18011 30490
rect 18011 30438 18023 30490
rect 18023 30438 18053 30490
rect 18077 30438 18087 30490
rect 18087 30438 18133 30490
rect 17837 30436 17893 30438
rect 17917 30436 17973 30438
rect 17997 30436 18053 30438
rect 18077 30436 18133 30438
rect 17837 29402 17893 29404
rect 17917 29402 17973 29404
rect 17997 29402 18053 29404
rect 18077 29402 18133 29404
rect 17837 29350 17883 29402
rect 17883 29350 17893 29402
rect 17917 29350 17947 29402
rect 17947 29350 17959 29402
rect 17959 29350 17973 29402
rect 17997 29350 18011 29402
rect 18011 29350 18023 29402
rect 18023 29350 18053 29402
rect 18077 29350 18087 29402
rect 18087 29350 18133 29402
rect 17837 29348 17893 29350
rect 17917 29348 17973 29350
rect 17997 29348 18053 29350
rect 18077 29348 18133 29350
rect 22058 32122 22114 32124
rect 22138 32122 22194 32124
rect 22218 32122 22274 32124
rect 22298 32122 22354 32124
rect 22058 32070 22104 32122
rect 22104 32070 22114 32122
rect 22138 32070 22168 32122
rect 22168 32070 22180 32122
rect 22180 32070 22194 32122
rect 22218 32070 22232 32122
rect 22232 32070 22244 32122
rect 22244 32070 22274 32122
rect 22298 32070 22308 32122
rect 22308 32070 22354 32122
rect 22058 32068 22114 32070
rect 22138 32068 22194 32070
rect 22218 32068 22274 32070
rect 22298 32068 22354 32070
rect 30499 33210 30555 33212
rect 30579 33210 30635 33212
rect 30659 33210 30715 33212
rect 30739 33210 30795 33212
rect 30499 33158 30545 33210
rect 30545 33158 30555 33210
rect 30579 33158 30609 33210
rect 30609 33158 30621 33210
rect 30621 33158 30635 33210
rect 30659 33158 30673 33210
rect 30673 33158 30685 33210
rect 30685 33158 30715 33210
rect 30739 33158 30749 33210
rect 30749 33158 30795 33210
rect 30499 33156 30555 33158
rect 30579 33156 30635 33158
rect 30659 33156 30715 33158
rect 30739 33156 30795 33158
rect 26278 32666 26334 32668
rect 26358 32666 26414 32668
rect 26438 32666 26494 32668
rect 26518 32666 26574 32668
rect 26278 32614 26324 32666
rect 26324 32614 26334 32666
rect 26358 32614 26388 32666
rect 26388 32614 26400 32666
rect 26400 32614 26414 32666
rect 26438 32614 26452 32666
rect 26452 32614 26464 32666
rect 26464 32614 26494 32666
rect 26518 32614 26528 32666
rect 26528 32614 26574 32666
rect 26278 32612 26334 32614
rect 26358 32612 26414 32614
rect 26438 32612 26494 32614
rect 26518 32612 26574 32614
rect 34719 32666 34775 32668
rect 34799 32666 34855 32668
rect 34879 32666 34935 32668
rect 34959 32666 35015 32668
rect 34719 32614 34765 32666
rect 34765 32614 34775 32666
rect 34799 32614 34829 32666
rect 34829 32614 34841 32666
rect 34841 32614 34855 32666
rect 34879 32614 34893 32666
rect 34893 32614 34905 32666
rect 34905 32614 34935 32666
rect 34959 32614 34969 32666
rect 34969 32614 35015 32666
rect 34719 32612 34775 32614
rect 34799 32612 34855 32614
rect 34879 32612 34935 32614
rect 34959 32612 35015 32614
rect 17837 28314 17893 28316
rect 17917 28314 17973 28316
rect 17997 28314 18053 28316
rect 18077 28314 18133 28316
rect 17837 28262 17883 28314
rect 17883 28262 17893 28314
rect 17917 28262 17947 28314
rect 17947 28262 17959 28314
rect 17959 28262 17973 28314
rect 17997 28262 18011 28314
rect 18011 28262 18023 28314
rect 18023 28262 18053 28314
rect 18077 28262 18087 28314
rect 18087 28262 18133 28314
rect 17837 28260 17893 28262
rect 17917 28260 17973 28262
rect 17997 28260 18053 28262
rect 18077 28260 18133 28262
rect 17837 27226 17893 27228
rect 17917 27226 17973 27228
rect 17997 27226 18053 27228
rect 18077 27226 18133 27228
rect 17837 27174 17883 27226
rect 17883 27174 17893 27226
rect 17917 27174 17947 27226
rect 17947 27174 17959 27226
rect 17959 27174 17973 27226
rect 17997 27174 18011 27226
rect 18011 27174 18023 27226
rect 18023 27174 18053 27226
rect 18077 27174 18087 27226
rect 18087 27174 18133 27226
rect 17837 27172 17893 27174
rect 17917 27172 17973 27174
rect 17997 27172 18053 27174
rect 18077 27172 18133 27174
rect 17837 26138 17893 26140
rect 17917 26138 17973 26140
rect 17997 26138 18053 26140
rect 18077 26138 18133 26140
rect 17837 26086 17883 26138
rect 17883 26086 17893 26138
rect 17917 26086 17947 26138
rect 17947 26086 17959 26138
rect 17959 26086 17973 26138
rect 17997 26086 18011 26138
rect 18011 26086 18023 26138
rect 18023 26086 18053 26138
rect 18077 26086 18087 26138
rect 18087 26086 18133 26138
rect 17837 26084 17893 26086
rect 17917 26084 17973 26086
rect 17997 26084 18053 26086
rect 18077 26084 18133 26086
rect 17837 25050 17893 25052
rect 17917 25050 17973 25052
rect 17997 25050 18053 25052
rect 18077 25050 18133 25052
rect 17837 24998 17883 25050
rect 17883 24998 17893 25050
rect 17917 24998 17947 25050
rect 17947 24998 17959 25050
rect 17959 24998 17973 25050
rect 17997 24998 18011 25050
rect 18011 24998 18023 25050
rect 18023 24998 18053 25050
rect 18077 24998 18087 25050
rect 18087 24998 18133 25050
rect 17837 24996 17893 24998
rect 17917 24996 17973 24998
rect 17997 24996 18053 24998
rect 18077 24996 18133 24998
rect 17837 23962 17893 23964
rect 17917 23962 17973 23964
rect 17997 23962 18053 23964
rect 18077 23962 18133 23964
rect 17837 23910 17883 23962
rect 17883 23910 17893 23962
rect 17917 23910 17947 23962
rect 17947 23910 17959 23962
rect 17959 23910 17973 23962
rect 17997 23910 18011 23962
rect 18011 23910 18023 23962
rect 18023 23910 18053 23962
rect 18077 23910 18087 23962
rect 18087 23910 18133 23962
rect 17837 23908 17893 23910
rect 17917 23908 17973 23910
rect 17997 23908 18053 23910
rect 18077 23908 18133 23910
rect 17837 22874 17893 22876
rect 17917 22874 17973 22876
rect 17997 22874 18053 22876
rect 18077 22874 18133 22876
rect 17837 22822 17883 22874
rect 17883 22822 17893 22874
rect 17917 22822 17947 22874
rect 17947 22822 17959 22874
rect 17959 22822 17973 22874
rect 17997 22822 18011 22874
rect 18011 22822 18023 22874
rect 18023 22822 18053 22874
rect 18077 22822 18087 22874
rect 18087 22822 18133 22874
rect 17837 22820 17893 22822
rect 17917 22820 17973 22822
rect 17997 22820 18053 22822
rect 18077 22820 18133 22822
rect 17837 21786 17893 21788
rect 17917 21786 17973 21788
rect 17997 21786 18053 21788
rect 18077 21786 18133 21788
rect 17837 21734 17883 21786
rect 17883 21734 17893 21786
rect 17917 21734 17947 21786
rect 17947 21734 17959 21786
rect 17959 21734 17973 21786
rect 17997 21734 18011 21786
rect 18011 21734 18023 21786
rect 18023 21734 18053 21786
rect 18077 21734 18087 21786
rect 18087 21734 18133 21786
rect 17837 21732 17893 21734
rect 17917 21732 17973 21734
rect 17997 21732 18053 21734
rect 18077 21732 18133 21734
rect 17837 20698 17893 20700
rect 17917 20698 17973 20700
rect 17997 20698 18053 20700
rect 18077 20698 18133 20700
rect 17837 20646 17883 20698
rect 17883 20646 17893 20698
rect 17917 20646 17947 20698
rect 17947 20646 17959 20698
rect 17959 20646 17973 20698
rect 17997 20646 18011 20698
rect 18011 20646 18023 20698
rect 18023 20646 18053 20698
rect 18077 20646 18087 20698
rect 18087 20646 18133 20698
rect 17837 20644 17893 20646
rect 17917 20644 17973 20646
rect 17997 20644 18053 20646
rect 18077 20644 18133 20646
rect 17837 19610 17893 19612
rect 17917 19610 17973 19612
rect 17997 19610 18053 19612
rect 18077 19610 18133 19612
rect 17837 19558 17883 19610
rect 17883 19558 17893 19610
rect 17917 19558 17947 19610
rect 17947 19558 17959 19610
rect 17959 19558 17973 19610
rect 17997 19558 18011 19610
rect 18011 19558 18023 19610
rect 18023 19558 18053 19610
rect 18077 19558 18087 19610
rect 18087 19558 18133 19610
rect 17837 19556 17893 19558
rect 17917 19556 17973 19558
rect 17997 19556 18053 19558
rect 18077 19556 18133 19558
rect 17837 18522 17893 18524
rect 17917 18522 17973 18524
rect 17997 18522 18053 18524
rect 18077 18522 18133 18524
rect 17837 18470 17883 18522
rect 17883 18470 17893 18522
rect 17917 18470 17947 18522
rect 17947 18470 17959 18522
rect 17959 18470 17973 18522
rect 17997 18470 18011 18522
rect 18011 18470 18023 18522
rect 18023 18470 18053 18522
rect 18077 18470 18087 18522
rect 18087 18470 18133 18522
rect 17837 18468 17893 18470
rect 17917 18468 17973 18470
rect 17997 18468 18053 18470
rect 18077 18468 18133 18470
rect 13617 11450 13673 11452
rect 13697 11450 13753 11452
rect 13777 11450 13833 11452
rect 13857 11450 13913 11452
rect 13617 11398 13663 11450
rect 13663 11398 13673 11450
rect 13697 11398 13727 11450
rect 13727 11398 13739 11450
rect 13739 11398 13753 11450
rect 13777 11398 13791 11450
rect 13791 11398 13803 11450
rect 13803 11398 13833 11450
rect 13857 11398 13867 11450
rect 13867 11398 13913 11450
rect 13617 11396 13673 11398
rect 13697 11396 13753 11398
rect 13777 11396 13833 11398
rect 13857 11396 13913 11398
rect 13617 10362 13673 10364
rect 13697 10362 13753 10364
rect 13777 10362 13833 10364
rect 13857 10362 13913 10364
rect 13617 10310 13663 10362
rect 13663 10310 13673 10362
rect 13697 10310 13727 10362
rect 13727 10310 13739 10362
rect 13739 10310 13753 10362
rect 13777 10310 13791 10362
rect 13791 10310 13803 10362
rect 13803 10310 13833 10362
rect 13857 10310 13867 10362
rect 13867 10310 13913 10362
rect 13617 10308 13673 10310
rect 13697 10308 13753 10310
rect 13777 10308 13833 10310
rect 13857 10308 13913 10310
rect 13617 9274 13673 9276
rect 13697 9274 13753 9276
rect 13777 9274 13833 9276
rect 13857 9274 13913 9276
rect 13617 9222 13663 9274
rect 13663 9222 13673 9274
rect 13697 9222 13727 9274
rect 13727 9222 13739 9274
rect 13739 9222 13753 9274
rect 13777 9222 13791 9274
rect 13791 9222 13803 9274
rect 13803 9222 13833 9274
rect 13857 9222 13867 9274
rect 13867 9222 13913 9274
rect 13617 9220 13673 9222
rect 13697 9220 13753 9222
rect 13777 9220 13833 9222
rect 13857 9220 13913 9222
rect 13617 8186 13673 8188
rect 13697 8186 13753 8188
rect 13777 8186 13833 8188
rect 13857 8186 13913 8188
rect 13617 8134 13663 8186
rect 13663 8134 13673 8186
rect 13697 8134 13727 8186
rect 13727 8134 13739 8186
rect 13739 8134 13753 8186
rect 13777 8134 13791 8186
rect 13791 8134 13803 8186
rect 13803 8134 13833 8186
rect 13857 8134 13867 8186
rect 13867 8134 13913 8186
rect 13617 8132 13673 8134
rect 13697 8132 13753 8134
rect 13777 8132 13833 8134
rect 13857 8132 13913 8134
rect 13617 7098 13673 7100
rect 13697 7098 13753 7100
rect 13777 7098 13833 7100
rect 13857 7098 13913 7100
rect 13617 7046 13663 7098
rect 13663 7046 13673 7098
rect 13697 7046 13727 7098
rect 13727 7046 13739 7098
rect 13739 7046 13753 7098
rect 13777 7046 13791 7098
rect 13791 7046 13803 7098
rect 13803 7046 13833 7098
rect 13857 7046 13867 7098
rect 13867 7046 13913 7098
rect 13617 7044 13673 7046
rect 13697 7044 13753 7046
rect 13777 7044 13833 7046
rect 13857 7044 13913 7046
rect 13617 6010 13673 6012
rect 13697 6010 13753 6012
rect 13777 6010 13833 6012
rect 13857 6010 13913 6012
rect 13617 5958 13663 6010
rect 13663 5958 13673 6010
rect 13697 5958 13727 6010
rect 13727 5958 13739 6010
rect 13739 5958 13753 6010
rect 13777 5958 13791 6010
rect 13791 5958 13803 6010
rect 13803 5958 13833 6010
rect 13857 5958 13867 6010
rect 13867 5958 13913 6010
rect 13617 5956 13673 5958
rect 13697 5956 13753 5958
rect 13777 5956 13833 5958
rect 13857 5956 13913 5958
rect 13617 4922 13673 4924
rect 13697 4922 13753 4924
rect 13777 4922 13833 4924
rect 13857 4922 13913 4924
rect 13617 4870 13663 4922
rect 13663 4870 13673 4922
rect 13697 4870 13727 4922
rect 13727 4870 13739 4922
rect 13739 4870 13753 4922
rect 13777 4870 13791 4922
rect 13791 4870 13803 4922
rect 13803 4870 13833 4922
rect 13857 4870 13867 4922
rect 13867 4870 13913 4922
rect 13617 4868 13673 4870
rect 13697 4868 13753 4870
rect 13777 4868 13833 4870
rect 13857 4868 13913 4870
rect 13617 3834 13673 3836
rect 13697 3834 13753 3836
rect 13777 3834 13833 3836
rect 13857 3834 13913 3836
rect 13617 3782 13663 3834
rect 13663 3782 13673 3834
rect 13697 3782 13727 3834
rect 13727 3782 13739 3834
rect 13739 3782 13753 3834
rect 13777 3782 13791 3834
rect 13791 3782 13803 3834
rect 13803 3782 13833 3834
rect 13857 3782 13867 3834
rect 13867 3782 13913 3834
rect 13617 3780 13673 3782
rect 13697 3780 13753 3782
rect 13777 3780 13833 3782
rect 13857 3780 13913 3782
rect 13617 2746 13673 2748
rect 13697 2746 13753 2748
rect 13777 2746 13833 2748
rect 13857 2746 13913 2748
rect 13617 2694 13663 2746
rect 13663 2694 13673 2746
rect 13697 2694 13727 2746
rect 13727 2694 13739 2746
rect 13739 2694 13753 2746
rect 13777 2694 13791 2746
rect 13791 2694 13803 2746
rect 13803 2694 13833 2746
rect 13857 2694 13867 2746
rect 13867 2694 13913 2746
rect 13617 2692 13673 2694
rect 13697 2692 13753 2694
rect 13777 2692 13833 2694
rect 13857 2692 13913 2694
rect 17837 17434 17893 17436
rect 17917 17434 17973 17436
rect 17997 17434 18053 17436
rect 18077 17434 18133 17436
rect 17837 17382 17883 17434
rect 17883 17382 17893 17434
rect 17917 17382 17947 17434
rect 17947 17382 17959 17434
rect 17959 17382 17973 17434
rect 17997 17382 18011 17434
rect 18011 17382 18023 17434
rect 18023 17382 18053 17434
rect 18077 17382 18087 17434
rect 18087 17382 18133 17434
rect 17837 17380 17893 17382
rect 17917 17380 17973 17382
rect 17997 17380 18053 17382
rect 18077 17380 18133 17382
rect 17406 12416 17462 12472
rect 17837 16346 17893 16348
rect 17917 16346 17973 16348
rect 17997 16346 18053 16348
rect 18077 16346 18133 16348
rect 17837 16294 17883 16346
rect 17883 16294 17893 16346
rect 17917 16294 17947 16346
rect 17947 16294 17959 16346
rect 17959 16294 17973 16346
rect 17997 16294 18011 16346
rect 18011 16294 18023 16346
rect 18023 16294 18053 16346
rect 18077 16294 18087 16346
rect 18087 16294 18133 16346
rect 17837 16292 17893 16294
rect 17917 16292 17973 16294
rect 17997 16292 18053 16294
rect 18077 16292 18133 16294
rect 17837 15258 17893 15260
rect 17917 15258 17973 15260
rect 17997 15258 18053 15260
rect 18077 15258 18133 15260
rect 17837 15206 17883 15258
rect 17883 15206 17893 15258
rect 17917 15206 17947 15258
rect 17947 15206 17959 15258
rect 17959 15206 17973 15258
rect 17997 15206 18011 15258
rect 18011 15206 18023 15258
rect 18023 15206 18053 15258
rect 18077 15206 18087 15258
rect 18087 15206 18133 15258
rect 17837 15204 17893 15206
rect 17917 15204 17973 15206
rect 17997 15204 18053 15206
rect 18077 15204 18133 15206
rect 17837 14170 17893 14172
rect 17917 14170 17973 14172
rect 17997 14170 18053 14172
rect 18077 14170 18133 14172
rect 17837 14118 17883 14170
rect 17883 14118 17893 14170
rect 17917 14118 17947 14170
rect 17947 14118 17959 14170
rect 17959 14118 17973 14170
rect 17997 14118 18011 14170
rect 18011 14118 18023 14170
rect 18023 14118 18053 14170
rect 18077 14118 18087 14170
rect 18087 14118 18133 14170
rect 17837 14116 17893 14118
rect 17917 14116 17973 14118
rect 17997 14116 18053 14118
rect 18077 14116 18133 14118
rect 17837 13082 17893 13084
rect 17917 13082 17973 13084
rect 17997 13082 18053 13084
rect 18077 13082 18133 13084
rect 17837 13030 17883 13082
rect 17883 13030 17893 13082
rect 17917 13030 17947 13082
rect 17947 13030 17959 13082
rect 17959 13030 17973 13082
rect 17997 13030 18011 13082
rect 18011 13030 18023 13082
rect 18023 13030 18053 13082
rect 18077 13030 18087 13082
rect 18087 13030 18133 13082
rect 17837 13028 17893 13030
rect 17917 13028 17973 13030
rect 17997 13028 18053 13030
rect 18077 13028 18133 13030
rect 17837 11994 17893 11996
rect 17917 11994 17973 11996
rect 17997 11994 18053 11996
rect 18077 11994 18133 11996
rect 17837 11942 17883 11994
rect 17883 11942 17893 11994
rect 17917 11942 17947 11994
rect 17947 11942 17959 11994
rect 17959 11942 17973 11994
rect 17997 11942 18011 11994
rect 18011 11942 18023 11994
rect 18023 11942 18053 11994
rect 18077 11942 18087 11994
rect 18087 11942 18133 11994
rect 17837 11940 17893 11942
rect 17917 11940 17973 11942
rect 17997 11940 18053 11942
rect 18077 11940 18133 11942
rect 17837 10906 17893 10908
rect 17917 10906 17973 10908
rect 17997 10906 18053 10908
rect 18077 10906 18133 10908
rect 17837 10854 17883 10906
rect 17883 10854 17893 10906
rect 17917 10854 17947 10906
rect 17947 10854 17959 10906
rect 17959 10854 17973 10906
rect 17997 10854 18011 10906
rect 18011 10854 18023 10906
rect 18023 10854 18053 10906
rect 18077 10854 18087 10906
rect 18087 10854 18133 10906
rect 17837 10852 17893 10854
rect 17917 10852 17973 10854
rect 17997 10852 18053 10854
rect 18077 10852 18133 10854
rect 22058 31034 22114 31036
rect 22138 31034 22194 31036
rect 22218 31034 22274 31036
rect 22298 31034 22354 31036
rect 22058 30982 22104 31034
rect 22104 30982 22114 31034
rect 22138 30982 22168 31034
rect 22168 30982 22180 31034
rect 22180 30982 22194 31034
rect 22218 30982 22232 31034
rect 22232 30982 22244 31034
rect 22244 30982 22274 31034
rect 22298 30982 22308 31034
rect 22308 30982 22354 31034
rect 22058 30980 22114 30982
rect 22138 30980 22194 30982
rect 22218 30980 22274 30982
rect 22298 30980 22354 30982
rect 22058 29946 22114 29948
rect 22138 29946 22194 29948
rect 22218 29946 22274 29948
rect 22298 29946 22354 29948
rect 22058 29894 22104 29946
rect 22104 29894 22114 29946
rect 22138 29894 22168 29946
rect 22168 29894 22180 29946
rect 22180 29894 22194 29946
rect 22218 29894 22232 29946
rect 22232 29894 22244 29946
rect 22244 29894 22274 29946
rect 22298 29894 22308 29946
rect 22308 29894 22354 29946
rect 22058 29892 22114 29894
rect 22138 29892 22194 29894
rect 22218 29892 22274 29894
rect 22298 29892 22354 29894
rect 22058 28858 22114 28860
rect 22138 28858 22194 28860
rect 22218 28858 22274 28860
rect 22298 28858 22354 28860
rect 22058 28806 22104 28858
rect 22104 28806 22114 28858
rect 22138 28806 22168 28858
rect 22168 28806 22180 28858
rect 22180 28806 22194 28858
rect 22218 28806 22232 28858
rect 22232 28806 22244 28858
rect 22244 28806 22274 28858
rect 22298 28806 22308 28858
rect 22308 28806 22354 28858
rect 22058 28804 22114 28806
rect 22138 28804 22194 28806
rect 22218 28804 22274 28806
rect 22298 28804 22354 28806
rect 21914 28056 21970 28112
rect 22058 27770 22114 27772
rect 22138 27770 22194 27772
rect 22218 27770 22274 27772
rect 22298 27770 22354 27772
rect 22058 27718 22104 27770
rect 22104 27718 22114 27770
rect 22138 27718 22168 27770
rect 22168 27718 22180 27770
rect 22180 27718 22194 27770
rect 22218 27718 22232 27770
rect 22232 27718 22244 27770
rect 22244 27718 22274 27770
rect 22298 27718 22308 27770
rect 22308 27718 22354 27770
rect 22058 27716 22114 27718
rect 22138 27716 22194 27718
rect 22218 27716 22274 27718
rect 22298 27716 22354 27718
rect 22058 26682 22114 26684
rect 22138 26682 22194 26684
rect 22218 26682 22274 26684
rect 22298 26682 22354 26684
rect 22058 26630 22104 26682
rect 22104 26630 22114 26682
rect 22138 26630 22168 26682
rect 22168 26630 22180 26682
rect 22180 26630 22194 26682
rect 22218 26630 22232 26682
rect 22232 26630 22244 26682
rect 22244 26630 22274 26682
rect 22298 26630 22308 26682
rect 22308 26630 22354 26682
rect 22058 26628 22114 26630
rect 22138 26628 22194 26630
rect 22218 26628 22274 26630
rect 22298 26628 22354 26630
rect 22058 25594 22114 25596
rect 22138 25594 22194 25596
rect 22218 25594 22274 25596
rect 22298 25594 22354 25596
rect 22058 25542 22104 25594
rect 22104 25542 22114 25594
rect 22138 25542 22168 25594
rect 22168 25542 22180 25594
rect 22180 25542 22194 25594
rect 22218 25542 22232 25594
rect 22232 25542 22244 25594
rect 22244 25542 22274 25594
rect 22298 25542 22308 25594
rect 22308 25542 22354 25594
rect 22058 25540 22114 25542
rect 22138 25540 22194 25542
rect 22218 25540 22274 25542
rect 22298 25540 22354 25542
rect 19798 20984 19854 21040
rect 17837 9818 17893 9820
rect 17917 9818 17973 9820
rect 17997 9818 18053 9820
rect 18077 9818 18133 9820
rect 17837 9766 17883 9818
rect 17883 9766 17893 9818
rect 17917 9766 17947 9818
rect 17947 9766 17959 9818
rect 17959 9766 17973 9818
rect 17997 9766 18011 9818
rect 18011 9766 18023 9818
rect 18023 9766 18053 9818
rect 18077 9766 18087 9818
rect 18087 9766 18133 9818
rect 17837 9764 17893 9766
rect 17917 9764 17973 9766
rect 17997 9764 18053 9766
rect 18077 9764 18133 9766
rect 17837 8730 17893 8732
rect 17917 8730 17973 8732
rect 17997 8730 18053 8732
rect 18077 8730 18133 8732
rect 17837 8678 17883 8730
rect 17883 8678 17893 8730
rect 17917 8678 17947 8730
rect 17947 8678 17959 8730
rect 17959 8678 17973 8730
rect 17997 8678 18011 8730
rect 18011 8678 18023 8730
rect 18023 8678 18053 8730
rect 18077 8678 18087 8730
rect 18087 8678 18133 8730
rect 17837 8676 17893 8678
rect 17917 8676 17973 8678
rect 17997 8676 18053 8678
rect 18077 8676 18133 8678
rect 17837 7642 17893 7644
rect 17917 7642 17973 7644
rect 17997 7642 18053 7644
rect 18077 7642 18133 7644
rect 17837 7590 17883 7642
rect 17883 7590 17893 7642
rect 17917 7590 17947 7642
rect 17947 7590 17959 7642
rect 17959 7590 17973 7642
rect 17997 7590 18011 7642
rect 18011 7590 18023 7642
rect 18023 7590 18053 7642
rect 18077 7590 18087 7642
rect 18087 7590 18133 7642
rect 17837 7588 17893 7590
rect 17917 7588 17973 7590
rect 17997 7588 18053 7590
rect 18077 7588 18133 7590
rect 17837 6554 17893 6556
rect 17917 6554 17973 6556
rect 17997 6554 18053 6556
rect 18077 6554 18133 6556
rect 17837 6502 17883 6554
rect 17883 6502 17893 6554
rect 17917 6502 17947 6554
rect 17947 6502 17959 6554
rect 17959 6502 17973 6554
rect 17997 6502 18011 6554
rect 18011 6502 18023 6554
rect 18023 6502 18053 6554
rect 18077 6502 18087 6554
rect 18087 6502 18133 6554
rect 17837 6500 17893 6502
rect 17917 6500 17973 6502
rect 17997 6500 18053 6502
rect 18077 6500 18133 6502
rect 17837 5466 17893 5468
rect 17917 5466 17973 5468
rect 17997 5466 18053 5468
rect 18077 5466 18133 5468
rect 17837 5414 17883 5466
rect 17883 5414 17893 5466
rect 17917 5414 17947 5466
rect 17947 5414 17959 5466
rect 17959 5414 17973 5466
rect 17997 5414 18011 5466
rect 18011 5414 18023 5466
rect 18023 5414 18053 5466
rect 18077 5414 18087 5466
rect 18087 5414 18133 5466
rect 17837 5412 17893 5414
rect 17917 5412 17973 5414
rect 17997 5412 18053 5414
rect 18077 5412 18133 5414
rect 26278 31578 26334 31580
rect 26358 31578 26414 31580
rect 26438 31578 26494 31580
rect 26518 31578 26574 31580
rect 26278 31526 26324 31578
rect 26324 31526 26334 31578
rect 26358 31526 26388 31578
rect 26388 31526 26400 31578
rect 26400 31526 26414 31578
rect 26438 31526 26452 31578
rect 26452 31526 26464 31578
rect 26464 31526 26494 31578
rect 26518 31526 26528 31578
rect 26528 31526 26574 31578
rect 26278 31524 26334 31526
rect 26358 31524 26414 31526
rect 26438 31524 26494 31526
rect 26518 31524 26574 31526
rect 24858 28076 24914 28112
rect 26278 30490 26334 30492
rect 26358 30490 26414 30492
rect 26438 30490 26494 30492
rect 26518 30490 26574 30492
rect 26278 30438 26324 30490
rect 26324 30438 26334 30490
rect 26358 30438 26388 30490
rect 26388 30438 26400 30490
rect 26400 30438 26414 30490
rect 26438 30438 26452 30490
rect 26452 30438 26464 30490
rect 26464 30438 26494 30490
rect 26518 30438 26528 30490
rect 26528 30438 26574 30490
rect 26278 30436 26334 30438
rect 26358 30436 26414 30438
rect 26438 30436 26494 30438
rect 26518 30436 26574 30438
rect 24858 28056 24860 28076
rect 24860 28056 24912 28076
rect 24912 28056 24914 28076
rect 26278 29402 26334 29404
rect 26358 29402 26414 29404
rect 26438 29402 26494 29404
rect 26518 29402 26574 29404
rect 26278 29350 26324 29402
rect 26324 29350 26334 29402
rect 26358 29350 26388 29402
rect 26388 29350 26400 29402
rect 26400 29350 26414 29402
rect 26438 29350 26452 29402
rect 26452 29350 26464 29402
rect 26464 29350 26494 29402
rect 26518 29350 26528 29402
rect 26528 29350 26574 29402
rect 26278 29348 26334 29350
rect 26358 29348 26414 29350
rect 26438 29348 26494 29350
rect 26518 29348 26574 29350
rect 26278 28314 26334 28316
rect 26358 28314 26414 28316
rect 26438 28314 26494 28316
rect 26518 28314 26574 28316
rect 26278 28262 26324 28314
rect 26324 28262 26334 28314
rect 26358 28262 26388 28314
rect 26388 28262 26400 28314
rect 26400 28262 26414 28314
rect 26438 28262 26452 28314
rect 26452 28262 26464 28314
rect 26464 28262 26494 28314
rect 26518 28262 26528 28314
rect 26528 28262 26574 28314
rect 26278 28260 26334 28262
rect 26358 28260 26414 28262
rect 26438 28260 26494 28262
rect 26518 28260 26574 28262
rect 22058 24506 22114 24508
rect 22138 24506 22194 24508
rect 22218 24506 22274 24508
rect 22298 24506 22354 24508
rect 22058 24454 22104 24506
rect 22104 24454 22114 24506
rect 22138 24454 22168 24506
rect 22168 24454 22180 24506
rect 22180 24454 22194 24506
rect 22218 24454 22232 24506
rect 22232 24454 22244 24506
rect 22244 24454 22274 24506
rect 22298 24454 22308 24506
rect 22308 24454 22354 24506
rect 22058 24452 22114 24454
rect 22138 24452 22194 24454
rect 22218 24452 22274 24454
rect 22298 24452 22354 24454
rect 22058 23418 22114 23420
rect 22138 23418 22194 23420
rect 22218 23418 22274 23420
rect 22298 23418 22354 23420
rect 22058 23366 22104 23418
rect 22104 23366 22114 23418
rect 22138 23366 22168 23418
rect 22168 23366 22180 23418
rect 22180 23366 22194 23418
rect 22218 23366 22232 23418
rect 22232 23366 22244 23418
rect 22244 23366 22274 23418
rect 22298 23366 22308 23418
rect 22308 23366 22354 23418
rect 22058 23364 22114 23366
rect 22138 23364 22194 23366
rect 22218 23364 22274 23366
rect 22298 23364 22354 23366
rect 22058 22330 22114 22332
rect 22138 22330 22194 22332
rect 22218 22330 22274 22332
rect 22298 22330 22354 22332
rect 22058 22278 22104 22330
rect 22104 22278 22114 22330
rect 22138 22278 22168 22330
rect 22168 22278 22180 22330
rect 22180 22278 22194 22330
rect 22218 22278 22232 22330
rect 22232 22278 22244 22330
rect 22244 22278 22274 22330
rect 22298 22278 22308 22330
rect 22308 22278 22354 22330
rect 22058 22276 22114 22278
rect 22138 22276 22194 22278
rect 22218 22276 22274 22278
rect 22298 22276 22354 22278
rect 22058 21242 22114 21244
rect 22138 21242 22194 21244
rect 22218 21242 22274 21244
rect 22298 21242 22354 21244
rect 22058 21190 22104 21242
rect 22104 21190 22114 21242
rect 22138 21190 22168 21242
rect 22168 21190 22180 21242
rect 22180 21190 22194 21242
rect 22218 21190 22232 21242
rect 22232 21190 22244 21242
rect 22244 21190 22274 21242
rect 22298 21190 22308 21242
rect 22308 21190 22354 21242
rect 22058 21188 22114 21190
rect 22138 21188 22194 21190
rect 22218 21188 22274 21190
rect 22298 21188 22354 21190
rect 22058 20154 22114 20156
rect 22138 20154 22194 20156
rect 22218 20154 22274 20156
rect 22298 20154 22354 20156
rect 22058 20102 22104 20154
rect 22104 20102 22114 20154
rect 22138 20102 22168 20154
rect 22168 20102 22180 20154
rect 22180 20102 22194 20154
rect 22218 20102 22232 20154
rect 22232 20102 22244 20154
rect 22244 20102 22274 20154
rect 22298 20102 22308 20154
rect 22308 20102 22354 20154
rect 22058 20100 22114 20102
rect 22138 20100 22194 20102
rect 22218 20100 22274 20102
rect 22298 20100 22354 20102
rect 22058 19066 22114 19068
rect 22138 19066 22194 19068
rect 22218 19066 22274 19068
rect 22298 19066 22354 19068
rect 22058 19014 22104 19066
rect 22104 19014 22114 19066
rect 22138 19014 22168 19066
rect 22168 19014 22180 19066
rect 22180 19014 22194 19066
rect 22218 19014 22232 19066
rect 22232 19014 22244 19066
rect 22244 19014 22274 19066
rect 22298 19014 22308 19066
rect 22308 19014 22354 19066
rect 22058 19012 22114 19014
rect 22138 19012 22194 19014
rect 22218 19012 22274 19014
rect 22298 19012 22354 19014
rect 22058 17978 22114 17980
rect 22138 17978 22194 17980
rect 22218 17978 22274 17980
rect 22298 17978 22354 17980
rect 22058 17926 22104 17978
rect 22104 17926 22114 17978
rect 22138 17926 22168 17978
rect 22168 17926 22180 17978
rect 22180 17926 22194 17978
rect 22218 17926 22232 17978
rect 22232 17926 22244 17978
rect 22244 17926 22274 17978
rect 22298 17926 22308 17978
rect 22308 17926 22354 17978
rect 22058 17924 22114 17926
rect 22138 17924 22194 17926
rect 22218 17924 22274 17926
rect 22298 17924 22354 17926
rect 22058 16890 22114 16892
rect 22138 16890 22194 16892
rect 22218 16890 22274 16892
rect 22298 16890 22354 16892
rect 22058 16838 22104 16890
rect 22104 16838 22114 16890
rect 22138 16838 22168 16890
rect 22168 16838 22180 16890
rect 22180 16838 22194 16890
rect 22218 16838 22232 16890
rect 22232 16838 22244 16890
rect 22244 16838 22274 16890
rect 22298 16838 22308 16890
rect 22308 16838 22354 16890
rect 22058 16836 22114 16838
rect 22138 16836 22194 16838
rect 22218 16836 22274 16838
rect 22298 16836 22354 16838
rect 22058 15802 22114 15804
rect 22138 15802 22194 15804
rect 22218 15802 22274 15804
rect 22298 15802 22354 15804
rect 22058 15750 22104 15802
rect 22104 15750 22114 15802
rect 22138 15750 22168 15802
rect 22168 15750 22180 15802
rect 22180 15750 22194 15802
rect 22218 15750 22232 15802
rect 22232 15750 22244 15802
rect 22244 15750 22274 15802
rect 22298 15750 22308 15802
rect 22308 15750 22354 15802
rect 22058 15748 22114 15750
rect 22138 15748 22194 15750
rect 22218 15748 22274 15750
rect 22298 15748 22354 15750
rect 21270 12416 21326 12472
rect 22058 14714 22114 14716
rect 22138 14714 22194 14716
rect 22218 14714 22274 14716
rect 22298 14714 22354 14716
rect 22058 14662 22104 14714
rect 22104 14662 22114 14714
rect 22138 14662 22168 14714
rect 22168 14662 22180 14714
rect 22180 14662 22194 14714
rect 22218 14662 22232 14714
rect 22232 14662 22244 14714
rect 22244 14662 22274 14714
rect 22298 14662 22308 14714
rect 22308 14662 22354 14714
rect 22058 14660 22114 14662
rect 22138 14660 22194 14662
rect 22218 14660 22274 14662
rect 22298 14660 22354 14662
rect 26278 27226 26334 27228
rect 26358 27226 26414 27228
rect 26438 27226 26494 27228
rect 26518 27226 26574 27228
rect 26278 27174 26324 27226
rect 26324 27174 26334 27226
rect 26358 27174 26388 27226
rect 26388 27174 26400 27226
rect 26400 27174 26414 27226
rect 26438 27174 26452 27226
rect 26452 27174 26464 27226
rect 26464 27174 26494 27226
rect 26518 27174 26528 27226
rect 26528 27174 26574 27226
rect 26278 27172 26334 27174
rect 26358 27172 26414 27174
rect 26438 27172 26494 27174
rect 26518 27172 26574 27174
rect 22098 13912 22154 13968
rect 22058 13626 22114 13628
rect 22138 13626 22194 13628
rect 22218 13626 22274 13628
rect 22298 13626 22354 13628
rect 22058 13574 22104 13626
rect 22104 13574 22114 13626
rect 22138 13574 22168 13626
rect 22168 13574 22180 13626
rect 22180 13574 22194 13626
rect 22218 13574 22232 13626
rect 22232 13574 22244 13626
rect 22244 13574 22274 13626
rect 22298 13574 22308 13626
rect 22308 13574 22354 13626
rect 22058 13572 22114 13574
rect 22138 13572 22194 13574
rect 22218 13572 22274 13574
rect 22298 13572 22354 13574
rect 22058 12538 22114 12540
rect 22138 12538 22194 12540
rect 22218 12538 22274 12540
rect 22298 12538 22354 12540
rect 22058 12486 22104 12538
rect 22104 12486 22114 12538
rect 22138 12486 22168 12538
rect 22168 12486 22180 12538
rect 22180 12486 22194 12538
rect 22218 12486 22232 12538
rect 22232 12486 22244 12538
rect 22244 12486 22274 12538
rect 22298 12486 22308 12538
rect 22308 12486 22354 12538
rect 22058 12484 22114 12486
rect 22138 12484 22194 12486
rect 22218 12484 22274 12486
rect 22298 12484 22354 12486
rect 26606 26324 26608 26344
rect 26608 26324 26660 26344
rect 26660 26324 26662 26344
rect 26606 26288 26662 26324
rect 26278 26138 26334 26140
rect 26358 26138 26414 26140
rect 26438 26138 26494 26140
rect 26518 26138 26574 26140
rect 26278 26086 26324 26138
rect 26324 26086 26334 26138
rect 26358 26086 26388 26138
rect 26388 26086 26400 26138
rect 26400 26086 26414 26138
rect 26438 26086 26452 26138
rect 26452 26086 26464 26138
rect 26464 26086 26494 26138
rect 26518 26086 26528 26138
rect 26528 26086 26574 26138
rect 26278 26084 26334 26086
rect 26358 26084 26414 26086
rect 26438 26084 26494 26086
rect 26518 26084 26574 26086
rect 26278 25050 26334 25052
rect 26358 25050 26414 25052
rect 26438 25050 26494 25052
rect 26518 25050 26574 25052
rect 26278 24998 26324 25050
rect 26324 24998 26334 25050
rect 26358 24998 26388 25050
rect 26388 24998 26400 25050
rect 26400 24998 26414 25050
rect 26438 24998 26452 25050
rect 26452 24998 26464 25050
rect 26464 24998 26494 25050
rect 26518 24998 26528 25050
rect 26528 24998 26574 25050
rect 26278 24996 26334 24998
rect 26358 24996 26414 24998
rect 26438 24996 26494 24998
rect 26518 24996 26574 24998
rect 26278 23962 26334 23964
rect 26358 23962 26414 23964
rect 26438 23962 26494 23964
rect 26518 23962 26574 23964
rect 26278 23910 26324 23962
rect 26324 23910 26334 23962
rect 26358 23910 26388 23962
rect 26388 23910 26400 23962
rect 26400 23910 26414 23962
rect 26438 23910 26452 23962
rect 26452 23910 26464 23962
rect 26464 23910 26494 23962
rect 26518 23910 26528 23962
rect 26528 23910 26574 23962
rect 26278 23908 26334 23910
rect 26358 23908 26414 23910
rect 26438 23908 26494 23910
rect 26518 23908 26574 23910
rect 26278 22874 26334 22876
rect 26358 22874 26414 22876
rect 26438 22874 26494 22876
rect 26518 22874 26574 22876
rect 26278 22822 26324 22874
rect 26324 22822 26334 22874
rect 26358 22822 26388 22874
rect 26388 22822 26400 22874
rect 26400 22822 26414 22874
rect 26438 22822 26452 22874
rect 26452 22822 26464 22874
rect 26464 22822 26494 22874
rect 26518 22822 26528 22874
rect 26528 22822 26574 22874
rect 26278 22820 26334 22822
rect 26358 22820 26414 22822
rect 26438 22820 26494 22822
rect 26518 22820 26574 22822
rect 27618 26288 27674 26344
rect 26278 21786 26334 21788
rect 26358 21786 26414 21788
rect 26438 21786 26494 21788
rect 26518 21786 26574 21788
rect 26278 21734 26324 21786
rect 26324 21734 26334 21786
rect 26358 21734 26388 21786
rect 26388 21734 26400 21786
rect 26400 21734 26414 21786
rect 26438 21734 26452 21786
rect 26452 21734 26464 21786
rect 26464 21734 26494 21786
rect 26518 21734 26528 21786
rect 26528 21734 26574 21786
rect 26278 21732 26334 21734
rect 26358 21732 26414 21734
rect 26438 21732 26494 21734
rect 26518 21732 26574 21734
rect 26278 20698 26334 20700
rect 26358 20698 26414 20700
rect 26438 20698 26494 20700
rect 26518 20698 26574 20700
rect 26278 20646 26324 20698
rect 26324 20646 26334 20698
rect 26358 20646 26388 20698
rect 26388 20646 26400 20698
rect 26400 20646 26414 20698
rect 26438 20646 26452 20698
rect 26452 20646 26464 20698
rect 26464 20646 26494 20698
rect 26518 20646 26528 20698
rect 26528 20646 26574 20698
rect 26278 20644 26334 20646
rect 26358 20644 26414 20646
rect 26438 20644 26494 20646
rect 26518 20644 26574 20646
rect 26278 19610 26334 19612
rect 26358 19610 26414 19612
rect 26438 19610 26494 19612
rect 26518 19610 26574 19612
rect 26278 19558 26324 19610
rect 26324 19558 26334 19610
rect 26358 19558 26388 19610
rect 26388 19558 26400 19610
rect 26400 19558 26414 19610
rect 26438 19558 26452 19610
rect 26452 19558 26464 19610
rect 26464 19558 26494 19610
rect 26518 19558 26528 19610
rect 26528 19558 26574 19610
rect 26278 19556 26334 19558
rect 26358 19556 26414 19558
rect 26438 19556 26494 19558
rect 26518 19556 26574 19558
rect 22058 11450 22114 11452
rect 22138 11450 22194 11452
rect 22218 11450 22274 11452
rect 22298 11450 22354 11452
rect 22058 11398 22104 11450
rect 22104 11398 22114 11450
rect 22138 11398 22168 11450
rect 22168 11398 22180 11450
rect 22180 11398 22194 11450
rect 22218 11398 22232 11450
rect 22232 11398 22244 11450
rect 22244 11398 22274 11450
rect 22298 11398 22308 11450
rect 22308 11398 22354 11450
rect 22058 11396 22114 11398
rect 22138 11396 22194 11398
rect 22218 11396 22274 11398
rect 22298 11396 22354 11398
rect 22058 10362 22114 10364
rect 22138 10362 22194 10364
rect 22218 10362 22274 10364
rect 22298 10362 22354 10364
rect 22058 10310 22104 10362
rect 22104 10310 22114 10362
rect 22138 10310 22168 10362
rect 22168 10310 22180 10362
rect 22180 10310 22194 10362
rect 22218 10310 22232 10362
rect 22232 10310 22244 10362
rect 22244 10310 22274 10362
rect 22298 10310 22308 10362
rect 22308 10310 22354 10362
rect 22058 10308 22114 10310
rect 22138 10308 22194 10310
rect 22218 10308 22274 10310
rect 22298 10308 22354 10310
rect 22058 9274 22114 9276
rect 22138 9274 22194 9276
rect 22218 9274 22274 9276
rect 22298 9274 22354 9276
rect 22058 9222 22104 9274
rect 22104 9222 22114 9274
rect 22138 9222 22168 9274
rect 22168 9222 22180 9274
rect 22180 9222 22194 9274
rect 22218 9222 22232 9274
rect 22232 9222 22244 9274
rect 22244 9222 22274 9274
rect 22298 9222 22308 9274
rect 22308 9222 22354 9274
rect 22058 9220 22114 9222
rect 22138 9220 22194 9222
rect 22218 9220 22274 9222
rect 22298 9220 22354 9222
rect 22058 8186 22114 8188
rect 22138 8186 22194 8188
rect 22218 8186 22274 8188
rect 22298 8186 22354 8188
rect 22058 8134 22104 8186
rect 22104 8134 22114 8186
rect 22138 8134 22168 8186
rect 22168 8134 22180 8186
rect 22180 8134 22194 8186
rect 22218 8134 22232 8186
rect 22232 8134 22244 8186
rect 22244 8134 22274 8186
rect 22298 8134 22308 8186
rect 22308 8134 22354 8186
rect 22058 8132 22114 8134
rect 22138 8132 22194 8134
rect 22218 8132 22274 8134
rect 22298 8132 22354 8134
rect 22058 7098 22114 7100
rect 22138 7098 22194 7100
rect 22218 7098 22274 7100
rect 22298 7098 22354 7100
rect 22058 7046 22104 7098
rect 22104 7046 22114 7098
rect 22138 7046 22168 7098
rect 22168 7046 22180 7098
rect 22180 7046 22194 7098
rect 22218 7046 22232 7098
rect 22232 7046 22244 7098
rect 22244 7046 22274 7098
rect 22298 7046 22308 7098
rect 22308 7046 22354 7098
rect 22058 7044 22114 7046
rect 22138 7044 22194 7046
rect 22218 7044 22274 7046
rect 22298 7044 22354 7046
rect 26278 18522 26334 18524
rect 26358 18522 26414 18524
rect 26438 18522 26494 18524
rect 26518 18522 26574 18524
rect 26278 18470 26324 18522
rect 26324 18470 26334 18522
rect 26358 18470 26388 18522
rect 26388 18470 26400 18522
rect 26400 18470 26414 18522
rect 26438 18470 26452 18522
rect 26452 18470 26464 18522
rect 26464 18470 26494 18522
rect 26518 18470 26528 18522
rect 26528 18470 26574 18522
rect 26278 18468 26334 18470
rect 26358 18468 26414 18470
rect 26438 18468 26494 18470
rect 26518 18468 26574 18470
rect 26278 17434 26334 17436
rect 26358 17434 26414 17436
rect 26438 17434 26494 17436
rect 26518 17434 26574 17436
rect 26278 17382 26324 17434
rect 26324 17382 26334 17434
rect 26358 17382 26388 17434
rect 26388 17382 26400 17434
rect 26400 17382 26414 17434
rect 26438 17382 26452 17434
rect 26452 17382 26464 17434
rect 26464 17382 26494 17434
rect 26518 17382 26528 17434
rect 26528 17382 26574 17434
rect 26278 17380 26334 17382
rect 26358 17380 26414 17382
rect 26438 17380 26494 17382
rect 26518 17380 26574 17382
rect 26278 16346 26334 16348
rect 26358 16346 26414 16348
rect 26438 16346 26494 16348
rect 26518 16346 26574 16348
rect 26278 16294 26324 16346
rect 26324 16294 26334 16346
rect 26358 16294 26388 16346
rect 26388 16294 26400 16346
rect 26400 16294 26414 16346
rect 26438 16294 26452 16346
rect 26452 16294 26464 16346
rect 26464 16294 26494 16346
rect 26518 16294 26528 16346
rect 26528 16294 26574 16346
rect 26278 16292 26334 16294
rect 26358 16292 26414 16294
rect 26438 16292 26494 16294
rect 26518 16292 26574 16294
rect 26278 15258 26334 15260
rect 26358 15258 26414 15260
rect 26438 15258 26494 15260
rect 26518 15258 26574 15260
rect 26278 15206 26324 15258
rect 26324 15206 26334 15258
rect 26358 15206 26388 15258
rect 26388 15206 26400 15258
rect 26400 15206 26414 15258
rect 26438 15206 26452 15258
rect 26452 15206 26464 15258
rect 26464 15206 26494 15258
rect 26518 15206 26528 15258
rect 26528 15206 26574 15258
rect 26278 15204 26334 15206
rect 26358 15204 26414 15206
rect 26438 15204 26494 15206
rect 26518 15204 26574 15206
rect 26278 14170 26334 14172
rect 26358 14170 26414 14172
rect 26438 14170 26494 14172
rect 26518 14170 26574 14172
rect 26278 14118 26324 14170
rect 26324 14118 26334 14170
rect 26358 14118 26388 14170
rect 26388 14118 26400 14170
rect 26400 14118 26414 14170
rect 26438 14118 26452 14170
rect 26452 14118 26464 14170
rect 26464 14118 26494 14170
rect 26518 14118 26528 14170
rect 26528 14118 26574 14170
rect 26278 14116 26334 14118
rect 26358 14116 26414 14118
rect 26438 14116 26494 14118
rect 26518 14116 26574 14118
rect 26278 13082 26334 13084
rect 26358 13082 26414 13084
rect 26438 13082 26494 13084
rect 26518 13082 26574 13084
rect 26278 13030 26324 13082
rect 26324 13030 26334 13082
rect 26358 13030 26388 13082
rect 26388 13030 26400 13082
rect 26400 13030 26414 13082
rect 26438 13030 26452 13082
rect 26452 13030 26464 13082
rect 26464 13030 26494 13082
rect 26518 13030 26528 13082
rect 26528 13030 26574 13082
rect 26278 13028 26334 13030
rect 26358 13028 26414 13030
rect 26438 13028 26494 13030
rect 26518 13028 26574 13030
rect 26278 11994 26334 11996
rect 26358 11994 26414 11996
rect 26438 11994 26494 11996
rect 26518 11994 26574 11996
rect 26278 11942 26324 11994
rect 26324 11942 26334 11994
rect 26358 11942 26388 11994
rect 26388 11942 26400 11994
rect 26400 11942 26414 11994
rect 26438 11942 26452 11994
rect 26452 11942 26464 11994
rect 26464 11942 26494 11994
rect 26518 11942 26528 11994
rect 26528 11942 26574 11994
rect 26278 11940 26334 11942
rect 26358 11940 26414 11942
rect 26438 11940 26494 11942
rect 26518 11940 26574 11942
rect 22058 6010 22114 6012
rect 22138 6010 22194 6012
rect 22218 6010 22274 6012
rect 22298 6010 22354 6012
rect 22058 5958 22104 6010
rect 22104 5958 22114 6010
rect 22138 5958 22168 6010
rect 22168 5958 22180 6010
rect 22180 5958 22194 6010
rect 22218 5958 22232 6010
rect 22232 5958 22244 6010
rect 22244 5958 22274 6010
rect 22298 5958 22308 6010
rect 22308 5958 22354 6010
rect 22058 5956 22114 5958
rect 22138 5956 22194 5958
rect 22218 5956 22274 5958
rect 22298 5956 22354 5958
rect 26278 10906 26334 10908
rect 26358 10906 26414 10908
rect 26438 10906 26494 10908
rect 26518 10906 26574 10908
rect 26278 10854 26324 10906
rect 26324 10854 26334 10906
rect 26358 10854 26388 10906
rect 26388 10854 26400 10906
rect 26400 10854 26414 10906
rect 26438 10854 26452 10906
rect 26452 10854 26464 10906
rect 26464 10854 26494 10906
rect 26518 10854 26528 10906
rect 26528 10854 26574 10906
rect 26278 10852 26334 10854
rect 26358 10852 26414 10854
rect 26438 10852 26494 10854
rect 26518 10852 26574 10854
rect 26278 9818 26334 9820
rect 26358 9818 26414 9820
rect 26438 9818 26494 9820
rect 26518 9818 26574 9820
rect 26278 9766 26324 9818
rect 26324 9766 26334 9818
rect 26358 9766 26388 9818
rect 26388 9766 26400 9818
rect 26400 9766 26414 9818
rect 26438 9766 26452 9818
rect 26452 9766 26464 9818
rect 26464 9766 26494 9818
rect 26518 9766 26528 9818
rect 26528 9766 26574 9818
rect 26278 9764 26334 9766
rect 26358 9764 26414 9766
rect 26438 9764 26494 9766
rect 26518 9764 26574 9766
rect 30102 22500 30158 22536
rect 30102 22480 30104 22500
rect 30104 22480 30156 22500
rect 30156 22480 30158 22500
rect 30499 32122 30555 32124
rect 30579 32122 30635 32124
rect 30659 32122 30715 32124
rect 30739 32122 30795 32124
rect 30499 32070 30545 32122
rect 30545 32070 30555 32122
rect 30579 32070 30609 32122
rect 30609 32070 30621 32122
rect 30621 32070 30635 32122
rect 30659 32070 30673 32122
rect 30673 32070 30685 32122
rect 30685 32070 30715 32122
rect 30739 32070 30749 32122
rect 30749 32070 30795 32122
rect 30499 32068 30555 32070
rect 30579 32068 30635 32070
rect 30659 32068 30715 32070
rect 30739 32068 30795 32070
rect 30499 31034 30555 31036
rect 30579 31034 30635 31036
rect 30659 31034 30715 31036
rect 30739 31034 30795 31036
rect 30499 30982 30545 31034
rect 30545 30982 30555 31034
rect 30579 30982 30609 31034
rect 30609 30982 30621 31034
rect 30621 30982 30635 31034
rect 30659 30982 30673 31034
rect 30673 30982 30685 31034
rect 30685 30982 30715 31034
rect 30739 30982 30749 31034
rect 30749 30982 30795 31034
rect 30499 30980 30555 30982
rect 30579 30980 30635 30982
rect 30659 30980 30715 30982
rect 30739 30980 30795 30982
rect 30499 29946 30555 29948
rect 30579 29946 30635 29948
rect 30659 29946 30715 29948
rect 30739 29946 30795 29948
rect 30499 29894 30545 29946
rect 30545 29894 30555 29946
rect 30579 29894 30609 29946
rect 30609 29894 30621 29946
rect 30621 29894 30635 29946
rect 30659 29894 30673 29946
rect 30673 29894 30685 29946
rect 30685 29894 30715 29946
rect 30739 29894 30749 29946
rect 30749 29894 30795 29946
rect 30499 29892 30555 29894
rect 30579 29892 30635 29894
rect 30659 29892 30715 29894
rect 30739 29892 30795 29894
rect 30499 28858 30555 28860
rect 30579 28858 30635 28860
rect 30659 28858 30715 28860
rect 30739 28858 30795 28860
rect 30499 28806 30545 28858
rect 30545 28806 30555 28858
rect 30579 28806 30609 28858
rect 30609 28806 30621 28858
rect 30621 28806 30635 28858
rect 30659 28806 30673 28858
rect 30673 28806 30685 28858
rect 30685 28806 30715 28858
rect 30739 28806 30749 28858
rect 30749 28806 30795 28858
rect 30499 28804 30555 28806
rect 30579 28804 30635 28806
rect 30659 28804 30715 28806
rect 30739 28804 30795 28806
rect 30499 27770 30555 27772
rect 30579 27770 30635 27772
rect 30659 27770 30715 27772
rect 30739 27770 30795 27772
rect 30499 27718 30545 27770
rect 30545 27718 30555 27770
rect 30579 27718 30609 27770
rect 30609 27718 30621 27770
rect 30621 27718 30635 27770
rect 30659 27718 30673 27770
rect 30673 27718 30685 27770
rect 30685 27718 30715 27770
rect 30739 27718 30749 27770
rect 30749 27718 30795 27770
rect 30499 27716 30555 27718
rect 30579 27716 30635 27718
rect 30659 27716 30715 27718
rect 30739 27716 30795 27718
rect 30499 26682 30555 26684
rect 30579 26682 30635 26684
rect 30659 26682 30715 26684
rect 30739 26682 30795 26684
rect 30499 26630 30545 26682
rect 30545 26630 30555 26682
rect 30579 26630 30609 26682
rect 30609 26630 30621 26682
rect 30621 26630 30635 26682
rect 30659 26630 30673 26682
rect 30673 26630 30685 26682
rect 30685 26630 30715 26682
rect 30739 26630 30749 26682
rect 30749 26630 30795 26682
rect 30499 26628 30555 26630
rect 30579 26628 30635 26630
rect 30659 26628 30715 26630
rect 30739 26628 30795 26630
rect 30499 25594 30555 25596
rect 30579 25594 30635 25596
rect 30659 25594 30715 25596
rect 30739 25594 30795 25596
rect 30499 25542 30545 25594
rect 30545 25542 30555 25594
rect 30579 25542 30609 25594
rect 30609 25542 30621 25594
rect 30621 25542 30635 25594
rect 30659 25542 30673 25594
rect 30673 25542 30685 25594
rect 30685 25542 30715 25594
rect 30739 25542 30749 25594
rect 30749 25542 30795 25594
rect 30499 25540 30555 25542
rect 30579 25540 30635 25542
rect 30659 25540 30715 25542
rect 30739 25540 30795 25542
rect 30499 24506 30555 24508
rect 30579 24506 30635 24508
rect 30659 24506 30715 24508
rect 30739 24506 30795 24508
rect 30499 24454 30545 24506
rect 30545 24454 30555 24506
rect 30579 24454 30609 24506
rect 30609 24454 30621 24506
rect 30621 24454 30635 24506
rect 30659 24454 30673 24506
rect 30673 24454 30685 24506
rect 30685 24454 30715 24506
rect 30739 24454 30749 24506
rect 30749 24454 30795 24506
rect 30499 24452 30555 24454
rect 30579 24452 30635 24454
rect 30659 24452 30715 24454
rect 30739 24452 30795 24454
rect 30499 23418 30555 23420
rect 30579 23418 30635 23420
rect 30659 23418 30715 23420
rect 30739 23418 30795 23420
rect 30499 23366 30545 23418
rect 30545 23366 30555 23418
rect 30579 23366 30609 23418
rect 30609 23366 30621 23418
rect 30621 23366 30635 23418
rect 30659 23366 30673 23418
rect 30673 23366 30685 23418
rect 30685 23366 30715 23418
rect 30739 23366 30749 23418
rect 30749 23366 30795 23418
rect 30499 23364 30555 23366
rect 30579 23364 30635 23366
rect 30659 23364 30715 23366
rect 30739 23364 30795 23366
rect 30499 22330 30555 22332
rect 30579 22330 30635 22332
rect 30659 22330 30715 22332
rect 30739 22330 30795 22332
rect 30499 22278 30545 22330
rect 30545 22278 30555 22330
rect 30579 22278 30609 22330
rect 30609 22278 30621 22330
rect 30621 22278 30635 22330
rect 30659 22278 30673 22330
rect 30673 22278 30685 22330
rect 30685 22278 30715 22330
rect 30739 22278 30749 22330
rect 30749 22278 30795 22330
rect 30499 22276 30555 22278
rect 30579 22276 30635 22278
rect 30659 22276 30715 22278
rect 30739 22276 30795 22278
rect 28446 20984 28502 21040
rect 30499 21242 30555 21244
rect 30579 21242 30635 21244
rect 30659 21242 30715 21244
rect 30739 21242 30795 21244
rect 30499 21190 30545 21242
rect 30545 21190 30555 21242
rect 30579 21190 30609 21242
rect 30609 21190 30621 21242
rect 30621 21190 30635 21242
rect 30659 21190 30673 21242
rect 30673 21190 30685 21242
rect 30685 21190 30715 21242
rect 30739 21190 30749 21242
rect 30749 21190 30795 21242
rect 30499 21188 30555 21190
rect 30579 21188 30635 21190
rect 30659 21188 30715 21190
rect 30739 21188 30795 21190
rect 31298 22516 31300 22536
rect 31300 22516 31352 22536
rect 31352 22516 31354 22536
rect 31298 22480 31354 22516
rect 34719 31578 34775 31580
rect 34799 31578 34855 31580
rect 34879 31578 34935 31580
rect 34959 31578 35015 31580
rect 34719 31526 34765 31578
rect 34765 31526 34775 31578
rect 34799 31526 34829 31578
rect 34829 31526 34841 31578
rect 34841 31526 34855 31578
rect 34879 31526 34893 31578
rect 34893 31526 34905 31578
rect 34905 31526 34935 31578
rect 34959 31526 34969 31578
rect 34969 31526 35015 31578
rect 34719 31524 34775 31526
rect 34799 31524 34855 31526
rect 34879 31524 34935 31526
rect 34959 31524 35015 31526
rect 34719 30490 34775 30492
rect 34799 30490 34855 30492
rect 34879 30490 34935 30492
rect 34959 30490 35015 30492
rect 34719 30438 34765 30490
rect 34765 30438 34775 30490
rect 34799 30438 34829 30490
rect 34829 30438 34841 30490
rect 34841 30438 34855 30490
rect 34879 30438 34893 30490
rect 34893 30438 34905 30490
rect 34905 30438 34935 30490
rect 34959 30438 34969 30490
rect 34969 30438 35015 30490
rect 34719 30436 34775 30438
rect 34799 30436 34855 30438
rect 34879 30436 34935 30438
rect 34959 30436 35015 30438
rect 34719 29402 34775 29404
rect 34799 29402 34855 29404
rect 34879 29402 34935 29404
rect 34959 29402 35015 29404
rect 34719 29350 34765 29402
rect 34765 29350 34775 29402
rect 34799 29350 34829 29402
rect 34829 29350 34841 29402
rect 34841 29350 34855 29402
rect 34879 29350 34893 29402
rect 34893 29350 34905 29402
rect 34905 29350 34935 29402
rect 34959 29350 34969 29402
rect 34969 29350 35015 29402
rect 34719 29348 34775 29350
rect 34799 29348 34855 29350
rect 34879 29348 34935 29350
rect 34959 29348 35015 29350
rect 34719 28314 34775 28316
rect 34799 28314 34855 28316
rect 34879 28314 34935 28316
rect 34959 28314 35015 28316
rect 34719 28262 34765 28314
rect 34765 28262 34775 28314
rect 34799 28262 34829 28314
rect 34829 28262 34841 28314
rect 34841 28262 34855 28314
rect 34879 28262 34893 28314
rect 34893 28262 34905 28314
rect 34905 28262 34935 28314
rect 34959 28262 34969 28314
rect 34969 28262 35015 28314
rect 34719 28260 34775 28262
rect 34799 28260 34855 28262
rect 34879 28260 34935 28262
rect 34959 28260 35015 28262
rect 34719 27226 34775 27228
rect 34799 27226 34855 27228
rect 34879 27226 34935 27228
rect 34959 27226 35015 27228
rect 34719 27174 34765 27226
rect 34765 27174 34775 27226
rect 34799 27174 34829 27226
rect 34829 27174 34841 27226
rect 34841 27174 34855 27226
rect 34879 27174 34893 27226
rect 34893 27174 34905 27226
rect 34905 27174 34935 27226
rect 34959 27174 34969 27226
rect 34969 27174 35015 27226
rect 34719 27172 34775 27174
rect 34799 27172 34855 27174
rect 34879 27172 34935 27174
rect 34959 27172 35015 27174
rect 34719 26138 34775 26140
rect 34799 26138 34855 26140
rect 34879 26138 34935 26140
rect 34959 26138 35015 26140
rect 34719 26086 34765 26138
rect 34765 26086 34775 26138
rect 34799 26086 34829 26138
rect 34829 26086 34841 26138
rect 34841 26086 34855 26138
rect 34879 26086 34893 26138
rect 34893 26086 34905 26138
rect 34905 26086 34935 26138
rect 34959 26086 34969 26138
rect 34969 26086 35015 26138
rect 34719 26084 34775 26086
rect 34799 26084 34855 26086
rect 34879 26084 34935 26086
rect 34959 26084 35015 26086
rect 34719 25050 34775 25052
rect 34799 25050 34855 25052
rect 34879 25050 34935 25052
rect 34959 25050 35015 25052
rect 34719 24998 34765 25050
rect 34765 24998 34775 25050
rect 34799 24998 34829 25050
rect 34829 24998 34841 25050
rect 34841 24998 34855 25050
rect 34879 24998 34893 25050
rect 34893 24998 34905 25050
rect 34905 24998 34935 25050
rect 34959 24998 34969 25050
rect 34969 24998 35015 25050
rect 34719 24996 34775 24998
rect 34799 24996 34855 24998
rect 34879 24996 34935 24998
rect 34959 24996 35015 24998
rect 34719 23962 34775 23964
rect 34799 23962 34855 23964
rect 34879 23962 34935 23964
rect 34959 23962 35015 23964
rect 34719 23910 34765 23962
rect 34765 23910 34775 23962
rect 34799 23910 34829 23962
rect 34829 23910 34841 23962
rect 34841 23910 34855 23962
rect 34879 23910 34893 23962
rect 34893 23910 34905 23962
rect 34905 23910 34935 23962
rect 34959 23910 34969 23962
rect 34969 23910 35015 23962
rect 34719 23908 34775 23910
rect 34799 23908 34855 23910
rect 34879 23908 34935 23910
rect 34959 23908 35015 23910
rect 30499 20154 30555 20156
rect 30579 20154 30635 20156
rect 30659 20154 30715 20156
rect 30739 20154 30795 20156
rect 30499 20102 30545 20154
rect 30545 20102 30555 20154
rect 30579 20102 30609 20154
rect 30609 20102 30621 20154
rect 30621 20102 30635 20154
rect 30659 20102 30673 20154
rect 30673 20102 30685 20154
rect 30685 20102 30715 20154
rect 30739 20102 30749 20154
rect 30749 20102 30795 20154
rect 30499 20100 30555 20102
rect 30579 20100 30635 20102
rect 30659 20100 30715 20102
rect 30739 20100 30795 20102
rect 30499 19066 30555 19068
rect 30579 19066 30635 19068
rect 30659 19066 30715 19068
rect 30739 19066 30795 19068
rect 30499 19014 30545 19066
rect 30545 19014 30555 19066
rect 30579 19014 30609 19066
rect 30609 19014 30621 19066
rect 30621 19014 30635 19066
rect 30659 19014 30673 19066
rect 30673 19014 30685 19066
rect 30685 19014 30715 19066
rect 30739 19014 30749 19066
rect 30749 19014 30795 19066
rect 30499 19012 30555 19014
rect 30579 19012 30635 19014
rect 30659 19012 30715 19014
rect 30739 19012 30795 19014
rect 30499 17978 30555 17980
rect 30579 17978 30635 17980
rect 30659 17978 30715 17980
rect 30739 17978 30795 17980
rect 30499 17926 30545 17978
rect 30545 17926 30555 17978
rect 30579 17926 30609 17978
rect 30609 17926 30621 17978
rect 30621 17926 30635 17978
rect 30659 17926 30673 17978
rect 30673 17926 30685 17978
rect 30685 17926 30715 17978
rect 30739 17926 30749 17978
rect 30749 17926 30795 17978
rect 30499 17924 30555 17926
rect 30579 17924 30635 17926
rect 30659 17924 30715 17926
rect 30739 17924 30795 17926
rect 30499 16890 30555 16892
rect 30579 16890 30635 16892
rect 30659 16890 30715 16892
rect 30739 16890 30795 16892
rect 30499 16838 30545 16890
rect 30545 16838 30555 16890
rect 30579 16838 30609 16890
rect 30609 16838 30621 16890
rect 30621 16838 30635 16890
rect 30659 16838 30673 16890
rect 30673 16838 30685 16890
rect 30685 16838 30715 16890
rect 30739 16838 30749 16890
rect 30749 16838 30795 16890
rect 30499 16836 30555 16838
rect 30579 16836 30635 16838
rect 30659 16836 30715 16838
rect 30739 16836 30795 16838
rect 27802 13932 27858 13968
rect 27802 13912 27804 13932
rect 27804 13912 27856 13932
rect 27856 13912 27858 13932
rect 26278 8730 26334 8732
rect 26358 8730 26414 8732
rect 26438 8730 26494 8732
rect 26518 8730 26574 8732
rect 26278 8678 26324 8730
rect 26324 8678 26334 8730
rect 26358 8678 26388 8730
rect 26388 8678 26400 8730
rect 26400 8678 26414 8730
rect 26438 8678 26452 8730
rect 26452 8678 26464 8730
rect 26464 8678 26494 8730
rect 26518 8678 26528 8730
rect 26528 8678 26574 8730
rect 26278 8676 26334 8678
rect 26358 8676 26414 8678
rect 26438 8676 26494 8678
rect 26518 8676 26574 8678
rect 26278 7642 26334 7644
rect 26358 7642 26414 7644
rect 26438 7642 26494 7644
rect 26518 7642 26574 7644
rect 26278 7590 26324 7642
rect 26324 7590 26334 7642
rect 26358 7590 26388 7642
rect 26388 7590 26400 7642
rect 26400 7590 26414 7642
rect 26438 7590 26452 7642
rect 26452 7590 26464 7642
rect 26464 7590 26494 7642
rect 26518 7590 26528 7642
rect 26528 7590 26574 7642
rect 26278 7588 26334 7590
rect 26358 7588 26414 7590
rect 26438 7588 26494 7590
rect 26518 7588 26574 7590
rect 26278 6554 26334 6556
rect 26358 6554 26414 6556
rect 26438 6554 26494 6556
rect 26518 6554 26574 6556
rect 26278 6502 26324 6554
rect 26324 6502 26334 6554
rect 26358 6502 26388 6554
rect 26388 6502 26400 6554
rect 26400 6502 26414 6554
rect 26438 6502 26452 6554
rect 26452 6502 26464 6554
rect 26464 6502 26494 6554
rect 26518 6502 26528 6554
rect 26528 6502 26574 6554
rect 26278 6500 26334 6502
rect 26358 6500 26414 6502
rect 26438 6500 26494 6502
rect 26518 6500 26574 6502
rect 26278 5466 26334 5468
rect 26358 5466 26414 5468
rect 26438 5466 26494 5468
rect 26518 5466 26574 5468
rect 26278 5414 26324 5466
rect 26324 5414 26334 5466
rect 26358 5414 26388 5466
rect 26388 5414 26400 5466
rect 26400 5414 26414 5466
rect 26438 5414 26452 5466
rect 26452 5414 26464 5466
rect 26464 5414 26494 5466
rect 26518 5414 26528 5466
rect 26528 5414 26574 5466
rect 26278 5412 26334 5414
rect 26358 5412 26414 5414
rect 26438 5412 26494 5414
rect 26518 5412 26574 5414
rect 22058 4922 22114 4924
rect 22138 4922 22194 4924
rect 22218 4922 22274 4924
rect 22298 4922 22354 4924
rect 22058 4870 22104 4922
rect 22104 4870 22114 4922
rect 22138 4870 22168 4922
rect 22168 4870 22180 4922
rect 22180 4870 22194 4922
rect 22218 4870 22232 4922
rect 22232 4870 22244 4922
rect 22244 4870 22274 4922
rect 22298 4870 22308 4922
rect 22308 4870 22354 4922
rect 22058 4868 22114 4870
rect 22138 4868 22194 4870
rect 22218 4868 22274 4870
rect 22298 4868 22354 4870
rect 17837 4378 17893 4380
rect 17917 4378 17973 4380
rect 17997 4378 18053 4380
rect 18077 4378 18133 4380
rect 17837 4326 17883 4378
rect 17883 4326 17893 4378
rect 17917 4326 17947 4378
rect 17947 4326 17959 4378
rect 17959 4326 17973 4378
rect 17997 4326 18011 4378
rect 18011 4326 18023 4378
rect 18023 4326 18053 4378
rect 18077 4326 18087 4378
rect 18087 4326 18133 4378
rect 17837 4324 17893 4326
rect 17917 4324 17973 4326
rect 17997 4324 18053 4326
rect 18077 4324 18133 4326
rect 17837 3290 17893 3292
rect 17917 3290 17973 3292
rect 17997 3290 18053 3292
rect 18077 3290 18133 3292
rect 17837 3238 17883 3290
rect 17883 3238 17893 3290
rect 17917 3238 17947 3290
rect 17947 3238 17959 3290
rect 17959 3238 17973 3290
rect 17997 3238 18011 3290
rect 18011 3238 18023 3290
rect 18023 3238 18053 3290
rect 18077 3238 18087 3290
rect 18087 3238 18133 3290
rect 17837 3236 17893 3238
rect 17917 3236 17973 3238
rect 17997 3236 18053 3238
rect 18077 3236 18133 3238
rect 22058 3834 22114 3836
rect 22138 3834 22194 3836
rect 22218 3834 22274 3836
rect 22298 3834 22354 3836
rect 22058 3782 22104 3834
rect 22104 3782 22114 3834
rect 22138 3782 22168 3834
rect 22168 3782 22180 3834
rect 22180 3782 22194 3834
rect 22218 3782 22232 3834
rect 22232 3782 22244 3834
rect 22244 3782 22274 3834
rect 22298 3782 22308 3834
rect 22308 3782 22354 3834
rect 22058 3780 22114 3782
rect 22138 3780 22194 3782
rect 22218 3780 22274 3782
rect 22298 3780 22354 3782
rect 22058 2746 22114 2748
rect 22138 2746 22194 2748
rect 22218 2746 22274 2748
rect 22298 2746 22354 2748
rect 22058 2694 22104 2746
rect 22104 2694 22114 2746
rect 22138 2694 22168 2746
rect 22168 2694 22180 2746
rect 22180 2694 22194 2746
rect 22218 2694 22232 2746
rect 22232 2694 22244 2746
rect 22244 2694 22274 2746
rect 22298 2694 22308 2746
rect 22308 2694 22354 2746
rect 22058 2692 22114 2694
rect 22138 2692 22194 2694
rect 22218 2692 22274 2694
rect 22298 2692 22354 2694
rect 26278 4378 26334 4380
rect 26358 4378 26414 4380
rect 26438 4378 26494 4380
rect 26518 4378 26574 4380
rect 26278 4326 26324 4378
rect 26324 4326 26334 4378
rect 26358 4326 26388 4378
rect 26388 4326 26400 4378
rect 26400 4326 26414 4378
rect 26438 4326 26452 4378
rect 26452 4326 26464 4378
rect 26464 4326 26494 4378
rect 26518 4326 26528 4378
rect 26528 4326 26574 4378
rect 26278 4324 26334 4326
rect 26358 4324 26414 4326
rect 26438 4324 26494 4326
rect 26518 4324 26574 4326
rect 30499 15802 30555 15804
rect 30579 15802 30635 15804
rect 30659 15802 30715 15804
rect 30739 15802 30795 15804
rect 30499 15750 30545 15802
rect 30545 15750 30555 15802
rect 30579 15750 30609 15802
rect 30609 15750 30621 15802
rect 30621 15750 30635 15802
rect 30659 15750 30673 15802
rect 30673 15750 30685 15802
rect 30685 15750 30715 15802
rect 30739 15750 30749 15802
rect 30749 15750 30795 15802
rect 30499 15748 30555 15750
rect 30579 15748 30635 15750
rect 30659 15748 30715 15750
rect 30739 15748 30795 15750
rect 28906 13948 28908 13968
rect 28908 13948 28960 13968
rect 28960 13948 28962 13968
rect 28906 13912 28962 13948
rect 30499 14714 30555 14716
rect 30579 14714 30635 14716
rect 30659 14714 30715 14716
rect 30739 14714 30795 14716
rect 30499 14662 30545 14714
rect 30545 14662 30555 14714
rect 30579 14662 30609 14714
rect 30609 14662 30621 14714
rect 30621 14662 30635 14714
rect 30659 14662 30673 14714
rect 30673 14662 30685 14714
rect 30685 14662 30715 14714
rect 30739 14662 30749 14714
rect 30749 14662 30795 14714
rect 30499 14660 30555 14662
rect 30579 14660 30635 14662
rect 30659 14660 30715 14662
rect 30739 14660 30795 14662
rect 30499 13626 30555 13628
rect 30579 13626 30635 13628
rect 30659 13626 30715 13628
rect 30739 13626 30795 13628
rect 30499 13574 30545 13626
rect 30545 13574 30555 13626
rect 30579 13574 30609 13626
rect 30609 13574 30621 13626
rect 30621 13574 30635 13626
rect 30659 13574 30673 13626
rect 30673 13574 30685 13626
rect 30685 13574 30715 13626
rect 30739 13574 30749 13626
rect 30749 13574 30795 13626
rect 30499 13572 30555 13574
rect 30579 13572 30635 13574
rect 30659 13572 30715 13574
rect 30739 13572 30795 13574
rect 30499 12538 30555 12540
rect 30579 12538 30635 12540
rect 30659 12538 30715 12540
rect 30739 12538 30795 12540
rect 30499 12486 30545 12538
rect 30545 12486 30555 12538
rect 30579 12486 30609 12538
rect 30609 12486 30621 12538
rect 30621 12486 30635 12538
rect 30659 12486 30673 12538
rect 30673 12486 30685 12538
rect 30685 12486 30715 12538
rect 30739 12486 30749 12538
rect 30749 12486 30795 12538
rect 30499 12484 30555 12486
rect 30579 12484 30635 12486
rect 30659 12484 30715 12486
rect 30739 12484 30795 12486
rect 30499 11450 30555 11452
rect 30579 11450 30635 11452
rect 30659 11450 30715 11452
rect 30739 11450 30795 11452
rect 30499 11398 30545 11450
rect 30545 11398 30555 11450
rect 30579 11398 30609 11450
rect 30609 11398 30621 11450
rect 30621 11398 30635 11450
rect 30659 11398 30673 11450
rect 30673 11398 30685 11450
rect 30685 11398 30715 11450
rect 30739 11398 30749 11450
rect 30749 11398 30795 11450
rect 30499 11396 30555 11398
rect 30579 11396 30635 11398
rect 30659 11396 30715 11398
rect 30739 11396 30795 11398
rect 34719 22874 34775 22876
rect 34799 22874 34855 22876
rect 34879 22874 34935 22876
rect 34959 22874 35015 22876
rect 34719 22822 34765 22874
rect 34765 22822 34775 22874
rect 34799 22822 34829 22874
rect 34829 22822 34841 22874
rect 34841 22822 34855 22874
rect 34879 22822 34893 22874
rect 34893 22822 34905 22874
rect 34905 22822 34935 22874
rect 34959 22822 34969 22874
rect 34969 22822 35015 22874
rect 34719 22820 34775 22822
rect 34799 22820 34855 22822
rect 34879 22820 34935 22822
rect 34959 22820 35015 22822
rect 34719 21786 34775 21788
rect 34799 21786 34855 21788
rect 34879 21786 34935 21788
rect 34959 21786 35015 21788
rect 34719 21734 34765 21786
rect 34765 21734 34775 21786
rect 34799 21734 34829 21786
rect 34829 21734 34841 21786
rect 34841 21734 34855 21786
rect 34879 21734 34893 21786
rect 34893 21734 34905 21786
rect 34905 21734 34935 21786
rect 34959 21734 34969 21786
rect 34969 21734 35015 21786
rect 34719 21732 34775 21734
rect 34799 21732 34855 21734
rect 34879 21732 34935 21734
rect 34959 21732 35015 21734
rect 34719 20698 34775 20700
rect 34799 20698 34855 20700
rect 34879 20698 34935 20700
rect 34959 20698 35015 20700
rect 34719 20646 34765 20698
rect 34765 20646 34775 20698
rect 34799 20646 34829 20698
rect 34829 20646 34841 20698
rect 34841 20646 34855 20698
rect 34879 20646 34893 20698
rect 34893 20646 34905 20698
rect 34905 20646 34935 20698
rect 34959 20646 34969 20698
rect 34969 20646 35015 20698
rect 34719 20644 34775 20646
rect 34799 20644 34855 20646
rect 34879 20644 34935 20646
rect 34959 20644 35015 20646
rect 34719 19610 34775 19612
rect 34799 19610 34855 19612
rect 34879 19610 34935 19612
rect 34959 19610 35015 19612
rect 34719 19558 34765 19610
rect 34765 19558 34775 19610
rect 34799 19558 34829 19610
rect 34829 19558 34841 19610
rect 34841 19558 34855 19610
rect 34879 19558 34893 19610
rect 34893 19558 34905 19610
rect 34905 19558 34935 19610
rect 34959 19558 34969 19610
rect 34969 19558 35015 19610
rect 34719 19556 34775 19558
rect 34799 19556 34855 19558
rect 34879 19556 34935 19558
rect 34959 19556 35015 19558
rect 34719 18522 34775 18524
rect 34799 18522 34855 18524
rect 34879 18522 34935 18524
rect 34959 18522 35015 18524
rect 34719 18470 34765 18522
rect 34765 18470 34775 18522
rect 34799 18470 34829 18522
rect 34829 18470 34841 18522
rect 34841 18470 34855 18522
rect 34879 18470 34893 18522
rect 34893 18470 34905 18522
rect 34905 18470 34935 18522
rect 34959 18470 34969 18522
rect 34969 18470 35015 18522
rect 34719 18468 34775 18470
rect 34799 18468 34855 18470
rect 34879 18468 34935 18470
rect 34959 18468 35015 18470
rect 34334 17856 34390 17912
rect 34719 17434 34775 17436
rect 34799 17434 34855 17436
rect 34879 17434 34935 17436
rect 34959 17434 35015 17436
rect 34719 17382 34765 17434
rect 34765 17382 34775 17434
rect 34799 17382 34829 17434
rect 34829 17382 34841 17434
rect 34841 17382 34855 17434
rect 34879 17382 34893 17434
rect 34893 17382 34905 17434
rect 34905 17382 34935 17434
rect 34959 17382 34969 17434
rect 34969 17382 35015 17434
rect 34719 17380 34775 17382
rect 34799 17380 34855 17382
rect 34879 17380 34935 17382
rect 34959 17380 35015 17382
rect 34719 16346 34775 16348
rect 34799 16346 34855 16348
rect 34879 16346 34935 16348
rect 34959 16346 35015 16348
rect 34719 16294 34765 16346
rect 34765 16294 34775 16346
rect 34799 16294 34829 16346
rect 34829 16294 34841 16346
rect 34841 16294 34855 16346
rect 34879 16294 34893 16346
rect 34893 16294 34905 16346
rect 34905 16294 34935 16346
rect 34959 16294 34969 16346
rect 34969 16294 35015 16346
rect 34719 16292 34775 16294
rect 34799 16292 34855 16294
rect 34879 16292 34935 16294
rect 34959 16292 35015 16294
rect 34719 15258 34775 15260
rect 34799 15258 34855 15260
rect 34879 15258 34935 15260
rect 34959 15258 35015 15260
rect 34719 15206 34765 15258
rect 34765 15206 34775 15258
rect 34799 15206 34829 15258
rect 34829 15206 34841 15258
rect 34841 15206 34855 15258
rect 34879 15206 34893 15258
rect 34893 15206 34905 15258
rect 34905 15206 34935 15258
rect 34959 15206 34969 15258
rect 34969 15206 35015 15258
rect 34719 15204 34775 15206
rect 34799 15204 34855 15206
rect 34879 15204 34935 15206
rect 34959 15204 35015 15206
rect 34719 14170 34775 14172
rect 34799 14170 34855 14172
rect 34879 14170 34935 14172
rect 34959 14170 35015 14172
rect 34719 14118 34765 14170
rect 34765 14118 34775 14170
rect 34799 14118 34829 14170
rect 34829 14118 34841 14170
rect 34841 14118 34855 14170
rect 34879 14118 34893 14170
rect 34893 14118 34905 14170
rect 34905 14118 34935 14170
rect 34959 14118 34969 14170
rect 34969 14118 35015 14170
rect 34719 14116 34775 14118
rect 34799 14116 34855 14118
rect 34879 14116 34935 14118
rect 34959 14116 35015 14118
rect 30499 10362 30555 10364
rect 30579 10362 30635 10364
rect 30659 10362 30715 10364
rect 30739 10362 30795 10364
rect 30499 10310 30545 10362
rect 30545 10310 30555 10362
rect 30579 10310 30609 10362
rect 30609 10310 30621 10362
rect 30621 10310 30635 10362
rect 30659 10310 30673 10362
rect 30673 10310 30685 10362
rect 30685 10310 30715 10362
rect 30739 10310 30749 10362
rect 30749 10310 30795 10362
rect 30499 10308 30555 10310
rect 30579 10308 30635 10310
rect 30659 10308 30715 10310
rect 30739 10308 30795 10310
rect 30499 9274 30555 9276
rect 30579 9274 30635 9276
rect 30659 9274 30715 9276
rect 30739 9274 30795 9276
rect 30499 9222 30545 9274
rect 30545 9222 30555 9274
rect 30579 9222 30609 9274
rect 30609 9222 30621 9274
rect 30621 9222 30635 9274
rect 30659 9222 30673 9274
rect 30673 9222 30685 9274
rect 30685 9222 30715 9274
rect 30739 9222 30749 9274
rect 30749 9222 30795 9274
rect 30499 9220 30555 9222
rect 30579 9220 30635 9222
rect 30659 9220 30715 9222
rect 30739 9220 30795 9222
rect 34719 13082 34775 13084
rect 34799 13082 34855 13084
rect 34879 13082 34935 13084
rect 34959 13082 35015 13084
rect 34719 13030 34765 13082
rect 34765 13030 34775 13082
rect 34799 13030 34829 13082
rect 34829 13030 34841 13082
rect 34841 13030 34855 13082
rect 34879 13030 34893 13082
rect 34893 13030 34905 13082
rect 34905 13030 34935 13082
rect 34959 13030 34969 13082
rect 34969 13030 35015 13082
rect 34719 13028 34775 13030
rect 34799 13028 34855 13030
rect 34879 13028 34935 13030
rect 34959 13028 35015 13030
rect 34719 11994 34775 11996
rect 34799 11994 34855 11996
rect 34879 11994 34935 11996
rect 34959 11994 35015 11996
rect 34719 11942 34765 11994
rect 34765 11942 34775 11994
rect 34799 11942 34829 11994
rect 34829 11942 34841 11994
rect 34841 11942 34855 11994
rect 34879 11942 34893 11994
rect 34893 11942 34905 11994
rect 34905 11942 34935 11994
rect 34959 11942 34969 11994
rect 34969 11942 35015 11994
rect 34719 11940 34775 11942
rect 34799 11940 34855 11942
rect 34879 11940 34935 11942
rect 34959 11940 35015 11942
rect 34719 10906 34775 10908
rect 34799 10906 34855 10908
rect 34879 10906 34935 10908
rect 34959 10906 35015 10908
rect 34719 10854 34765 10906
rect 34765 10854 34775 10906
rect 34799 10854 34829 10906
rect 34829 10854 34841 10906
rect 34841 10854 34855 10906
rect 34879 10854 34893 10906
rect 34893 10854 34905 10906
rect 34905 10854 34935 10906
rect 34959 10854 34969 10906
rect 34969 10854 35015 10906
rect 34719 10852 34775 10854
rect 34799 10852 34855 10854
rect 34879 10852 34935 10854
rect 34959 10852 35015 10854
rect 30499 8186 30555 8188
rect 30579 8186 30635 8188
rect 30659 8186 30715 8188
rect 30739 8186 30795 8188
rect 30499 8134 30545 8186
rect 30545 8134 30555 8186
rect 30579 8134 30609 8186
rect 30609 8134 30621 8186
rect 30621 8134 30635 8186
rect 30659 8134 30673 8186
rect 30673 8134 30685 8186
rect 30685 8134 30715 8186
rect 30739 8134 30749 8186
rect 30749 8134 30795 8186
rect 30499 8132 30555 8134
rect 30579 8132 30635 8134
rect 30659 8132 30715 8134
rect 30739 8132 30795 8134
rect 26278 3290 26334 3292
rect 26358 3290 26414 3292
rect 26438 3290 26494 3292
rect 26518 3290 26574 3292
rect 26278 3238 26324 3290
rect 26324 3238 26334 3290
rect 26358 3238 26388 3290
rect 26388 3238 26400 3290
rect 26400 3238 26414 3290
rect 26438 3238 26452 3290
rect 26452 3238 26464 3290
rect 26464 3238 26494 3290
rect 26518 3238 26528 3290
rect 26528 3238 26574 3290
rect 26278 3236 26334 3238
rect 26358 3236 26414 3238
rect 26438 3236 26494 3238
rect 26518 3236 26574 3238
rect 30499 7098 30555 7100
rect 30579 7098 30635 7100
rect 30659 7098 30715 7100
rect 30739 7098 30795 7100
rect 30499 7046 30545 7098
rect 30545 7046 30555 7098
rect 30579 7046 30609 7098
rect 30609 7046 30621 7098
rect 30621 7046 30635 7098
rect 30659 7046 30673 7098
rect 30673 7046 30685 7098
rect 30685 7046 30715 7098
rect 30739 7046 30749 7098
rect 30749 7046 30795 7098
rect 30499 7044 30555 7046
rect 30579 7044 30635 7046
rect 30659 7044 30715 7046
rect 30739 7044 30795 7046
rect 34719 9818 34775 9820
rect 34799 9818 34855 9820
rect 34879 9818 34935 9820
rect 34959 9818 35015 9820
rect 34719 9766 34765 9818
rect 34765 9766 34775 9818
rect 34799 9766 34829 9818
rect 34829 9766 34841 9818
rect 34841 9766 34855 9818
rect 34879 9766 34893 9818
rect 34893 9766 34905 9818
rect 34905 9766 34935 9818
rect 34959 9766 34969 9818
rect 34969 9766 35015 9818
rect 34719 9764 34775 9766
rect 34799 9764 34855 9766
rect 34879 9764 34935 9766
rect 34959 9764 35015 9766
rect 34719 8730 34775 8732
rect 34799 8730 34855 8732
rect 34879 8730 34935 8732
rect 34959 8730 35015 8732
rect 34719 8678 34765 8730
rect 34765 8678 34775 8730
rect 34799 8678 34829 8730
rect 34829 8678 34841 8730
rect 34841 8678 34855 8730
rect 34879 8678 34893 8730
rect 34893 8678 34905 8730
rect 34905 8678 34935 8730
rect 34959 8678 34969 8730
rect 34969 8678 35015 8730
rect 34719 8676 34775 8678
rect 34799 8676 34855 8678
rect 34879 8676 34935 8678
rect 34959 8676 35015 8678
rect 34719 7642 34775 7644
rect 34799 7642 34855 7644
rect 34879 7642 34935 7644
rect 34959 7642 35015 7644
rect 34719 7590 34765 7642
rect 34765 7590 34775 7642
rect 34799 7590 34829 7642
rect 34829 7590 34841 7642
rect 34841 7590 34855 7642
rect 34879 7590 34893 7642
rect 34893 7590 34905 7642
rect 34905 7590 34935 7642
rect 34959 7590 34969 7642
rect 34969 7590 35015 7642
rect 34719 7588 34775 7590
rect 34799 7588 34855 7590
rect 34879 7588 34935 7590
rect 34959 7588 35015 7590
rect 34719 6554 34775 6556
rect 34799 6554 34855 6556
rect 34879 6554 34935 6556
rect 34959 6554 35015 6556
rect 34719 6502 34765 6554
rect 34765 6502 34775 6554
rect 34799 6502 34829 6554
rect 34829 6502 34841 6554
rect 34841 6502 34855 6554
rect 34879 6502 34893 6554
rect 34893 6502 34905 6554
rect 34905 6502 34935 6554
rect 34959 6502 34969 6554
rect 34969 6502 35015 6554
rect 34719 6500 34775 6502
rect 34799 6500 34855 6502
rect 34879 6500 34935 6502
rect 34959 6500 35015 6502
rect 30499 6010 30555 6012
rect 30579 6010 30635 6012
rect 30659 6010 30715 6012
rect 30739 6010 30795 6012
rect 30499 5958 30545 6010
rect 30545 5958 30555 6010
rect 30579 5958 30609 6010
rect 30609 5958 30621 6010
rect 30621 5958 30635 6010
rect 30659 5958 30673 6010
rect 30673 5958 30685 6010
rect 30685 5958 30715 6010
rect 30739 5958 30749 6010
rect 30749 5958 30795 6010
rect 30499 5956 30555 5958
rect 30579 5956 30635 5958
rect 30659 5956 30715 5958
rect 30739 5956 30795 5958
rect 34719 5466 34775 5468
rect 34799 5466 34855 5468
rect 34879 5466 34935 5468
rect 34959 5466 35015 5468
rect 34719 5414 34765 5466
rect 34765 5414 34775 5466
rect 34799 5414 34829 5466
rect 34829 5414 34841 5466
rect 34841 5414 34855 5466
rect 34879 5414 34893 5466
rect 34893 5414 34905 5466
rect 34905 5414 34935 5466
rect 34959 5414 34969 5466
rect 34969 5414 35015 5466
rect 34719 5412 34775 5414
rect 34799 5412 34855 5414
rect 34879 5412 34935 5414
rect 34959 5412 35015 5414
rect 30499 4922 30555 4924
rect 30579 4922 30635 4924
rect 30659 4922 30715 4924
rect 30739 4922 30795 4924
rect 30499 4870 30545 4922
rect 30545 4870 30555 4922
rect 30579 4870 30609 4922
rect 30609 4870 30621 4922
rect 30621 4870 30635 4922
rect 30659 4870 30673 4922
rect 30673 4870 30685 4922
rect 30685 4870 30715 4922
rect 30739 4870 30749 4922
rect 30749 4870 30795 4922
rect 30499 4868 30555 4870
rect 30579 4868 30635 4870
rect 30659 4868 30715 4870
rect 30739 4868 30795 4870
rect 34719 4378 34775 4380
rect 34799 4378 34855 4380
rect 34879 4378 34935 4380
rect 34959 4378 35015 4380
rect 34719 4326 34765 4378
rect 34765 4326 34775 4378
rect 34799 4326 34829 4378
rect 34829 4326 34841 4378
rect 34841 4326 34855 4378
rect 34879 4326 34893 4378
rect 34893 4326 34905 4378
rect 34905 4326 34935 4378
rect 34959 4326 34969 4378
rect 34969 4326 35015 4378
rect 34719 4324 34775 4326
rect 34799 4324 34855 4326
rect 34879 4324 34935 4326
rect 34959 4324 35015 4326
rect 30499 3834 30555 3836
rect 30579 3834 30635 3836
rect 30659 3834 30715 3836
rect 30739 3834 30795 3836
rect 30499 3782 30545 3834
rect 30545 3782 30555 3834
rect 30579 3782 30609 3834
rect 30609 3782 30621 3834
rect 30621 3782 30635 3834
rect 30659 3782 30673 3834
rect 30673 3782 30685 3834
rect 30685 3782 30715 3834
rect 30739 3782 30749 3834
rect 30749 3782 30795 3834
rect 30499 3780 30555 3782
rect 30579 3780 30635 3782
rect 30659 3780 30715 3782
rect 30739 3780 30795 3782
rect 34719 3290 34775 3292
rect 34799 3290 34855 3292
rect 34879 3290 34935 3292
rect 34959 3290 35015 3292
rect 34719 3238 34765 3290
rect 34765 3238 34775 3290
rect 34799 3238 34829 3290
rect 34829 3238 34841 3290
rect 34841 3238 34855 3290
rect 34879 3238 34893 3290
rect 34893 3238 34905 3290
rect 34905 3238 34935 3290
rect 34959 3238 34969 3290
rect 34969 3238 35015 3290
rect 34719 3236 34775 3238
rect 34799 3236 34855 3238
rect 34879 3236 34935 3238
rect 34959 3236 35015 3238
rect 30499 2746 30555 2748
rect 30579 2746 30635 2748
rect 30659 2746 30715 2748
rect 30739 2746 30795 2748
rect 30499 2694 30545 2746
rect 30545 2694 30555 2746
rect 30579 2694 30609 2746
rect 30609 2694 30621 2746
rect 30621 2694 30635 2746
rect 30659 2694 30673 2746
rect 30673 2694 30685 2746
rect 30685 2694 30715 2746
rect 30739 2694 30749 2746
rect 30749 2694 30795 2746
rect 30499 2692 30555 2694
rect 30579 2692 30635 2694
rect 30659 2692 30715 2694
rect 30739 2692 30795 2694
rect 9396 2202 9452 2204
rect 9476 2202 9532 2204
rect 9556 2202 9612 2204
rect 9636 2202 9692 2204
rect 9396 2150 9442 2202
rect 9442 2150 9452 2202
rect 9476 2150 9506 2202
rect 9506 2150 9518 2202
rect 9518 2150 9532 2202
rect 9556 2150 9570 2202
rect 9570 2150 9582 2202
rect 9582 2150 9612 2202
rect 9636 2150 9646 2202
rect 9646 2150 9692 2202
rect 9396 2148 9452 2150
rect 9476 2148 9532 2150
rect 9556 2148 9612 2150
rect 9636 2148 9692 2150
rect 17837 2202 17893 2204
rect 17917 2202 17973 2204
rect 17997 2202 18053 2204
rect 18077 2202 18133 2204
rect 17837 2150 17883 2202
rect 17883 2150 17893 2202
rect 17917 2150 17947 2202
rect 17947 2150 17959 2202
rect 17959 2150 17973 2202
rect 17997 2150 18011 2202
rect 18011 2150 18023 2202
rect 18023 2150 18053 2202
rect 18077 2150 18087 2202
rect 18087 2150 18133 2202
rect 17837 2148 17893 2150
rect 17917 2148 17973 2150
rect 17997 2148 18053 2150
rect 18077 2148 18133 2150
rect 26278 2202 26334 2204
rect 26358 2202 26414 2204
rect 26438 2202 26494 2204
rect 26518 2202 26574 2204
rect 26278 2150 26324 2202
rect 26324 2150 26334 2202
rect 26358 2150 26388 2202
rect 26388 2150 26400 2202
rect 26400 2150 26414 2202
rect 26438 2150 26452 2202
rect 26452 2150 26464 2202
rect 26464 2150 26494 2202
rect 26518 2150 26528 2202
rect 26528 2150 26574 2202
rect 26278 2148 26334 2150
rect 26358 2148 26414 2150
rect 26438 2148 26494 2150
rect 26518 2148 26574 2150
rect 34719 2202 34775 2204
rect 34799 2202 34855 2204
rect 34879 2202 34935 2204
rect 34959 2202 35015 2204
rect 34719 2150 34765 2202
rect 34765 2150 34775 2202
rect 34799 2150 34829 2202
rect 34829 2150 34841 2202
rect 34841 2150 34855 2202
rect 34879 2150 34893 2202
rect 34893 2150 34905 2202
rect 34905 2150 34935 2202
rect 34959 2150 34969 2202
rect 34969 2150 35015 2202
rect 34719 2148 34775 2150
rect 34799 2148 34855 2150
rect 34879 2148 34935 2150
rect 34959 2148 35015 2150
<< metal3 >>
rect 9386 33760 9702 33761
rect 9386 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9702 33760
rect 9386 33695 9702 33696
rect 17827 33760 18143 33761
rect 17827 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18143 33760
rect 17827 33695 18143 33696
rect 26268 33760 26584 33761
rect 26268 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26584 33760
rect 26268 33695 26584 33696
rect 34709 33760 35025 33761
rect 34709 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35025 33760
rect 34709 33695 35025 33696
rect 5166 33216 5482 33217
rect 5166 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5482 33216
rect 5166 33151 5482 33152
rect 13607 33216 13923 33217
rect 13607 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13923 33216
rect 13607 33151 13923 33152
rect 22048 33216 22364 33217
rect 22048 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22364 33216
rect 22048 33151 22364 33152
rect 30489 33216 30805 33217
rect 30489 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30805 33216
rect 30489 33151 30805 33152
rect 9386 32672 9702 32673
rect 9386 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9702 32672
rect 9386 32607 9702 32608
rect 17827 32672 18143 32673
rect 17827 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18143 32672
rect 17827 32607 18143 32608
rect 26268 32672 26584 32673
rect 26268 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26584 32672
rect 26268 32607 26584 32608
rect 34709 32672 35025 32673
rect 34709 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35025 32672
rect 34709 32607 35025 32608
rect 5166 32128 5482 32129
rect 5166 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5482 32128
rect 5166 32063 5482 32064
rect 13607 32128 13923 32129
rect 13607 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13923 32128
rect 13607 32063 13923 32064
rect 22048 32128 22364 32129
rect 22048 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22364 32128
rect 22048 32063 22364 32064
rect 30489 32128 30805 32129
rect 30489 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30805 32128
rect 30489 32063 30805 32064
rect 9386 31584 9702 31585
rect 9386 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9702 31584
rect 9386 31519 9702 31520
rect 17827 31584 18143 31585
rect 17827 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18143 31584
rect 17827 31519 18143 31520
rect 26268 31584 26584 31585
rect 26268 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26584 31584
rect 26268 31519 26584 31520
rect 34709 31584 35025 31585
rect 34709 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35025 31584
rect 34709 31519 35025 31520
rect 5166 31040 5482 31041
rect 5166 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5482 31040
rect 5166 30975 5482 30976
rect 13607 31040 13923 31041
rect 13607 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13923 31040
rect 13607 30975 13923 30976
rect 22048 31040 22364 31041
rect 22048 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22364 31040
rect 22048 30975 22364 30976
rect 30489 31040 30805 31041
rect 30489 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30805 31040
rect 30489 30975 30805 30976
rect 9386 30496 9702 30497
rect 9386 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9702 30496
rect 9386 30431 9702 30432
rect 17827 30496 18143 30497
rect 17827 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18143 30496
rect 17827 30431 18143 30432
rect 26268 30496 26584 30497
rect 26268 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26584 30496
rect 26268 30431 26584 30432
rect 34709 30496 35025 30497
rect 34709 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35025 30496
rect 34709 30431 35025 30432
rect 5166 29952 5482 29953
rect 5166 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5482 29952
rect 5166 29887 5482 29888
rect 13607 29952 13923 29953
rect 13607 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13923 29952
rect 13607 29887 13923 29888
rect 22048 29952 22364 29953
rect 22048 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22364 29952
rect 22048 29887 22364 29888
rect 30489 29952 30805 29953
rect 30489 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30805 29952
rect 30489 29887 30805 29888
rect 9386 29408 9702 29409
rect 9386 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9702 29408
rect 9386 29343 9702 29344
rect 17827 29408 18143 29409
rect 17827 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18143 29408
rect 17827 29343 18143 29344
rect 26268 29408 26584 29409
rect 26268 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26584 29408
rect 26268 29343 26584 29344
rect 34709 29408 35025 29409
rect 34709 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35025 29408
rect 34709 29343 35025 29344
rect 5166 28864 5482 28865
rect 5166 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5482 28864
rect 5166 28799 5482 28800
rect 13607 28864 13923 28865
rect 13607 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13923 28864
rect 13607 28799 13923 28800
rect 22048 28864 22364 28865
rect 22048 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22364 28864
rect 22048 28799 22364 28800
rect 30489 28864 30805 28865
rect 30489 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30805 28864
rect 30489 28799 30805 28800
rect 9386 28320 9702 28321
rect 9386 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9702 28320
rect 9386 28255 9702 28256
rect 17827 28320 18143 28321
rect 17827 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18143 28320
rect 17827 28255 18143 28256
rect 26268 28320 26584 28321
rect 26268 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26584 28320
rect 26268 28255 26584 28256
rect 34709 28320 35025 28321
rect 34709 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35025 28320
rect 34709 28255 35025 28256
rect 21909 28114 21975 28117
rect 24853 28114 24919 28117
rect 21909 28112 24919 28114
rect 21909 28056 21914 28112
rect 21970 28056 24858 28112
rect 24914 28056 24919 28112
rect 21909 28054 24919 28056
rect 21909 28051 21975 28054
rect 24853 28051 24919 28054
rect 5166 27776 5482 27777
rect 5166 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5482 27776
rect 5166 27711 5482 27712
rect 13607 27776 13923 27777
rect 13607 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13923 27776
rect 13607 27711 13923 27712
rect 22048 27776 22364 27777
rect 22048 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22364 27776
rect 22048 27711 22364 27712
rect 30489 27776 30805 27777
rect 30489 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30805 27776
rect 30489 27711 30805 27712
rect 9386 27232 9702 27233
rect 9386 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9702 27232
rect 9386 27167 9702 27168
rect 17827 27232 18143 27233
rect 17827 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18143 27232
rect 17827 27167 18143 27168
rect 26268 27232 26584 27233
rect 26268 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26584 27232
rect 26268 27167 26584 27168
rect 34709 27232 35025 27233
rect 34709 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35025 27232
rect 34709 27167 35025 27168
rect 5166 26688 5482 26689
rect 5166 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5482 26688
rect 5166 26623 5482 26624
rect 13607 26688 13923 26689
rect 13607 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13923 26688
rect 13607 26623 13923 26624
rect 22048 26688 22364 26689
rect 22048 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22364 26688
rect 22048 26623 22364 26624
rect 30489 26688 30805 26689
rect 30489 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30805 26688
rect 30489 26623 30805 26624
rect 26601 26346 26667 26349
rect 27613 26346 27679 26349
rect 26601 26344 27679 26346
rect 26601 26288 26606 26344
rect 26662 26288 27618 26344
rect 27674 26288 27679 26344
rect 26601 26286 27679 26288
rect 26601 26283 26667 26286
rect 27613 26283 27679 26286
rect 9386 26144 9702 26145
rect 9386 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9702 26144
rect 9386 26079 9702 26080
rect 17827 26144 18143 26145
rect 17827 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18143 26144
rect 17827 26079 18143 26080
rect 26268 26144 26584 26145
rect 26268 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26584 26144
rect 26268 26079 26584 26080
rect 34709 26144 35025 26145
rect 34709 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35025 26144
rect 34709 26079 35025 26080
rect 5166 25600 5482 25601
rect 5166 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5482 25600
rect 5166 25535 5482 25536
rect 13607 25600 13923 25601
rect 13607 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13923 25600
rect 13607 25535 13923 25536
rect 22048 25600 22364 25601
rect 22048 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22364 25600
rect 22048 25535 22364 25536
rect 30489 25600 30805 25601
rect 30489 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30805 25600
rect 30489 25535 30805 25536
rect 9386 25056 9702 25057
rect 9386 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9702 25056
rect 9386 24991 9702 24992
rect 17827 25056 18143 25057
rect 17827 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18143 25056
rect 17827 24991 18143 24992
rect 26268 25056 26584 25057
rect 26268 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26584 25056
rect 26268 24991 26584 24992
rect 34709 25056 35025 25057
rect 34709 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35025 25056
rect 34709 24991 35025 24992
rect 5166 24512 5482 24513
rect 5166 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5482 24512
rect 5166 24447 5482 24448
rect 13607 24512 13923 24513
rect 13607 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13923 24512
rect 13607 24447 13923 24448
rect 22048 24512 22364 24513
rect 22048 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22364 24512
rect 22048 24447 22364 24448
rect 30489 24512 30805 24513
rect 30489 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30805 24512
rect 30489 24447 30805 24448
rect 9386 23968 9702 23969
rect 9386 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9702 23968
rect 9386 23903 9702 23904
rect 17827 23968 18143 23969
rect 17827 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18143 23968
rect 17827 23903 18143 23904
rect 26268 23968 26584 23969
rect 26268 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26584 23968
rect 26268 23903 26584 23904
rect 34709 23968 35025 23969
rect 34709 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35025 23968
rect 34709 23903 35025 23904
rect 5166 23424 5482 23425
rect 5166 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5482 23424
rect 5166 23359 5482 23360
rect 13607 23424 13923 23425
rect 13607 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13923 23424
rect 13607 23359 13923 23360
rect 22048 23424 22364 23425
rect 22048 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22364 23424
rect 22048 23359 22364 23360
rect 30489 23424 30805 23425
rect 30489 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30805 23424
rect 30489 23359 30805 23360
rect 9386 22880 9702 22881
rect 9386 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9702 22880
rect 9386 22815 9702 22816
rect 17827 22880 18143 22881
rect 17827 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18143 22880
rect 17827 22815 18143 22816
rect 26268 22880 26584 22881
rect 26268 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26584 22880
rect 26268 22815 26584 22816
rect 34709 22880 35025 22881
rect 34709 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35025 22880
rect 34709 22815 35025 22816
rect 30097 22538 30163 22541
rect 31293 22538 31359 22541
rect 30097 22536 31359 22538
rect 30097 22480 30102 22536
rect 30158 22480 31298 22536
rect 31354 22480 31359 22536
rect 30097 22478 31359 22480
rect 30097 22475 30163 22478
rect 31293 22475 31359 22478
rect 5166 22336 5482 22337
rect 5166 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5482 22336
rect 5166 22271 5482 22272
rect 13607 22336 13923 22337
rect 13607 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13923 22336
rect 13607 22271 13923 22272
rect 22048 22336 22364 22337
rect 22048 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22364 22336
rect 22048 22271 22364 22272
rect 30489 22336 30805 22337
rect 30489 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30805 22336
rect 30489 22271 30805 22272
rect 9386 21792 9702 21793
rect 9386 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9702 21792
rect 9386 21727 9702 21728
rect 17827 21792 18143 21793
rect 17827 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18143 21792
rect 17827 21727 18143 21728
rect 26268 21792 26584 21793
rect 26268 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26584 21792
rect 26268 21727 26584 21728
rect 34709 21792 35025 21793
rect 34709 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35025 21792
rect 34709 21727 35025 21728
rect 5166 21248 5482 21249
rect 5166 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5482 21248
rect 5166 21183 5482 21184
rect 13607 21248 13923 21249
rect 13607 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13923 21248
rect 13607 21183 13923 21184
rect 22048 21248 22364 21249
rect 22048 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22364 21248
rect 22048 21183 22364 21184
rect 30489 21248 30805 21249
rect 30489 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30805 21248
rect 30489 21183 30805 21184
rect 19793 21042 19859 21045
rect 28441 21042 28507 21045
rect 19793 21040 28507 21042
rect 19793 20984 19798 21040
rect 19854 20984 28446 21040
rect 28502 20984 28507 21040
rect 19793 20982 28507 20984
rect 19793 20979 19859 20982
rect 28441 20979 28507 20982
rect 9386 20704 9702 20705
rect 9386 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9702 20704
rect 9386 20639 9702 20640
rect 17827 20704 18143 20705
rect 17827 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18143 20704
rect 17827 20639 18143 20640
rect 26268 20704 26584 20705
rect 26268 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26584 20704
rect 26268 20639 26584 20640
rect 34709 20704 35025 20705
rect 34709 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35025 20704
rect 34709 20639 35025 20640
rect 5166 20160 5482 20161
rect 5166 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5482 20160
rect 5166 20095 5482 20096
rect 13607 20160 13923 20161
rect 13607 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13923 20160
rect 13607 20095 13923 20096
rect 22048 20160 22364 20161
rect 22048 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22364 20160
rect 22048 20095 22364 20096
rect 30489 20160 30805 20161
rect 30489 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30805 20160
rect 30489 20095 30805 20096
rect 4153 19954 4219 19957
rect 5349 19954 5415 19957
rect 4153 19952 5415 19954
rect 4153 19896 4158 19952
rect 4214 19896 5354 19952
rect 5410 19896 5415 19952
rect 4153 19894 5415 19896
rect 4153 19891 4219 19894
rect 5349 19891 5415 19894
rect 3693 19818 3759 19821
rect 4889 19818 4955 19821
rect 3693 19816 4955 19818
rect 3693 19760 3698 19816
rect 3754 19760 4894 19816
rect 4950 19760 4955 19816
rect 3693 19758 4955 19760
rect 3693 19755 3759 19758
rect 4889 19755 4955 19758
rect 9386 19616 9702 19617
rect 9386 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9702 19616
rect 9386 19551 9702 19552
rect 17827 19616 18143 19617
rect 17827 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18143 19616
rect 17827 19551 18143 19552
rect 26268 19616 26584 19617
rect 26268 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26584 19616
rect 26268 19551 26584 19552
rect 34709 19616 35025 19617
rect 34709 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35025 19616
rect 34709 19551 35025 19552
rect 5166 19072 5482 19073
rect 5166 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5482 19072
rect 5166 19007 5482 19008
rect 13607 19072 13923 19073
rect 13607 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13923 19072
rect 13607 19007 13923 19008
rect 22048 19072 22364 19073
rect 22048 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22364 19072
rect 22048 19007 22364 19008
rect 30489 19072 30805 19073
rect 30489 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30805 19072
rect 30489 19007 30805 19008
rect 9386 18528 9702 18529
rect 9386 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9702 18528
rect 9386 18463 9702 18464
rect 17827 18528 18143 18529
rect 17827 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18143 18528
rect 17827 18463 18143 18464
rect 26268 18528 26584 18529
rect 26268 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26584 18528
rect 26268 18463 26584 18464
rect 34709 18528 35025 18529
rect 34709 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35025 18528
rect 34709 18463 35025 18464
rect 5166 17984 5482 17985
rect 5166 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5482 17984
rect 5166 17919 5482 17920
rect 13607 17984 13923 17985
rect 13607 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13923 17984
rect 13607 17919 13923 17920
rect 22048 17984 22364 17985
rect 22048 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22364 17984
rect 22048 17919 22364 17920
rect 30489 17984 30805 17985
rect 30489 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30805 17984
rect 30489 17919 30805 17920
rect 34329 17914 34395 17917
rect 35200 17914 36000 17944
rect 34329 17912 36000 17914
rect 34329 17856 34334 17912
rect 34390 17856 36000 17912
rect 34329 17854 36000 17856
rect 34329 17851 34395 17854
rect 35200 17824 36000 17854
rect 9386 17440 9702 17441
rect 9386 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9702 17440
rect 9386 17375 9702 17376
rect 17827 17440 18143 17441
rect 17827 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18143 17440
rect 17827 17375 18143 17376
rect 26268 17440 26584 17441
rect 26268 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26584 17440
rect 26268 17375 26584 17376
rect 34709 17440 35025 17441
rect 34709 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35025 17440
rect 34709 17375 35025 17376
rect 5166 16896 5482 16897
rect 5166 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5482 16896
rect 5166 16831 5482 16832
rect 13607 16896 13923 16897
rect 13607 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13923 16896
rect 13607 16831 13923 16832
rect 22048 16896 22364 16897
rect 22048 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22364 16896
rect 22048 16831 22364 16832
rect 30489 16896 30805 16897
rect 30489 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30805 16896
rect 30489 16831 30805 16832
rect 9386 16352 9702 16353
rect 9386 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9702 16352
rect 9386 16287 9702 16288
rect 17827 16352 18143 16353
rect 17827 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18143 16352
rect 17827 16287 18143 16288
rect 26268 16352 26584 16353
rect 26268 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26584 16352
rect 26268 16287 26584 16288
rect 34709 16352 35025 16353
rect 34709 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35025 16352
rect 34709 16287 35025 16288
rect 5166 15808 5482 15809
rect 5166 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5482 15808
rect 5166 15743 5482 15744
rect 13607 15808 13923 15809
rect 13607 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13923 15808
rect 13607 15743 13923 15744
rect 22048 15808 22364 15809
rect 22048 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22364 15808
rect 22048 15743 22364 15744
rect 30489 15808 30805 15809
rect 30489 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30805 15808
rect 30489 15743 30805 15744
rect 9386 15264 9702 15265
rect 9386 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9702 15264
rect 9386 15199 9702 15200
rect 17827 15264 18143 15265
rect 17827 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18143 15264
rect 17827 15199 18143 15200
rect 26268 15264 26584 15265
rect 26268 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26584 15264
rect 26268 15199 26584 15200
rect 34709 15264 35025 15265
rect 34709 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35025 15264
rect 34709 15199 35025 15200
rect 5166 14720 5482 14721
rect 5166 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5482 14720
rect 5166 14655 5482 14656
rect 13607 14720 13923 14721
rect 13607 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13923 14720
rect 13607 14655 13923 14656
rect 22048 14720 22364 14721
rect 22048 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22364 14720
rect 22048 14655 22364 14656
rect 30489 14720 30805 14721
rect 30489 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30805 14720
rect 30489 14655 30805 14656
rect 9386 14176 9702 14177
rect 9386 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9702 14176
rect 9386 14111 9702 14112
rect 17827 14176 18143 14177
rect 17827 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18143 14176
rect 17827 14111 18143 14112
rect 26268 14176 26584 14177
rect 26268 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26584 14176
rect 26268 14111 26584 14112
rect 34709 14176 35025 14177
rect 34709 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35025 14176
rect 34709 14111 35025 14112
rect 22093 13970 22159 13973
rect 27797 13970 27863 13973
rect 28901 13970 28967 13973
rect 22093 13968 28967 13970
rect 22093 13912 22098 13968
rect 22154 13912 27802 13968
rect 27858 13912 28906 13968
rect 28962 13912 28967 13968
rect 22093 13910 28967 13912
rect 22093 13907 22159 13910
rect 27797 13907 27863 13910
rect 28901 13907 28967 13910
rect 5166 13632 5482 13633
rect 5166 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5482 13632
rect 5166 13567 5482 13568
rect 13607 13632 13923 13633
rect 13607 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13923 13632
rect 13607 13567 13923 13568
rect 22048 13632 22364 13633
rect 22048 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22364 13632
rect 22048 13567 22364 13568
rect 30489 13632 30805 13633
rect 30489 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30805 13632
rect 30489 13567 30805 13568
rect 9386 13088 9702 13089
rect 9386 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9702 13088
rect 9386 13023 9702 13024
rect 17827 13088 18143 13089
rect 17827 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18143 13088
rect 17827 13023 18143 13024
rect 26268 13088 26584 13089
rect 26268 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26584 13088
rect 26268 13023 26584 13024
rect 34709 13088 35025 13089
rect 34709 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35025 13088
rect 34709 13023 35025 13024
rect 5166 12544 5482 12545
rect 5166 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5482 12544
rect 5166 12479 5482 12480
rect 13607 12544 13923 12545
rect 13607 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13923 12544
rect 13607 12479 13923 12480
rect 22048 12544 22364 12545
rect 22048 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22364 12544
rect 22048 12479 22364 12480
rect 30489 12544 30805 12545
rect 30489 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30805 12544
rect 30489 12479 30805 12480
rect 17401 12474 17467 12477
rect 21265 12474 21331 12477
rect 17401 12472 21331 12474
rect 17401 12416 17406 12472
rect 17462 12416 21270 12472
rect 21326 12416 21331 12472
rect 17401 12414 21331 12416
rect 17401 12411 17467 12414
rect 21265 12411 21331 12414
rect 9386 12000 9702 12001
rect 9386 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9702 12000
rect 9386 11935 9702 11936
rect 17827 12000 18143 12001
rect 17827 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18143 12000
rect 17827 11935 18143 11936
rect 26268 12000 26584 12001
rect 26268 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26584 12000
rect 26268 11935 26584 11936
rect 34709 12000 35025 12001
rect 34709 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35025 12000
rect 34709 11935 35025 11936
rect 5166 11456 5482 11457
rect 5166 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5482 11456
rect 5166 11391 5482 11392
rect 13607 11456 13923 11457
rect 13607 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13923 11456
rect 13607 11391 13923 11392
rect 22048 11456 22364 11457
rect 22048 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22364 11456
rect 22048 11391 22364 11392
rect 30489 11456 30805 11457
rect 30489 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30805 11456
rect 30489 11391 30805 11392
rect 9386 10912 9702 10913
rect 9386 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9702 10912
rect 9386 10847 9702 10848
rect 17827 10912 18143 10913
rect 17827 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18143 10912
rect 17827 10847 18143 10848
rect 26268 10912 26584 10913
rect 26268 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26584 10912
rect 26268 10847 26584 10848
rect 34709 10912 35025 10913
rect 34709 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35025 10912
rect 34709 10847 35025 10848
rect 5166 10368 5482 10369
rect 5166 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5482 10368
rect 5166 10303 5482 10304
rect 13607 10368 13923 10369
rect 13607 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13923 10368
rect 13607 10303 13923 10304
rect 22048 10368 22364 10369
rect 22048 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22364 10368
rect 22048 10303 22364 10304
rect 30489 10368 30805 10369
rect 30489 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30805 10368
rect 30489 10303 30805 10304
rect 9386 9824 9702 9825
rect 9386 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9702 9824
rect 9386 9759 9702 9760
rect 17827 9824 18143 9825
rect 17827 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18143 9824
rect 17827 9759 18143 9760
rect 26268 9824 26584 9825
rect 26268 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26584 9824
rect 26268 9759 26584 9760
rect 34709 9824 35025 9825
rect 34709 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35025 9824
rect 34709 9759 35025 9760
rect 5166 9280 5482 9281
rect 5166 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5482 9280
rect 5166 9215 5482 9216
rect 13607 9280 13923 9281
rect 13607 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13923 9280
rect 13607 9215 13923 9216
rect 22048 9280 22364 9281
rect 22048 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22364 9280
rect 22048 9215 22364 9216
rect 30489 9280 30805 9281
rect 30489 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30805 9280
rect 30489 9215 30805 9216
rect 9386 8736 9702 8737
rect 9386 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9702 8736
rect 9386 8671 9702 8672
rect 17827 8736 18143 8737
rect 17827 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18143 8736
rect 17827 8671 18143 8672
rect 26268 8736 26584 8737
rect 26268 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26584 8736
rect 26268 8671 26584 8672
rect 34709 8736 35025 8737
rect 34709 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35025 8736
rect 34709 8671 35025 8672
rect 5166 8192 5482 8193
rect 5166 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5482 8192
rect 5166 8127 5482 8128
rect 13607 8192 13923 8193
rect 13607 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13923 8192
rect 13607 8127 13923 8128
rect 22048 8192 22364 8193
rect 22048 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22364 8192
rect 22048 8127 22364 8128
rect 30489 8192 30805 8193
rect 30489 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30805 8192
rect 30489 8127 30805 8128
rect 9386 7648 9702 7649
rect 9386 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9702 7648
rect 9386 7583 9702 7584
rect 17827 7648 18143 7649
rect 17827 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18143 7648
rect 17827 7583 18143 7584
rect 26268 7648 26584 7649
rect 26268 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26584 7648
rect 26268 7583 26584 7584
rect 34709 7648 35025 7649
rect 34709 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35025 7648
rect 34709 7583 35025 7584
rect 5166 7104 5482 7105
rect 5166 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5482 7104
rect 5166 7039 5482 7040
rect 13607 7104 13923 7105
rect 13607 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13923 7104
rect 13607 7039 13923 7040
rect 22048 7104 22364 7105
rect 22048 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22364 7104
rect 22048 7039 22364 7040
rect 30489 7104 30805 7105
rect 30489 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30805 7104
rect 30489 7039 30805 7040
rect 9386 6560 9702 6561
rect 9386 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9702 6560
rect 9386 6495 9702 6496
rect 17827 6560 18143 6561
rect 17827 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18143 6560
rect 17827 6495 18143 6496
rect 26268 6560 26584 6561
rect 26268 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26584 6560
rect 26268 6495 26584 6496
rect 34709 6560 35025 6561
rect 34709 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35025 6560
rect 34709 6495 35025 6496
rect 5166 6016 5482 6017
rect 5166 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5482 6016
rect 5166 5951 5482 5952
rect 13607 6016 13923 6017
rect 13607 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13923 6016
rect 13607 5951 13923 5952
rect 22048 6016 22364 6017
rect 22048 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22364 6016
rect 22048 5951 22364 5952
rect 30489 6016 30805 6017
rect 30489 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30805 6016
rect 30489 5951 30805 5952
rect 9386 5472 9702 5473
rect 9386 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9702 5472
rect 9386 5407 9702 5408
rect 17827 5472 18143 5473
rect 17827 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18143 5472
rect 17827 5407 18143 5408
rect 26268 5472 26584 5473
rect 26268 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26584 5472
rect 26268 5407 26584 5408
rect 34709 5472 35025 5473
rect 34709 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35025 5472
rect 34709 5407 35025 5408
rect 5166 4928 5482 4929
rect 5166 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5482 4928
rect 5166 4863 5482 4864
rect 13607 4928 13923 4929
rect 13607 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13923 4928
rect 13607 4863 13923 4864
rect 22048 4928 22364 4929
rect 22048 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22364 4928
rect 22048 4863 22364 4864
rect 30489 4928 30805 4929
rect 30489 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30805 4928
rect 30489 4863 30805 4864
rect 9386 4384 9702 4385
rect 9386 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9702 4384
rect 9386 4319 9702 4320
rect 17827 4384 18143 4385
rect 17827 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18143 4384
rect 17827 4319 18143 4320
rect 26268 4384 26584 4385
rect 26268 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26584 4384
rect 26268 4319 26584 4320
rect 34709 4384 35025 4385
rect 34709 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35025 4384
rect 34709 4319 35025 4320
rect 5166 3840 5482 3841
rect 5166 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5482 3840
rect 5166 3775 5482 3776
rect 13607 3840 13923 3841
rect 13607 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13923 3840
rect 13607 3775 13923 3776
rect 22048 3840 22364 3841
rect 22048 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22364 3840
rect 22048 3775 22364 3776
rect 30489 3840 30805 3841
rect 30489 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30805 3840
rect 30489 3775 30805 3776
rect 9386 3296 9702 3297
rect 9386 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9702 3296
rect 9386 3231 9702 3232
rect 17827 3296 18143 3297
rect 17827 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18143 3296
rect 17827 3231 18143 3232
rect 26268 3296 26584 3297
rect 26268 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26584 3296
rect 26268 3231 26584 3232
rect 34709 3296 35025 3297
rect 34709 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35025 3296
rect 34709 3231 35025 3232
rect 5166 2752 5482 2753
rect 5166 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5482 2752
rect 5166 2687 5482 2688
rect 13607 2752 13923 2753
rect 13607 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13923 2752
rect 13607 2687 13923 2688
rect 22048 2752 22364 2753
rect 22048 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22364 2752
rect 22048 2687 22364 2688
rect 30489 2752 30805 2753
rect 30489 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30805 2752
rect 30489 2687 30805 2688
rect 9386 2208 9702 2209
rect 9386 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9702 2208
rect 9386 2143 9702 2144
rect 17827 2208 18143 2209
rect 17827 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18143 2208
rect 17827 2143 18143 2144
rect 26268 2208 26584 2209
rect 26268 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26584 2208
rect 26268 2143 26584 2144
rect 34709 2208 35025 2209
rect 34709 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35025 2208
rect 34709 2143 35025 2144
<< via3 >>
rect 9392 33756 9456 33760
rect 9392 33700 9396 33756
rect 9396 33700 9452 33756
rect 9452 33700 9456 33756
rect 9392 33696 9456 33700
rect 9472 33756 9536 33760
rect 9472 33700 9476 33756
rect 9476 33700 9532 33756
rect 9532 33700 9536 33756
rect 9472 33696 9536 33700
rect 9552 33756 9616 33760
rect 9552 33700 9556 33756
rect 9556 33700 9612 33756
rect 9612 33700 9616 33756
rect 9552 33696 9616 33700
rect 9632 33756 9696 33760
rect 9632 33700 9636 33756
rect 9636 33700 9692 33756
rect 9692 33700 9696 33756
rect 9632 33696 9696 33700
rect 17833 33756 17897 33760
rect 17833 33700 17837 33756
rect 17837 33700 17893 33756
rect 17893 33700 17897 33756
rect 17833 33696 17897 33700
rect 17913 33756 17977 33760
rect 17913 33700 17917 33756
rect 17917 33700 17973 33756
rect 17973 33700 17977 33756
rect 17913 33696 17977 33700
rect 17993 33756 18057 33760
rect 17993 33700 17997 33756
rect 17997 33700 18053 33756
rect 18053 33700 18057 33756
rect 17993 33696 18057 33700
rect 18073 33756 18137 33760
rect 18073 33700 18077 33756
rect 18077 33700 18133 33756
rect 18133 33700 18137 33756
rect 18073 33696 18137 33700
rect 26274 33756 26338 33760
rect 26274 33700 26278 33756
rect 26278 33700 26334 33756
rect 26334 33700 26338 33756
rect 26274 33696 26338 33700
rect 26354 33756 26418 33760
rect 26354 33700 26358 33756
rect 26358 33700 26414 33756
rect 26414 33700 26418 33756
rect 26354 33696 26418 33700
rect 26434 33756 26498 33760
rect 26434 33700 26438 33756
rect 26438 33700 26494 33756
rect 26494 33700 26498 33756
rect 26434 33696 26498 33700
rect 26514 33756 26578 33760
rect 26514 33700 26518 33756
rect 26518 33700 26574 33756
rect 26574 33700 26578 33756
rect 26514 33696 26578 33700
rect 34715 33756 34779 33760
rect 34715 33700 34719 33756
rect 34719 33700 34775 33756
rect 34775 33700 34779 33756
rect 34715 33696 34779 33700
rect 34795 33756 34859 33760
rect 34795 33700 34799 33756
rect 34799 33700 34855 33756
rect 34855 33700 34859 33756
rect 34795 33696 34859 33700
rect 34875 33756 34939 33760
rect 34875 33700 34879 33756
rect 34879 33700 34935 33756
rect 34935 33700 34939 33756
rect 34875 33696 34939 33700
rect 34955 33756 35019 33760
rect 34955 33700 34959 33756
rect 34959 33700 35015 33756
rect 35015 33700 35019 33756
rect 34955 33696 35019 33700
rect 5172 33212 5236 33216
rect 5172 33156 5176 33212
rect 5176 33156 5232 33212
rect 5232 33156 5236 33212
rect 5172 33152 5236 33156
rect 5252 33212 5316 33216
rect 5252 33156 5256 33212
rect 5256 33156 5312 33212
rect 5312 33156 5316 33212
rect 5252 33152 5316 33156
rect 5332 33212 5396 33216
rect 5332 33156 5336 33212
rect 5336 33156 5392 33212
rect 5392 33156 5396 33212
rect 5332 33152 5396 33156
rect 5412 33212 5476 33216
rect 5412 33156 5416 33212
rect 5416 33156 5472 33212
rect 5472 33156 5476 33212
rect 5412 33152 5476 33156
rect 13613 33212 13677 33216
rect 13613 33156 13617 33212
rect 13617 33156 13673 33212
rect 13673 33156 13677 33212
rect 13613 33152 13677 33156
rect 13693 33212 13757 33216
rect 13693 33156 13697 33212
rect 13697 33156 13753 33212
rect 13753 33156 13757 33212
rect 13693 33152 13757 33156
rect 13773 33212 13837 33216
rect 13773 33156 13777 33212
rect 13777 33156 13833 33212
rect 13833 33156 13837 33212
rect 13773 33152 13837 33156
rect 13853 33212 13917 33216
rect 13853 33156 13857 33212
rect 13857 33156 13913 33212
rect 13913 33156 13917 33212
rect 13853 33152 13917 33156
rect 22054 33212 22118 33216
rect 22054 33156 22058 33212
rect 22058 33156 22114 33212
rect 22114 33156 22118 33212
rect 22054 33152 22118 33156
rect 22134 33212 22198 33216
rect 22134 33156 22138 33212
rect 22138 33156 22194 33212
rect 22194 33156 22198 33212
rect 22134 33152 22198 33156
rect 22214 33212 22278 33216
rect 22214 33156 22218 33212
rect 22218 33156 22274 33212
rect 22274 33156 22278 33212
rect 22214 33152 22278 33156
rect 22294 33212 22358 33216
rect 22294 33156 22298 33212
rect 22298 33156 22354 33212
rect 22354 33156 22358 33212
rect 22294 33152 22358 33156
rect 30495 33212 30559 33216
rect 30495 33156 30499 33212
rect 30499 33156 30555 33212
rect 30555 33156 30559 33212
rect 30495 33152 30559 33156
rect 30575 33212 30639 33216
rect 30575 33156 30579 33212
rect 30579 33156 30635 33212
rect 30635 33156 30639 33212
rect 30575 33152 30639 33156
rect 30655 33212 30719 33216
rect 30655 33156 30659 33212
rect 30659 33156 30715 33212
rect 30715 33156 30719 33212
rect 30655 33152 30719 33156
rect 30735 33212 30799 33216
rect 30735 33156 30739 33212
rect 30739 33156 30795 33212
rect 30795 33156 30799 33212
rect 30735 33152 30799 33156
rect 9392 32668 9456 32672
rect 9392 32612 9396 32668
rect 9396 32612 9452 32668
rect 9452 32612 9456 32668
rect 9392 32608 9456 32612
rect 9472 32668 9536 32672
rect 9472 32612 9476 32668
rect 9476 32612 9532 32668
rect 9532 32612 9536 32668
rect 9472 32608 9536 32612
rect 9552 32668 9616 32672
rect 9552 32612 9556 32668
rect 9556 32612 9612 32668
rect 9612 32612 9616 32668
rect 9552 32608 9616 32612
rect 9632 32668 9696 32672
rect 9632 32612 9636 32668
rect 9636 32612 9692 32668
rect 9692 32612 9696 32668
rect 9632 32608 9696 32612
rect 17833 32668 17897 32672
rect 17833 32612 17837 32668
rect 17837 32612 17893 32668
rect 17893 32612 17897 32668
rect 17833 32608 17897 32612
rect 17913 32668 17977 32672
rect 17913 32612 17917 32668
rect 17917 32612 17973 32668
rect 17973 32612 17977 32668
rect 17913 32608 17977 32612
rect 17993 32668 18057 32672
rect 17993 32612 17997 32668
rect 17997 32612 18053 32668
rect 18053 32612 18057 32668
rect 17993 32608 18057 32612
rect 18073 32668 18137 32672
rect 18073 32612 18077 32668
rect 18077 32612 18133 32668
rect 18133 32612 18137 32668
rect 18073 32608 18137 32612
rect 26274 32668 26338 32672
rect 26274 32612 26278 32668
rect 26278 32612 26334 32668
rect 26334 32612 26338 32668
rect 26274 32608 26338 32612
rect 26354 32668 26418 32672
rect 26354 32612 26358 32668
rect 26358 32612 26414 32668
rect 26414 32612 26418 32668
rect 26354 32608 26418 32612
rect 26434 32668 26498 32672
rect 26434 32612 26438 32668
rect 26438 32612 26494 32668
rect 26494 32612 26498 32668
rect 26434 32608 26498 32612
rect 26514 32668 26578 32672
rect 26514 32612 26518 32668
rect 26518 32612 26574 32668
rect 26574 32612 26578 32668
rect 26514 32608 26578 32612
rect 34715 32668 34779 32672
rect 34715 32612 34719 32668
rect 34719 32612 34775 32668
rect 34775 32612 34779 32668
rect 34715 32608 34779 32612
rect 34795 32668 34859 32672
rect 34795 32612 34799 32668
rect 34799 32612 34855 32668
rect 34855 32612 34859 32668
rect 34795 32608 34859 32612
rect 34875 32668 34939 32672
rect 34875 32612 34879 32668
rect 34879 32612 34935 32668
rect 34935 32612 34939 32668
rect 34875 32608 34939 32612
rect 34955 32668 35019 32672
rect 34955 32612 34959 32668
rect 34959 32612 35015 32668
rect 35015 32612 35019 32668
rect 34955 32608 35019 32612
rect 5172 32124 5236 32128
rect 5172 32068 5176 32124
rect 5176 32068 5232 32124
rect 5232 32068 5236 32124
rect 5172 32064 5236 32068
rect 5252 32124 5316 32128
rect 5252 32068 5256 32124
rect 5256 32068 5312 32124
rect 5312 32068 5316 32124
rect 5252 32064 5316 32068
rect 5332 32124 5396 32128
rect 5332 32068 5336 32124
rect 5336 32068 5392 32124
rect 5392 32068 5396 32124
rect 5332 32064 5396 32068
rect 5412 32124 5476 32128
rect 5412 32068 5416 32124
rect 5416 32068 5472 32124
rect 5472 32068 5476 32124
rect 5412 32064 5476 32068
rect 13613 32124 13677 32128
rect 13613 32068 13617 32124
rect 13617 32068 13673 32124
rect 13673 32068 13677 32124
rect 13613 32064 13677 32068
rect 13693 32124 13757 32128
rect 13693 32068 13697 32124
rect 13697 32068 13753 32124
rect 13753 32068 13757 32124
rect 13693 32064 13757 32068
rect 13773 32124 13837 32128
rect 13773 32068 13777 32124
rect 13777 32068 13833 32124
rect 13833 32068 13837 32124
rect 13773 32064 13837 32068
rect 13853 32124 13917 32128
rect 13853 32068 13857 32124
rect 13857 32068 13913 32124
rect 13913 32068 13917 32124
rect 13853 32064 13917 32068
rect 22054 32124 22118 32128
rect 22054 32068 22058 32124
rect 22058 32068 22114 32124
rect 22114 32068 22118 32124
rect 22054 32064 22118 32068
rect 22134 32124 22198 32128
rect 22134 32068 22138 32124
rect 22138 32068 22194 32124
rect 22194 32068 22198 32124
rect 22134 32064 22198 32068
rect 22214 32124 22278 32128
rect 22214 32068 22218 32124
rect 22218 32068 22274 32124
rect 22274 32068 22278 32124
rect 22214 32064 22278 32068
rect 22294 32124 22358 32128
rect 22294 32068 22298 32124
rect 22298 32068 22354 32124
rect 22354 32068 22358 32124
rect 22294 32064 22358 32068
rect 30495 32124 30559 32128
rect 30495 32068 30499 32124
rect 30499 32068 30555 32124
rect 30555 32068 30559 32124
rect 30495 32064 30559 32068
rect 30575 32124 30639 32128
rect 30575 32068 30579 32124
rect 30579 32068 30635 32124
rect 30635 32068 30639 32124
rect 30575 32064 30639 32068
rect 30655 32124 30719 32128
rect 30655 32068 30659 32124
rect 30659 32068 30715 32124
rect 30715 32068 30719 32124
rect 30655 32064 30719 32068
rect 30735 32124 30799 32128
rect 30735 32068 30739 32124
rect 30739 32068 30795 32124
rect 30795 32068 30799 32124
rect 30735 32064 30799 32068
rect 9392 31580 9456 31584
rect 9392 31524 9396 31580
rect 9396 31524 9452 31580
rect 9452 31524 9456 31580
rect 9392 31520 9456 31524
rect 9472 31580 9536 31584
rect 9472 31524 9476 31580
rect 9476 31524 9532 31580
rect 9532 31524 9536 31580
rect 9472 31520 9536 31524
rect 9552 31580 9616 31584
rect 9552 31524 9556 31580
rect 9556 31524 9612 31580
rect 9612 31524 9616 31580
rect 9552 31520 9616 31524
rect 9632 31580 9696 31584
rect 9632 31524 9636 31580
rect 9636 31524 9692 31580
rect 9692 31524 9696 31580
rect 9632 31520 9696 31524
rect 17833 31580 17897 31584
rect 17833 31524 17837 31580
rect 17837 31524 17893 31580
rect 17893 31524 17897 31580
rect 17833 31520 17897 31524
rect 17913 31580 17977 31584
rect 17913 31524 17917 31580
rect 17917 31524 17973 31580
rect 17973 31524 17977 31580
rect 17913 31520 17977 31524
rect 17993 31580 18057 31584
rect 17993 31524 17997 31580
rect 17997 31524 18053 31580
rect 18053 31524 18057 31580
rect 17993 31520 18057 31524
rect 18073 31580 18137 31584
rect 18073 31524 18077 31580
rect 18077 31524 18133 31580
rect 18133 31524 18137 31580
rect 18073 31520 18137 31524
rect 26274 31580 26338 31584
rect 26274 31524 26278 31580
rect 26278 31524 26334 31580
rect 26334 31524 26338 31580
rect 26274 31520 26338 31524
rect 26354 31580 26418 31584
rect 26354 31524 26358 31580
rect 26358 31524 26414 31580
rect 26414 31524 26418 31580
rect 26354 31520 26418 31524
rect 26434 31580 26498 31584
rect 26434 31524 26438 31580
rect 26438 31524 26494 31580
rect 26494 31524 26498 31580
rect 26434 31520 26498 31524
rect 26514 31580 26578 31584
rect 26514 31524 26518 31580
rect 26518 31524 26574 31580
rect 26574 31524 26578 31580
rect 26514 31520 26578 31524
rect 34715 31580 34779 31584
rect 34715 31524 34719 31580
rect 34719 31524 34775 31580
rect 34775 31524 34779 31580
rect 34715 31520 34779 31524
rect 34795 31580 34859 31584
rect 34795 31524 34799 31580
rect 34799 31524 34855 31580
rect 34855 31524 34859 31580
rect 34795 31520 34859 31524
rect 34875 31580 34939 31584
rect 34875 31524 34879 31580
rect 34879 31524 34935 31580
rect 34935 31524 34939 31580
rect 34875 31520 34939 31524
rect 34955 31580 35019 31584
rect 34955 31524 34959 31580
rect 34959 31524 35015 31580
rect 35015 31524 35019 31580
rect 34955 31520 35019 31524
rect 5172 31036 5236 31040
rect 5172 30980 5176 31036
rect 5176 30980 5232 31036
rect 5232 30980 5236 31036
rect 5172 30976 5236 30980
rect 5252 31036 5316 31040
rect 5252 30980 5256 31036
rect 5256 30980 5312 31036
rect 5312 30980 5316 31036
rect 5252 30976 5316 30980
rect 5332 31036 5396 31040
rect 5332 30980 5336 31036
rect 5336 30980 5392 31036
rect 5392 30980 5396 31036
rect 5332 30976 5396 30980
rect 5412 31036 5476 31040
rect 5412 30980 5416 31036
rect 5416 30980 5472 31036
rect 5472 30980 5476 31036
rect 5412 30976 5476 30980
rect 13613 31036 13677 31040
rect 13613 30980 13617 31036
rect 13617 30980 13673 31036
rect 13673 30980 13677 31036
rect 13613 30976 13677 30980
rect 13693 31036 13757 31040
rect 13693 30980 13697 31036
rect 13697 30980 13753 31036
rect 13753 30980 13757 31036
rect 13693 30976 13757 30980
rect 13773 31036 13837 31040
rect 13773 30980 13777 31036
rect 13777 30980 13833 31036
rect 13833 30980 13837 31036
rect 13773 30976 13837 30980
rect 13853 31036 13917 31040
rect 13853 30980 13857 31036
rect 13857 30980 13913 31036
rect 13913 30980 13917 31036
rect 13853 30976 13917 30980
rect 22054 31036 22118 31040
rect 22054 30980 22058 31036
rect 22058 30980 22114 31036
rect 22114 30980 22118 31036
rect 22054 30976 22118 30980
rect 22134 31036 22198 31040
rect 22134 30980 22138 31036
rect 22138 30980 22194 31036
rect 22194 30980 22198 31036
rect 22134 30976 22198 30980
rect 22214 31036 22278 31040
rect 22214 30980 22218 31036
rect 22218 30980 22274 31036
rect 22274 30980 22278 31036
rect 22214 30976 22278 30980
rect 22294 31036 22358 31040
rect 22294 30980 22298 31036
rect 22298 30980 22354 31036
rect 22354 30980 22358 31036
rect 22294 30976 22358 30980
rect 30495 31036 30559 31040
rect 30495 30980 30499 31036
rect 30499 30980 30555 31036
rect 30555 30980 30559 31036
rect 30495 30976 30559 30980
rect 30575 31036 30639 31040
rect 30575 30980 30579 31036
rect 30579 30980 30635 31036
rect 30635 30980 30639 31036
rect 30575 30976 30639 30980
rect 30655 31036 30719 31040
rect 30655 30980 30659 31036
rect 30659 30980 30715 31036
rect 30715 30980 30719 31036
rect 30655 30976 30719 30980
rect 30735 31036 30799 31040
rect 30735 30980 30739 31036
rect 30739 30980 30795 31036
rect 30795 30980 30799 31036
rect 30735 30976 30799 30980
rect 9392 30492 9456 30496
rect 9392 30436 9396 30492
rect 9396 30436 9452 30492
rect 9452 30436 9456 30492
rect 9392 30432 9456 30436
rect 9472 30492 9536 30496
rect 9472 30436 9476 30492
rect 9476 30436 9532 30492
rect 9532 30436 9536 30492
rect 9472 30432 9536 30436
rect 9552 30492 9616 30496
rect 9552 30436 9556 30492
rect 9556 30436 9612 30492
rect 9612 30436 9616 30492
rect 9552 30432 9616 30436
rect 9632 30492 9696 30496
rect 9632 30436 9636 30492
rect 9636 30436 9692 30492
rect 9692 30436 9696 30492
rect 9632 30432 9696 30436
rect 17833 30492 17897 30496
rect 17833 30436 17837 30492
rect 17837 30436 17893 30492
rect 17893 30436 17897 30492
rect 17833 30432 17897 30436
rect 17913 30492 17977 30496
rect 17913 30436 17917 30492
rect 17917 30436 17973 30492
rect 17973 30436 17977 30492
rect 17913 30432 17977 30436
rect 17993 30492 18057 30496
rect 17993 30436 17997 30492
rect 17997 30436 18053 30492
rect 18053 30436 18057 30492
rect 17993 30432 18057 30436
rect 18073 30492 18137 30496
rect 18073 30436 18077 30492
rect 18077 30436 18133 30492
rect 18133 30436 18137 30492
rect 18073 30432 18137 30436
rect 26274 30492 26338 30496
rect 26274 30436 26278 30492
rect 26278 30436 26334 30492
rect 26334 30436 26338 30492
rect 26274 30432 26338 30436
rect 26354 30492 26418 30496
rect 26354 30436 26358 30492
rect 26358 30436 26414 30492
rect 26414 30436 26418 30492
rect 26354 30432 26418 30436
rect 26434 30492 26498 30496
rect 26434 30436 26438 30492
rect 26438 30436 26494 30492
rect 26494 30436 26498 30492
rect 26434 30432 26498 30436
rect 26514 30492 26578 30496
rect 26514 30436 26518 30492
rect 26518 30436 26574 30492
rect 26574 30436 26578 30492
rect 26514 30432 26578 30436
rect 34715 30492 34779 30496
rect 34715 30436 34719 30492
rect 34719 30436 34775 30492
rect 34775 30436 34779 30492
rect 34715 30432 34779 30436
rect 34795 30492 34859 30496
rect 34795 30436 34799 30492
rect 34799 30436 34855 30492
rect 34855 30436 34859 30492
rect 34795 30432 34859 30436
rect 34875 30492 34939 30496
rect 34875 30436 34879 30492
rect 34879 30436 34935 30492
rect 34935 30436 34939 30492
rect 34875 30432 34939 30436
rect 34955 30492 35019 30496
rect 34955 30436 34959 30492
rect 34959 30436 35015 30492
rect 35015 30436 35019 30492
rect 34955 30432 35019 30436
rect 5172 29948 5236 29952
rect 5172 29892 5176 29948
rect 5176 29892 5232 29948
rect 5232 29892 5236 29948
rect 5172 29888 5236 29892
rect 5252 29948 5316 29952
rect 5252 29892 5256 29948
rect 5256 29892 5312 29948
rect 5312 29892 5316 29948
rect 5252 29888 5316 29892
rect 5332 29948 5396 29952
rect 5332 29892 5336 29948
rect 5336 29892 5392 29948
rect 5392 29892 5396 29948
rect 5332 29888 5396 29892
rect 5412 29948 5476 29952
rect 5412 29892 5416 29948
rect 5416 29892 5472 29948
rect 5472 29892 5476 29948
rect 5412 29888 5476 29892
rect 13613 29948 13677 29952
rect 13613 29892 13617 29948
rect 13617 29892 13673 29948
rect 13673 29892 13677 29948
rect 13613 29888 13677 29892
rect 13693 29948 13757 29952
rect 13693 29892 13697 29948
rect 13697 29892 13753 29948
rect 13753 29892 13757 29948
rect 13693 29888 13757 29892
rect 13773 29948 13837 29952
rect 13773 29892 13777 29948
rect 13777 29892 13833 29948
rect 13833 29892 13837 29948
rect 13773 29888 13837 29892
rect 13853 29948 13917 29952
rect 13853 29892 13857 29948
rect 13857 29892 13913 29948
rect 13913 29892 13917 29948
rect 13853 29888 13917 29892
rect 22054 29948 22118 29952
rect 22054 29892 22058 29948
rect 22058 29892 22114 29948
rect 22114 29892 22118 29948
rect 22054 29888 22118 29892
rect 22134 29948 22198 29952
rect 22134 29892 22138 29948
rect 22138 29892 22194 29948
rect 22194 29892 22198 29948
rect 22134 29888 22198 29892
rect 22214 29948 22278 29952
rect 22214 29892 22218 29948
rect 22218 29892 22274 29948
rect 22274 29892 22278 29948
rect 22214 29888 22278 29892
rect 22294 29948 22358 29952
rect 22294 29892 22298 29948
rect 22298 29892 22354 29948
rect 22354 29892 22358 29948
rect 22294 29888 22358 29892
rect 30495 29948 30559 29952
rect 30495 29892 30499 29948
rect 30499 29892 30555 29948
rect 30555 29892 30559 29948
rect 30495 29888 30559 29892
rect 30575 29948 30639 29952
rect 30575 29892 30579 29948
rect 30579 29892 30635 29948
rect 30635 29892 30639 29948
rect 30575 29888 30639 29892
rect 30655 29948 30719 29952
rect 30655 29892 30659 29948
rect 30659 29892 30715 29948
rect 30715 29892 30719 29948
rect 30655 29888 30719 29892
rect 30735 29948 30799 29952
rect 30735 29892 30739 29948
rect 30739 29892 30795 29948
rect 30795 29892 30799 29948
rect 30735 29888 30799 29892
rect 9392 29404 9456 29408
rect 9392 29348 9396 29404
rect 9396 29348 9452 29404
rect 9452 29348 9456 29404
rect 9392 29344 9456 29348
rect 9472 29404 9536 29408
rect 9472 29348 9476 29404
rect 9476 29348 9532 29404
rect 9532 29348 9536 29404
rect 9472 29344 9536 29348
rect 9552 29404 9616 29408
rect 9552 29348 9556 29404
rect 9556 29348 9612 29404
rect 9612 29348 9616 29404
rect 9552 29344 9616 29348
rect 9632 29404 9696 29408
rect 9632 29348 9636 29404
rect 9636 29348 9692 29404
rect 9692 29348 9696 29404
rect 9632 29344 9696 29348
rect 17833 29404 17897 29408
rect 17833 29348 17837 29404
rect 17837 29348 17893 29404
rect 17893 29348 17897 29404
rect 17833 29344 17897 29348
rect 17913 29404 17977 29408
rect 17913 29348 17917 29404
rect 17917 29348 17973 29404
rect 17973 29348 17977 29404
rect 17913 29344 17977 29348
rect 17993 29404 18057 29408
rect 17993 29348 17997 29404
rect 17997 29348 18053 29404
rect 18053 29348 18057 29404
rect 17993 29344 18057 29348
rect 18073 29404 18137 29408
rect 18073 29348 18077 29404
rect 18077 29348 18133 29404
rect 18133 29348 18137 29404
rect 18073 29344 18137 29348
rect 26274 29404 26338 29408
rect 26274 29348 26278 29404
rect 26278 29348 26334 29404
rect 26334 29348 26338 29404
rect 26274 29344 26338 29348
rect 26354 29404 26418 29408
rect 26354 29348 26358 29404
rect 26358 29348 26414 29404
rect 26414 29348 26418 29404
rect 26354 29344 26418 29348
rect 26434 29404 26498 29408
rect 26434 29348 26438 29404
rect 26438 29348 26494 29404
rect 26494 29348 26498 29404
rect 26434 29344 26498 29348
rect 26514 29404 26578 29408
rect 26514 29348 26518 29404
rect 26518 29348 26574 29404
rect 26574 29348 26578 29404
rect 26514 29344 26578 29348
rect 34715 29404 34779 29408
rect 34715 29348 34719 29404
rect 34719 29348 34775 29404
rect 34775 29348 34779 29404
rect 34715 29344 34779 29348
rect 34795 29404 34859 29408
rect 34795 29348 34799 29404
rect 34799 29348 34855 29404
rect 34855 29348 34859 29404
rect 34795 29344 34859 29348
rect 34875 29404 34939 29408
rect 34875 29348 34879 29404
rect 34879 29348 34935 29404
rect 34935 29348 34939 29404
rect 34875 29344 34939 29348
rect 34955 29404 35019 29408
rect 34955 29348 34959 29404
rect 34959 29348 35015 29404
rect 35015 29348 35019 29404
rect 34955 29344 35019 29348
rect 5172 28860 5236 28864
rect 5172 28804 5176 28860
rect 5176 28804 5232 28860
rect 5232 28804 5236 28860
rect 5172 28800 5236 28804
rect 5252 28860 5316 28864
rect 5252 28804 5256 28860
rect 5256 28804 5312 28860
rect 5312 28804 5316 28860
rect 5252 28800 5316 28804
rect 5332 28860 5396 28864
rect 5332 28804 5336 28860
rect 5336 28804 5392 28860
rect 5392 28804 5396 28860
rect 5332 28800 5396 28804
rect 5412 28860 5476 28864
rect 5412 28804 5416 28860
rect 5416 28804 5472 28860
rect 5472 28804 5476 28860
rect 5412 28800 5476 28804
rect 13613 28860 13677 28864
rect 13613 28804 13617 28860
rect 13617 28804 13673 28860
rect 13673 28804 13677 28860
rect 13613 28800 13677 28804
rect 13693 28860 13757 28864
rect 13693 28804 13697 28860
rect 13697 28804 13753 28860
rect 13753 28804 13757 28860
rect 13693 28800 13757 28804
rect 13773 28860 13837 28864
rect 13773 28804 13777 28860
rect 13777 28804 13833 28860
rect 13833 28804 13837 28860
rect 13773 28800 13837 28804
rect 13853 28860 13917 28864
rect 13853 28804 13857 28860
rect 13857 28804 13913 28860
rect 13913 28804 13917 28860
rect 13853 28800 13917 28804
rect 22054 28860 22118 28864
rect 22054 28804 22058 28860
rect 22058 28804 22114 28860
rect 22114 28804 22118 28860
rect 22054 28800 22118 28804
rect 22134 28860 22198 28864
rect 22134 28804 22138 28860
rect 22138 28804 22194 28860
rect 22194 28804 22198 28860
rect 22134 28800 22198 28804
rect 22214 28860 22278 28864
rect 22214 28804 22218 28860
rect 22218 28804 22274 28860
rect 22274 28804 22278 28860
rect 22214 28800 22278 28804
rect 22294 28860 22358 28864
rect 22294 28804 22298 28860
rect 22298 28804 22354 28860
rect 22354 28804 22358 28860
rect 22294 28800 22358 28804
rect 30495 28860 30559 28864
rect 30495 28804 30499 28860
rect 30499 28804 30555 28860
rect 30555 28804 30559 28860
rect 30495 28800 30559 28804
rect 30575 28860 30639 28864
rect 30575 28804 30579 28860
rect 30579 28804 30635 28860
rect 30635 28804 30639 28860
rect 30575 28800 30639 28804
rect 30655 28860 30719 28864
rect 30655 28804 30659 28860
rect 30659 28804 30715 28860
rect 30715 28804 30719 28860
rect 30655 28800 30719 28804
rect 30735 28860 30799 28864
rect 30735 28804 30739 28860
rect 30739 28804 30795 28860
rect 30795 28804 30799 28860
rect 30735 28800 30799 28804
rect 9392 28316 9456 28320
rect 9392 28260 9396 28316
rect 9396 28260 9452 28316
rect 9452 28260 9456 28316
rect 9392 28256 9456 28260
rect 9472 28316 9536 28320
rect 9472 28260 9476 28316
rect 9476 28260 9532 28316
rect 9532 28260 9536 28316
rect 9472 28256 9536 28260
rect 9552 28316 9616 28320
rect 9552 28260 9556 28316
rect 9556 28260 9612 28316
rect 9612 28260 9616 28316
rect 9552 28256 9616 28260
rect 9632 28316 9696 28320
rect 9632 28260 9636 28316
rect 9636 28260 9692 28316
rect 9692 28260 9696 28316
rect 9632 28256 9696 28260
rect 17833 28316 17897 28320
rect 17833 28260 17837 28316
rect 17837 28260 17893 28316
rect 17893 28260 17897 28316
rect 17833 28256 17897 28260
rect 17913 28316 17977 28320
rect 17913 28260 17917 28316
rect 17917 28260 17973 28316
rect 17973 28260 17977 28316
rect 17913 28256 17977 28260
rect 17993 28316 18057 28320
rect 17993 28260 17997 28316
rect 17997 28260 18053 28316
rect 18053 28260 18057 28316
rect 17993 28256 18057 28260
rect 18073 28316 18137 28320
rect 18073 28260 18077 28316
rect 18077 28260 18133 28316
rect 18133 28260 18137 28316
rect 18073 28256 18137 28260
rect 26274 28316 26338 28320
rect 26274 28260 26278 28316
rect 26278 28260 26334 28316
rect 26334 28260 26338 28316
rect 26274 28256 26338 28260
rect 26354 28316 26418 28320
rect 26354 28260 26358 28316
rect 26358 28260 26414 28316
rect 26414 28260 26418 28316
rect 26354 28256 26418 28260
rect 26434 28316 26498 28320
rect 26434 28260 26438 28316
rect 26438 28260 26494 28316
rect 26494 28260 26498 28316
rect 26434 28256 26498 28260
rect 26514 28316 26578 28320
rect 26514 28260 26518 28316
rect 26518 28260 26574 28316
rect 26574 28260 26578 28316
rect 26514 28256 26578 28260
rect 34715 28316 34779 28320
rect 34715 28260 34719 28316
rect 34719 28260 34775 28316
rect 34775 28260 34779 28316
rect 34715 28256 34779 28260
rect 34795 28316 34859 28320
rect 34795 28260 34799 28316
rect 34799 28260 34855 28316
rect 34855 28260 34859 28316
rect 34795 28256 34859 28260
rect 34875 28316 34939 28320
rect 34875 28260 34879 28316
rect 34879 28260 34935 28316
rect 34935 28260 34939 28316
rect 34875 28256 34939 28260
rect 34955 28316 35019 28320
rect 34955 28260 34959 28316
rect 34959 28260 35015 28316
rect 35015 28260 35019 28316
rect 34955 28256 35019 28260
rect 5172 27772 5236 27776
rect 5172 27716 5176 27772
rect 5176 27716 5232 27772
rect 5232 27716 5236 27772
rect 5172 27712 5236 27716
rect 5252 27772 5316 27776
rect 5252 27716 5256 27772
rect 5256 27716 5312 27772
rect 5312 27716 5316 27772
rect 5252 27712 5316 27716
rect 5332 27772 5396 27776
rect 5332 27716 5336 27772
rect 5336 27716 5392 27772
rect 5392 27716 5396 27772
rect 5332 27712 5396 27716
rect 5412 27772 5476 27776
rect 5412 27716 5416 27772
rect 5416 27716 5472 27772
rect 5472 27716 5476 27772
rect 5412 27712 5476 27716
rect 13613 27772 13677 27776
rect 13613 27716 13617 27772
rect 13617 27716 13673 27772
rect 13673 27716 13677 27772
rect 13613 27712 13677 27716
rect 13693 27772 13757 27776
rect 13693 27716 13697 27772
rect 13697 27716 13753 27772
rect 13753 27716 13757 27772
rect 13693 27712 13757 27716
rect 13773 27772 13837 27776
rect 13773 27716 13777 27772
rect 13777 27716 13833 27772
rect 13833 27716 13837 27772
rect 13773 27712 13837 27716
rect 13853 27772 13917 27776
rect 13853 27716 13857 27772
rect 13857 27716 13913 27772
rect 13913 27716 13917 27772
rect 13853 27712 13917 27716
rect 22054 27772 22118 27776
rect 22054 27716 22058 27772
rect 22058 27716 22114 27772
rect 22114 27716 22118 27772
rect 22054 27712 22118 27716
rect 22134 27772 22198 27776
rect 22134 27716 22138 27772
rect 22138 27716 22194 27772
rect 22194 27716 22198 27772
rect 22134 27712 22198 27716
rect 22214 27772 22278 27776
rect 22214 27716 22218 27772
rect 22218 27716 22274 27772
rect 22274 27716 22278 27772
rect 22214 27712 22278 27716
rect 22294 27772 22358 27776
rect 22294 27716 22298 27772
rect 22298 27716 22354 27772
rect 22354 27716 22358 27772
rect 22294 27712 22358 27716
rect 30495 27772 30559 27776
rect 30495 27716 30499 27772
rect 30499 27716 30555 27772
rect 30555 27716 30559 27772
rect 30495 27712 30559 27716
rect 30575 27772 30639 27776
rect 30575 27716 30579 27772
rect 30579 27716 30635 27772
rect 30635 27716 30639 27772
rect 30575 27712 30639 27716
rect 30655 27772 30719 27776
rect 30655 27716 30659 27772
rect 30659 27716 30715 27772
rect 30715 27716 30719 27772
rect 30655 27712 30719 27716
rect 30735 27772 30799 27776
rect 30735 27716 30739 27772
rect 30739 27716 30795 27772
rect 30795 27716 30799 27772
rect 30735 27712 30799 27716
rect 9392 27228 9456 27232
rect 9392 27172 9396 27228
rect 9396 27172 9452 27228
rect 9452 27172 9456 27228
rect 9392 27168 9456 27172
rect 9472 27228 9536 27232
rect 9472 27172 9476 27228
rect 9476 27172 9532 27228
rect 9532 27172 9536 27228
rect 9472 27168 9536 27172
rect 9552 27228 9616 27232
rect 9552 27172 9556 27228
rect 9556 27172 9612 27228
rect 9612 27172 9616 27228
rect 9552 27168 9616 27172
rect 9632 27228 9696 27232
rect 9632 27172 9636 27228
rect 9636 27172 9692 27228
rect 9692 27172 9696 27228
rect 9632 27168 9696 27172
rect 17833 27228 17897 27232
rect 17833 27172 17837 27228
rect 17837 27172 17893 27228
rect 17893 27172 17897 27228
rect 17833 27168 17897 27172
rect 17913 27228 17977 27232
rect 17913 27172 17917 27228
rect 17917 27172 17973 27228
rect 17973 27172 17977 27228
rect 17913 27168 17977 27172
rect 17993 27228 18057 27232
rect 17993 27172 17997 27228
rect 17997 27172 18053 27228
rect 18053 27172 18057 27228
rect 17993 27168 18057 27172
rect 18073 27228 18137 27232
rect 18073 27172 18077 27228
rect 18077 27172 18133 27228
rect 18133 27172 18137 27228
rect 18073 27168 18137 27172
rect 26274 27228 26338 27232
rect 26274 27172 26278 27228
rect 26278 27172 26334 27228
rect 26334 27172 26338 27228
rect 26274 27168 26338 27172
rect 26354 27228 26418 27232
rect 26354 27172 26358 27228
rect 26358 27172 26414 27228
rect 26414 27172 26418 27228
rect 26354 27168 26418 27172
rect 26434 27228 26498 27232
rect 26434 27172 26438 27228
rect 26438 27172 26494 27228
rect 26494 27172 26498 27228
rect 26434 27168 26498 27172
rect 26514 27228 26578 27232
rect 26514 27172 26518 27228
rect 26518 27172 26574 27228
rect 26574 27172 26578 27228
rect 26514 27168 26578 27172
rect 34715 27228 34779 27232
rect 34715 27172 34719 27228
rect 34719 27172 34775 27228
rect 34775 27172 34779 27228
rect 34715 27168 34779 27172
rect 34795 27228 34859 27232
rect 34795 27172 34799 27228
rect 34799 27172 34855 27228
rect 34855 27172 34859 27228
rect 34795 27168 34859 27172
rect 34875 27228 34939 27232
rect 34875 27172 34879 27228
rect 34879 27172 34935 27228
rect 34935 27172 34939 27228
rect 34875 27168 34939 27172
rect 34955 27228 35019 27232
rect 34955 27172 34959 27228
rect 34959 27172 35015 27228
rect 35015 27172 35019 27228
rect 34955 27168 35019 27172
rect 5172 26684 5236 26688
rect 5172 26628 5176 26684
rect 5176 26628 5232 26684
rect 5232 26628 5236 26684
rect 5172 26624 5236 26628
rect 5252 26684 5316 26688
rect 5252 26628 5256 26684
rect 5256 26628 5312 26684
rect 5312 26628 5316 26684
rect 5252 26624 5316 26628
rect 5332 26684 5396 26688
rect 5332 26628 5336 26684
rect 5336 26628 5392 26684
rect 5392 26628 5396 26684
rect 5332 26624 5396 26628
rect 5412 26684 5476 26688
rect 5412 26628 5416 26684
rect 5416 26628 5472 26684
rect 5472 26628 5476 26684
rect 5412 26624 5476 26628
rect 13613 26684 13677 26688
rect 13613 26628 13617 26684
rect 13617 26628 13673 26684
rect 13673 26628 13677 26684
rect 13613 26624 13677 26628
rect 13693 26684 13757 26688
rect 13693 26628 13697 26684
rect 13697 26628 13753 26684
rect 13753 26628 13757 26684
rect 13693 26624 13757 26628
rect 13773 26684 13837 26688
rect 13773 26628 13777 26684
rect 13777 26628 13833 26684
rect 13833 26628 13837 26684
rect 13773 26624 13837 26628
rect 13853 26684 13917 26688
rect 13853 26628 13857 26684
rect 13857 26628 13913 26684
rect 13913 26628 13917 26684
rect 13853 26624 13917 26628
rect 22054 26684 22118 26688
rect 22054 26628 22058 26684
rect 22058 26628 22114 26684
rect 22114 26628 22118 26684
rect 22054 26624 22118 26628
rect 22134 26684 22198 26688
rect 22134 26628 22138 26684
rect 22138 26628 22194 26684
rect 22194 26628 22198 26684
rect 22134 26624 22198 26628
rect 22214 26684 22278 26688
rect 22214 26628 22218 26684
rect 22218 26628 22274 26684
rect 22274 26628 22278 26684
rect 22214 26624 22278 26628
rect 22294 26684 22358 26688
rect 22294 26628 22298 26684
rect 22298 26628 22354 26684
rect 22354 26628 22358 26684
rect 22294 26624 22358 26628
rect 30495 26684 30559 26688
rect 30495 26628 30499 26684
rect 30499 26628 30555 26684
rect 30555 26628 30559 26684
rect 30495 26624 30559 26628
rect 30575 26684 30639 26688
rect 30575 26628 30579 26684
rect 30579 26628 30635 26684
rect 30635 26628 30639 26684
rect 30575 26624 30639 26628
rect 30655 26684 30719 26688
rect 30655 26628 30659 26684
rect 30659 26628 30715 26684
rect 30715 26628 30719 26684
rect 30655 26624 30719 26628
rect 30735 26684 30799 26688
rect 30735 26628 30739 26684
rect 30739 26628 30795 26684
rect 30795 26628 30799 26684
rect 30735 26624 30799 26628
rect 9392 26140 9456 26144
rect 9392 26084 9396 26140
rect 9396 26084 9452 26140
rect 9452 26084 9456 26140
rect 9392 26080 9456 26084
rect 9472 26140 9536 26144
rect 9472 26084 9476 26140
rect 9476 26084 9532 26140
rect 9532 26084 9536 26140
rect 9472 26080 9536 26084
rect 9552 26140 9616 26144
rect 9552 26084 9556 26140
rect 9556 26084 9612 26140
rect 9612 26084 9616 26140
rect 9552 26080 9616 26084
rect 9632 26140 9696 26144
rect 9632 26084 9636 26140
rect 9636 26084 9692 26140
rect 9692 26084 9696 26140
rect 9632 26080 9696 26084
rect 17833 26140 17897 26144
rect 17833 26084 17837 26140
rect 17837 26084 17893 26140
rect 17893 26084 17897 26140
rect 17833 26080 17897 26084
rect 17913 26140 17977 26144
rect 17913 26084 17917 26140
rect 17917 26084 17973 26140
rect 17973 26084 17977 26140
rect 17913 26080 17977 26084
rect 17993 26140 18057 26144
rect 17993 26084 17997 26140
rect 17997 26084 18053 26140
rect 18053 26084 18057 26140
rect 17993 26080 18057 26084
rect 18073 26140 18137 26144
rect 18073 26084 18077 26140
rect 18077 26084 18133 26140
rect 18133 26084 18137 26140
rect 18073 26080 18137 26084
rect 26274 26140 26338 26144
rect 26274 26084 26278 26140
rect 26278 26084 26334 26140
rect 26334 26084 26338 26140
rect 26274 26080 26338 26084
rect 26354 26140 26418 26144
rect 26354 26084 26358 26140
rect 26358 26084 26414 26140
rect 26414 26084 26418 26140
rect 26354 26080 26418 26084
rect 26434 26140 26498 26144
rect 26434 26084 26438 26140
rect 26438 26084 26494 26140
rect 26494 26084 26498 26140
rect 26434 26080 26498 26084
rect 26514 26140 26578 26144
rect 26514 26084 26518 26140
rect 26518 26084 26574 26140
rect 26574 26084 26578 26140
rect 26514 26080 26578 26084
rect 34715 26140 34779 26144
rect 34715 26084 34719 26140
rect 34719 26084 34775 26140
rect 34775 26084 34779 26140
rect 34715 26080 34779 26084
rect 34795 26140 34859 26144
rect 34795 26084 34799 26140
rect 34799 26084 34855 26140
rect 34855 26084 34859 26140
rect 34795 26080 34859 26084
rect 34875 26140 34939 26144
rect 34875 26084 34879 26140
rect 34879 26084 34935 26140
rect 34935 26084 34939 26140
rect 34875 26080 34939 26084
rect 34955 26140 35019 26144
rect 34955 26084 34959 26140
rect 34959 26084 35015 26140
rect 35015 26084 35019 26140
rect 34955 26080 35019 26084
rect 5172 25596 5236 25600
rect 5172 25540 5176 25596
rect 5176 25540 5232 25596
rect 5232 25540 5236 25596
rect 5172 25536 5236 25540
rect 5252 25596 5316 25600
rect 5252 25540 5256 25596
rect 5256 25540 5312 25596
rect 5312 25540 5316 25596
rect 5252 25536 5316 25540
rect 5332 25596 5396 25600
rect 5332 25540 5336 25596
rect 5336 25540 5392 25596
rect 5392 25540 5396 25596
rect 5332 25536 5396 25540
rect 5412 25596 5476 25600
rect 5412 25540 5416 25596
rect 5416 25540 5472 25596
rect 5472 25540 5476 25596
rect 5412 25536 5476 25540
rect 13613 25596 13677 25600
rect 13613 25540 13617 25596
rect 13617 25540 13673 25596
rect 13673 25540 13677 25596
rect 13613 25536 13677 25540
rect 13693 25596 13757 25600
rect 13693 25540 13697 25596
rect 13697 25540 13753 25596
rect 13753 25540 13757 25596
rect 13693 25536 13757 25540
rect 13773 25596 13837 25600
rect 13773 25540 13777 25596
rect 13777 25540 13833 25596
rect 13833 25540 13837 25596
rect 13773 25536 13837 25540
rect 13853 25596 13917 25600
rect 13853 25540 13857 25596
rect 13857 25540 13913 25596
rect 13913 25540 13917 25596
rect 13853 25536 13917 25540
rect 22054 25596 22118 25600
rect 22054 25540 22058 25596
rect 22058 25540 22114 25596
rect 22114 25540 22118 25596
rect 22054 25536 22118 25540
rect 22134 25596 22198 25600
rect 22134 25540 22138 25596
rect 22138 25540 22194 25596
rect 22194 25540 22198 25596
rect 22134 25536 22198 25540
rect 22214 25596 22278 25600
rect 22214 25540 22218 25596
rect 22218 25540 22274 25596
rect 22274 25540 22278 25596
rect 22214 25536 22278 25540
rect 22294 25596 22358 25600
rect 22294 25540 22298 25596
rect 22298 25540 22354 25596
rect 22354 25540 22358 25596
rect 22294 25536 22358 25540
rect 30495 25596 30559 25600
rect 30495 25540 30499 25596
rect 30499 25540 30555 25596
rect 30555 25540 30559 25596
rect 30495 25536 30559 25540
rect 30575 25596 30639 25600
rect 30575 25540 30579 25596
rect 30579 25540 30635 25596
rect 30635 25540 30639 25596
rect 30575 25536 30639 25540
rect 30655 25596 30719 25600
rect 30655 25540 30659 25596
rect 30659 25540 30715 25596
rect 30715 25540 30719 25596
rect 30655 25536 30719 25540
rect 30735 25596 30799 25600
rect 30735 25540 30739 25596
rect 30739 25540 30795 25596
rect 30795 25540 30799 25596
rect 30735 25536 30799 25540
rect 9392 25052 9456 25056
rect 9392 24996 9396 25052
rect 9396 24996 9452 25052
rect 9452 24996 9456 25052
rect 9392 24992 9456 24996
rect 9472 25052 9536 25056
rect 9472 24996 9476 25052
rect 9476 24996 9532 25052
rect 9532 24996 9536 25052
rect 9472 24992 9536 24996
rect 9552 25052 9616 25056
rect 9552 24996 9556 25052
rect 9556 24996 9612 25052
rect 9612 24996 9616 25052
rect 9552 24992 9616 24996
rect 9632 25052 9696 25056
rect 9632 24996 9636 25052
rect 9636 24996 9692 25052
rect 9692 24996 9696 25052
rect 9632 24992 9696 24996
rect 17833 25052 17897 25056
rect 17833 24996 17837 25052
rect 17837 24996 17893 25052
rect 17893 24996 17897 25052
rect 17833 24992 17897 24996
rect 17913 25052 17977 25056
rect 17913 24996 17917 25052
rect 17917 24996 17973 25052
rect 17973 24996 17977 25052
rect 17913 24992 17977 24996
rect 17993 25052 18057 25056
rect 17993 24996 17997 25052
rect 17997 24996 18053 25052
rect 18053 24996 18057 25052
rect 17993 24992 18057 24996
rect 18073 25052 18137 25056
rect 18073 24996 18077 25052
rect 18077 24996 18133 25052
rect 18133 24996 18137 25052
rect 18073 24992 18137 24996
rect 26274 25052 26338 25056
rect 26274 24996 26278 25052
rect 26278 24996 26334 25052
rect 26334 24996 26338 25052
rect 26274 24992 26338 24996
rect 26354 25052 26418 25056
rect 26354 24996 26358 25052
rect 26358 24996 26414 25052
rect 26414 24996 26418 25052
rect 26354 24992 26418 24996
rect 26434 25052 26498 25056
rect 26434 24996 26438 25052
rect 26438 24996 26494 25052
rect 26494 24996 26498 25052
rect 26434 24992 26498 24996
rect 26514 25052 26578 25056
rect 26514 24996 26518 25052
rect 26518 24996 26574 25052
rect 26574 24996 26578 25052
rect 26514 24992 26578 24996
rect 34715 25052 34779 25056
rect 34715 24996 34719 25052
rect 34719 24996 34775 25052
rect 34775 24996 34779 25052
rect 34715 24992 34779 24996
rect 34795 25052 34859 25056
rect 34795 24996 34799 25052
rect 34799 24996 34855 25052
rect 34855 24996 34859 25052
rect 34795 24992 34859 24996
rect 34875 25052 34939 25056
rect 34875 24996 34879 25052
rect 34879 24996 34935 25052
rect 34935 24996 34939 25052
rect 34875 24992 34939 24996
rect 34955 25052 35019 25056
rect 34955 24996 34959 25052
rect 34959 24996 35015 25052
rect 35015 24996 35019 25052
rect 34955 24992 35019 24996
rect 5172 24508 5236 24512
rect 5172 24452 5176 24508
rect 5176 24452 5232 24508
rect 5232 24452 5236 24508
rect 5172 24448 5236 24452
rect 5252 24508 5316 24512
rect 5252 24452 5256 24508
rect 5256 24452 5312 24508
rect 5312 24452 5316 24508
rect 5252 24448 5316 24452
rect 5332 24508 5396 24512
rect 5332 24452 5336 24508
rect 5336 24452 5392 24508
rect 5392 24452 5396 24508
rect 5332 24448 5396 24452
rect 5412 24508 5476 24512
rect 5412 24452 5416 24508
rect 5416 24452 5472 24508
rect 5472 24452 5476 24508
rect 5412 24448 5476 24452
rect 13613 24508 13677 24512
rect 13613 24452 13617 24508
rect 13617 24452 13673 24508
rect 13673 24452 13677 24508
rect 13613 24448 13677 24452
rect 13693 24508 13757 24512
rect 13693 24452 13697 24508
rect 13697 24452 13753 24508
rect 13753 24452 13757 24508
rect 13693 24448 13757 24452
rect 13773 24508 13837 24512
rect 13773 24452 13777 24508
rect 13777 24452 13833 24508
rect 13833 24452 13837 24508
rect 13773 24448 13837 24452
rect 13853 24508 13917 24512
rect 13853 24452 13857 24508
rect 13857 24452 13913 24508
rect 13913 24452 13917 24508
rect 13853 24448 13917 24452
rect 22054 24508 22118 24512
rect 22054 24452 22058 24508
rect 22058 24452 22114 24508
rect 22114 24452 22118 24508
rect 22054 24448 22118 24452
rect 22134 24508 22198 24512
rect 22134 24452 22138 24508
rect 22138 24452 22194 24508
rect 22194 24452 22198 24508
rect 22134 24448 22198 24452
rect 22214 24508 22278 24512
rect 22214 24452 22218 24508
rect 22218 24452 22274 24508
rect 22274 24452 22278 24508
rect 22214 24448 22278 24452
rect 22294 24508 22358 24512
rect 22294 24452 22298 24508
rect 22298 24452 22354 24508
rect 22354 24452 22358 24508
rect 22294 24448 22358 24452
rect 30495 24508 30559 24512
rect 30495 24452 30499 24508
rect 30499 24452 30555 24508
rect 30555 24452 30559 24508
rect 30495 24448 30559 24452
rect 30575 24508 30639 24512
rect 30575 24452 30579 24508
rect 30579 24452 30635 24508
rect 30635 24452 30639 24508
rect 30575 24448 30639 24452
rect 30655 24508 30719 24512
rect 30655 24452 30659 24508
rect 30659 24452 30715 24508
rect 30715 24452 30719 24508
rect 30655 24448 30719 24452
rect 30735 24508 30799 24512
rect 30735 24452 30739 24508
rect 30739 24452 30795 24508
rect 30795 24452 30799 24508
rect 30735 24448 30799 24452
rect 9392 23964 9456 23968
rect 9392 23908 9396 23964
rect 9396 23908 9452 23964
rect 9452 23908 9456 23964
rect 9392 23904 9456 23908
rect 9472 23964 9536 23968
rect 9472 23908 9476 23964
rect 9476 23908 9532 23964
rect 9532 23908 9536 23964
rect 9472 23904 9536 23908
rect 9552 23964 9616 23968
rect 9552 23908 9556 23964
rect 9556 23908 9612 23964
rect 9612 23908 9616 23964
rect 9552 23904 9616 23908
rect 9632 23964 9696 23968
rect 9632 23908 9636 23964
rect 9636 23908 9692 23964
rect 9692 23908 9696 23964
rect 9632 23904 9696 23908
rect 17833 23964 17897 23968
rect 17833 23908 17837 23964
rect 17837 23908 17893 23964
rect 17893 23908 17897 23964
rect 17833 23904 17897 23908
rect 17913 23964 17977 23968
rect 17913 23908 17917 23964
rect 17917 23908 17973 23964
rect 17973 23908 17977 23964
rect 17913 23904 17977 23908
rect 17993 23964 18057 23968
rect 17993 23908 17997 23964
rect 17997 23908 18053 23964
rect 18053 23908 18057 23964
rect 17993 23904 18057 23908
rect 18073 23964 18137 23968
rect 18073 23908 18077 23964
rect 18077 23908 18133 23964
rect 18133 23908 18137 23964
rect 18073 23904 18137 23908
rect 26274 23964 26338 23968
rect 26274 23908 26278 23964
rect 26278 23908 26334 23964
rect 26334 23908 26338 23964
rect 26274 23904 26338 23908
rect 26354 23964 26418 23968
rect 26354 23908 26358 23964
rect 26358 23908 26414 23964
rect 26414 23908 26418 23964
rect 26354 23904 26418 23908
rect 26434 23964 26498 23968
rect 26434 23908 26438 23964
rect 26438 23908 26494 23964
rect 26494 23908 26498 23964
rect 26434 23904 26498 23908
rect 26514 23964 26578 23968
rect 26514 23908 26518 23964
rect 26518 23908 26574 23964
rect 26574 23908 26578 23964
rect 26514 23904 26578 23908
rect 34715 23964 34779 23968
rect 34715 23908 34719 23964
rect 34719 23908 34775 23964
rect 34775 23908 34779 23964
rect 34715 23904 34779 23908
rect 34795 23964 34859 23968
rect 34795 23908 34799 23964
rect 34799 23908 34855 23964
rect 34855 23908 34859 23964
rect 34795 23904 34859 23908
rect 34875 23964 34939 23968
rect 34875 23908 34879 23964
rect 34879 23908 34935 23964
rect 34935 23908 34939 23964
rect 34875 23904 34939 23908
rect 34955 23964 35019 23968
rect 34955 23908 34959 23964
rect 34959 23908 35015 23964
rect 35015 23908 35019 23964
rect 34955 23904 35019 23908
rect 5172 23420 5236 23424
rect 5172 23364 5176 23420
rect 5176 23364 5232 23420
rect 5232 23364 5236 23420
rect 5172 23360 5236 23364
rect 5252 23420 5316 23424
rect 5252 23364 5256 23420
rect 5256 23364 5312 23420
rect 5312 23364 5316 23420
rect 5252 23360 5316 23364
rect 5332 23420 5396 23424
rect 5332 23364 5336 23420
rect 5336 23364 5392 23420
rect 5392 23364 5396 23420
rect 5332 23360 5396 23364
rect 5412 23420 5476 23424
rect 5412 23364 5416 23420
rect 5416 23364 5472 23420
rect 5472 23364 5476 23420
rect 5412 23360 5476 23364
rect 13613 23420 13677 23424
rect 13613 23364 13617 23420
rect 13617 23364 13673 23420
rect 13673 23364 13677 23420
rect 13613 23360 13677 23364
rect 13693 23420 13757 23424
rect 13693 23364 13697 23420
rect 13697 23364 13753 23420
rect 13753 23364 13757 23420
rect 13693 23360 13757 23364
rect 13773 23420 13837 23424
rect 13773 23364 13777 23420
rect 13777 23364 13833 23420
rect 13833 23364 13837 23420
rect 13773 23360 13837 23364
rect 13853 23420 13917 23424
rect 13853 23364 13857 23420
rect 13857 23364 13913 23420
rect 13913 23364 13917 23420
rect 13853 23360 13917 23364
rect 22054 23420 22118 23424
rect 22054 23364 22058 23420
rect 22058 23364 22114 23420
rect 22114 23364 22118 23420
rect 22054 23360 22118 23364
rect 22134 23420 22198 23424
rect 22134 23364 22138 23420
rect 22138 23364 22194 23420
rect 22194 23364 22198 23420
rect 22134 23360 22198 23364
rect 22214 23420 22278 23424
rect 22214 23364 22218 23420
rect 22218 23364 22274 23420
rect 22274 23364 22278 23420
rect 22214 23360 22278 23364
rect 22294 23420 22358 23424
rect 22294 23364 22298 23420
rect 22298 23364 22354 23420
rect 22354 23364 22358 23420
rect 22294 23360 22358 23364
rect 30495 23420 30559 23424
rect 30495 23364 30499 23420
rect 30499 23364 30555 23420
rect 30555 23364 30559 23420
rect 30495 23360 30559 23364
rect 30575 23420 30639 23424
rect 30575 23364 30579 23420
rect 30579 23364 30635 23420
rect 30635 23364 30639 23420
rect 30575 23360 30639 23364
rect 30655 23420 30719 23424
rect 30655 23364 30659 23420
rect 30659 23364 30715 23420
rect 30715 23364 30719 23420
rect 30655 23360 30719 23364
rect 30735 23420 30799 23424
rect 30735 23364 30739 23420
rect 30739 23364 30795 23420
rect 30795 23364 30799 23420
rect 30735 23360 30799 23364
rect 9392 22876 9456 22880
rect 9392 22820 9396 22876
rect 9396 22820 9452 22876
rect 9452 22820 9456 22876
rect 9392 22816 9456 22820
rect 9472 22876 9536 22880
rect 9472 22820 9476 22876
rect 9476 22820 9532 22876
rect 9532 22820 9536 22876
rect 9472 22816 9536 22820
rect 9552 22876 9616 22880
rect 9552 22820 9556 22876
rect 9556 22820 9612 22876
rect 9612 22820 9616 22876
rect 9552 22816 9616 22820
rect 9632 22876 9696 22880
rect 9632 22820 9636 22876
rect 9636 22820 9692 22876
rect 9692 22820 9696 22876
rect 9632 22816 9696 22820
rect 17833 22876 17897 22880
rect 17833 22820 17837 22876
rect 17837 22820 17893 22876
rect 17893 22820 17897 22876
rect 17833 22816 17897 22820
rect 17913 22876 17977 22880
rect 17913 22820 17917 22876
rect 17917 22820 17973 22876
rect 17973 22820 17977 22876
rect 17913 22816 17977 22820
rect 17993 22876 18057 22880
rect 17993 22820 17997 22876
rect 17997 22820 18053 22876
rect 18053 22820 18057 22876
rect 17993 22816 18057 22820
rect 18073 22876 18137 22880
rect 18073 22820 18077 22876
rect 18077 22820 18133 22876
rect 18133 22820 18137 22876
rect 18073 22816 18137 22820
rect 26274 22876 26338 22880
rect 26274 22820 26278 22876
rect 26278 22820 26334 22876
rect 26334 22820 26338 22876
rect 26274 22816 26338 22820
rect 26354 22876 26418 22880
rect 26354 22820 26358 22876
rect 26358 22820 26414 22876
rect 26414 22820 26418 22876
rect 26354 22816 26418 22820
rect 26434 22876 26498 22880
rect 26434 22820 26438 22876
rect 26438 22820 26494 22876
rect 26494 22820 26498 22876
rect 26434 22816 26498 22820
rect 26514 22876 26578 22880
rect 26514 22820 26518 22876
rect 26518 22820 26574 22876
rect 26574 22820 26578 22876
rect 26514 22816 26578 22820
rect 34715 22876 34779 22880
rect 34715 22820 34719 22876
rect 34719 22820 34775 22876
rect 34775 22820 34779 22876
rect 34715 22816 34779 22820
rect 34795 22876 34859 22880
rect 34795 22820 34799 22876
rect 34799 22820 34855 22876
rect 34855 22820 34859 22876
rect 34795 22816 34859 22820
rect 34875 22876 34939 22880
rect 34875 22820 34879 22876
rect 34879 22820 34935 22876
rect 34935 22820 34939 22876
rect 34875 22816 34939 22820
rect 34955 22876 35019 22880
rect 34955 22820 34959 22876
rect 34959 22820 35015 22876
rect 35015 22820 35019 22876
rect 34955 22816 35019 22820
rect 5172 22332 5236 22336
rect 5172 22276 5176 22332
rect 5176 22276 5232 22332
rect 5232 22276 5236 22332
rect 5172 22272 5236 22276
rect 5252 22332 5316 22336
rect 5252 22276 5256 22332
rect 5256 22276 5312 22332
rect 5312 22276 5316 22332
rect 5252 22272 5316 22276
rect 5332 22332 5396 22336
rect 5332 22276 5336 22332
rect 5336 22276 5392 22332
rect 5392 22276 5396 22332
rect 5332 22272 5396 22276
rect 5412 22332 5476 22336
rect 5412 22276 5416 22332
rect 5416 22276 5472 22332
rect 5472 22276 5476 22332
rect 5412 22272 5476 22276
rect 13613 22332 13677 22336
rect 13613 22276 13617 22332
rect 13617 22276 13673 22332
rect 13673 22276 13677 22332
rect 13613 22272 13677 22276
rect 13693 22332 13757 22336
rect 13693 22276 13697 22332
rect 13697 22276 13753 22332
rect 13753 22276 13757 22332
rect 13693 22272 13757 22276
rect 13773 22332 13837 22336
rect 13773 22276 13777 22332
rect 13777 22276 13833 22332
rect 13833 22276 13837 22332
rect 13773 22272 13837 22276
rect 13853 22332 13917 22336
rect 13853 22276 13857 22332
rect 13857 22276 13913 22332
rect 13913 22276 13917 22332
rect 13853 22272 13917 22276
rect 22054 22332 22118 22336
rect 22054 22276 22058 22332
rect 22058 22276 22114 22332
rect 22114 22276 22118 22332
rect 22054 22272 22118 22276
rect 22134 22332 22198 22336
rect 22134 22276 22138 22332
rect 22138 22276 22194 22332
rect 22194 22276 22198 22332
rect 22134 22272 22198 22276
rect 22214 22332 22278 22336
rect 22214 22276 22218 22332
rect 22218 22276 22274 22332
rect 22274 22276 22278 22332
rect 22214 22272 22278 22276
rect 22294 22332 22358 22336
rect 22294 22276 22298 22332
rect 22298 22276 22354 22332
rect 22354 22276 22358 22332
rect 22294 22272 22358 22276
rect 30495 22332 30559 22336
rect 30495 22276 30499 22332
rect 30499 22276 30555 22332
rect 30555 22276 30559 22332
rect 30495 22272 30559 22276
rect 30575 22332 30639 22336
rect 30575 22276 30579 22332
rect 30579 22276 30635 22332
rect 30635 22276 30639 22332
rect 30575 22272 30639 22276
rect 30655 22332 30719 22336
rect 30655 22276 30659 22332
rect 30659 22276 30715 22332
rect 30715 22276 30719 22332
rect 30655 22272 30719 22276
rect 30735 22332 30799 22336
rect 30735 22276 30739 22332
rect 30739 22276 30795 22332
rect 30795 22276 30799 22332
rect 30735 22272 30799 22276
rect 9392 21788 9456 21792
rect 9392 21732 9396 21788
rect 9396 21732 9452 21788
rect 9452 21732 9456 21788
rect 9392 21728 9456 21732
rect 9472 21788 9536 21792
rect 9472 21732 9476 21788
rect 9476 21732 9532 21788
rect 9532 21732 9536 21788
rect 9472 21728 9536 21732
rect 9552 21788 9616 21792
rect 9552 21732 9556 21788
rect 9556 21732 9612 21788
rect 9612 21732 9616 21788
rect 9552 21728 9616 21732
rect 9632 21788 9696 21792
rect 9632 21732 9636 21788
rect 9636 21732 9692 21788
rect 9692 21732 9696 21788
rect 9632 21728 9696 21732
rect 17833 21788 17897 21792
rect 17833 21732 17837 21788
rect 17837 21732 17893 21788
rect 17893 21732 17897 21788
rect 17833 21728 17897 21732
rect 17913 21788 17977 21792
rect 17913 21732 17917 21788
rect 17917 21732 17973 21788
rect 17973 21732 17977 21788
rect 17913 21728 17977 21732
rect 17993 21788 18057 21792
rect 17993 21732 17997 21788
rect 17997 21732 18053 21788
rect 18053 21732 18057 21788
rect 17993 21728 18057 21732
rect 18073 21788 18137 21792
rect 18073 21732 18077 21788
rect 18077 21732 18133 21788
rect 18133 21732 18137 21788
rect 18073 21728 18137 21732
rect 26274 21788 26338 21792
rect 26274 21732 26278 21788
rect 26278 21732 26334 21788
rect 26334 21732 26338 21788
rect 26274 21728 26338 21732
rect 26354 21788 26418 21792
rect 26354 21732 26358 21788
rect 26358 21732 26414 21788
rect 26414 21732 26418 21788
rect 26354 21728 26418 21732
rect 26434 21788 26498 21792
rect 26434 21732 26438 21788
rect 26438 21732 26494 21788
rect 26494 21732 26498 21788
rect 26434 21728 26498 21732
rect 26514 21788 26578 21792
rect 26514 21732 26518 21788
rect 26518 21732 26574 21788
rect 26574 21732 26578 21788
rect 26514 21728 26578 21732
rect 34715 21788 34779 21792
rect 34715 21732 34719 21788
rect 34719 21732 34775 21788
rect 34775 21732 34779 21788
rect 34715 21728 34779 21732
rect 34795 21788 34859 21792
rect 34795 21732 34799 21788
rect 34799 21732 34855 21788
rect 34855 21732 34859 21788
rect 34795 21728 34859 21732
rect 34875 21788 34939 21792
rect 34875 21732 34879 21788
rect 34879 21732 34935 21788
rect 34935 21732 34939 21788
rect 34875 21728 34939 21732
rect 34955 21788 35019 21792
rect 34955 21732 34959 21788
rect 34959 21732 35015 21788
rect 35015 21732 35019 21788
rect 34955 21728 35019 21732
rect 5172 21244 5236 21248
rect 5172 21188 5176 21244
rect 5176 21188 5232 21244
rect 5232 21188 5236 21244
rect 5172 21184 5236 21188
rect 5252 21244 5316 21248
rect 5252 21188 5256 21244
rect 5256 21188 5312 21244
rect 5312 21188 5316 21244
rect 5252 21184 5316 21188
rect 5332 21244 5396 21248
rect 5332 21188 5336 21244
rect 5336 21188 5392 21244
rect 5392 21188 5396 21244
rect 5332 21184 5396 21188
rect 5412 21244 5476 21248
rect 5412 21188 5416 21244
rect 5416 21188 5472 21244
rect 5472 21188 5476 21244
rect 5412 21184 5476 21188
rect 13613 21244 13677 21248
rect 13613 21188 13617 21244
rect 13617 21188 13673 21244
rect 13673 21188 13677 21244
rect 13613 21184 13677 21188
rect 13693 21244 13757 21248
rect 13693 21188 13697 21244
rect 13697 21188 13753 21244
rect 13753 21188 13757 21244
rect 13693 21184 13757 21188
rect 13773 21244 13837 21248
rect 13773 21188 13777 21244
rect 13777 21188 13833 21244
rect 13833 21188 13837 21244
rect 13773 21184 13837 21188
rect 13853 21244 13917 21248
rect 13853 21188 13857 21244
rect 13857 21188 13913 21244
rect 13913 21188 13917 21244
rect 13853 21184 13917 21188
rect 22054 21244 22118 21248
rect 22054 21188 22058 21244
rect 22058 21188 22114 21244
rect 22114 21188 22118 21244
rect 22054 21184 22118 21188
rect 22134 21244 22198 21248
rect 22134 21188 22138 21244
rect 22138 21188 22194 21244
rect 22194 21188 22198 21244
rect 22134 21184 22198 21188
rect 22214 21244 22278 21248
rect 22214 21188 22218 21244
rect 22218 21188 22274 21244
rect 22274 21188 22278 21244
rect 22214 21184 22278 21188
rect 22294 21244 22358 21248
rect 22294 21188 22298 21244
rect 22298 21188 22354 21244
rect 22354 21188 22358 21244
rect 22294 21184 22358 21188
rect 30495 21244 30559 21248
rect 30495 21188 30499 21244
rect 30499 21188 30555 21244
rect 30555 21188 30559 21244
rect 30495 21184 30559 21188
rect 30575 21244 30639 21248
rect 30575 21188 30579 21244
rect 30579 21188 30635 21244
rect 30635 21188 30639 21244
rect 30575 21184 30639 21188
rect 30655 21244 30719 21248
rect 30655 21188 30659 21244
rect 30659 21188 30715 21244
rect 30715 21188 30719 21244
rect 30655 21184 30719 21188
rect 30735 21244 30799 21248
rect 30735 21188 30739 21244
rect 30739 21188 30795 21244
rect 30795 21188 30799 21244
rect 30735 21184 30799 21188
rect 9392 20700 9456 20704
rect 9392 20644 9396 20700
rect 9396 20644 9452 20700
rect 9452 20644 9456 20700
rect 9392 20640 9456 20644
rect 9472 20700 9536 20704
rect 9472 20644 9476 20700
rect 9476 20644 9532 20700
rect 9532 20644 9536 20700
rect 9472 20640 9536 20644
rect 9552 20700 9616 20704
rect 9552 20644 9556 20700
rect 9556 20644 9612 20700
rect 9612 20644 9616 20700
rect 9552 20640 9616 20644
rect 9632 20700 9696 20704
rect 9632 20644 9636 20700
rect 9636 20644 9692 20700
rect 9692 20644 9696 20700
rect 9632 20640 9696 20644
rect 17833 20700 17897 20704
rect 17833 20644 17837 20700
rect 17837 20644 17893 20700
rect 17893 20644 17897 20700
rect 17833 20640 17897 20644
rect 17913 20700 17977 20704
rect 17913 20644 17917 20700
rect 17917 20644 17973 20700
rect 17973 20644 17977 20700
rect 17913 20640 17977 20644
rect 17993 20700 18057 20704
rect 17993 20644 17997 20700
rect 17997 20644 18053 20700
rect 18053 20644 18057 20700
rect 17993 20640 18057 20644
rect 18073 20700 18137 20704
rect 18073 20644 18077 20700
rect 18077 20644 18133 20700
rect 18133 20644 18137 20700
rect 18073 20640 18137 20644
rect 26274 20700 26338 20704
rect 26274 20644 26278 20700
rect 26278 20644 26334 20700
rect 26334 20644 26338 20700
rect 26274 20640 26338 20644
rect 26354 20700 26418 20704
rect 26354 20644 26358 20700
rect 26358 20644 26414 20700
rect 26414 20644 26418 20700
rect 26354 20640 26418 20644
rect 26434 20700 26498 20704
rect 26434 20644 26438 20700
rect 26438 20644 26494 20700
rect 26494 20644 26498 20700
rect 26434 20640 26498 20644
rect 26514 20700 26578 20704
rect 26514 20644 26518 20700
rect 26518 20644 26574 20700
rect 26574 20644 26578 20700
rect 26514 20640 26578 20644
rect 34715 20700 34779 20704
rect 34715 20644 34719 20700
rect 34719 20644 34775 20700
rect 34775 20644 34779 20700
rect 34715 20640 34779 20644
rect 34795 20700 34859 20704
rect 34795 20644 34799 20700
rect 34799 20644 34855 20700
rect 34855 20644 34859 20700
rect 34795 20640 34859 20644
rect 34875 20700 34939 20704
rect 34875 20644 34879 20700
rect 34879 20644 34935 20700
rect 34935 20644 34939 20700
rect 34875 20640 34939 20644
rect 34955 20700 35019 20704
rect 34955 20644 34959 20700
rect 34959 20644 35015 20700
rect 35015 20644 35019 20700
rect 34955 20640 35019 20644
rect 5172 20156 5236 20160
rect 5172 20100 5176 20156
rect 5176 20100 5232 20156
rect 5232 20100 5236 20156
rect 5172 20096 5236 20100
rect 5252 20156 5316 20160
rect 5252 20100 5256 20156
rect 5256 20100 5312 20156
rect 5312 20100 5316 20156
rect 5252 20096 5316 20100
rect 5332 20156 5396 20160
rect 5332 20100 5336 20156
rect 5336 20100 5392 20156
rect 5392 20100 5396 20156
rect 5332 20096 5396 20100
rect 5412 20156 5476 20160
rect 5412 20100 5416 20156
rect 5416 20100 5472 20156
rect 5472 20100 5476 20156
rect 5412 20096 5476 20100
rect 13613 20156 13677 20160
rect 13613 20100 13617 20156
rect 13617 20100 13673 20156
rect 13673 20100 13677 20156
rect 13613 20096 13677 20100
rect 13693 20156 13757 20160
rect 13693 20100 13697 20156
rect 13697 20100 13753 20156
rect 13753 20100 13757 20156
rect 13693 20096 13757 20100
rect 13773 20156 13837 20160
rect 13773 20100 13777 20156
rect 13777 20100 13833 20156
rect 13833 20100 13837 20156
rect 13773 20096 13837 20100
rect 13853 20156 13917 20160
rect 13853 20100 13857 20156
rect 13857 20100 13913 20156
rect 13913 20100 13917 20156
rect 13853 20096 13917 20100
rect 22054 20156 22118 20160
rect 22054 20100 22058 20156
rect 22058 20100 22114 20156
rect 22114 20100 22118 20156
rect 22054 20096 22118 20100
rect 22134 20156 22198 20160
rect 22134 20100 22138 20156
rect 22138 20100 22194 20156
rect 22194 20100 22198 20156
rect 22134 20096 22198 20100
rect 22214 20156 22278 20160
rect 22214 20100 22218 20156
rect 22218 20100 22274 20156
rect 22274 20100 22278 20156
rect 22214 20096 22278 20100
rect 22294 20156 22358 20160
rect 22294 20100 22298 20156
rect 22298 20100 22354 20156
rect 22354 20100 22358 20156
rect 22294 20096 22358 20100
rect 30495 20156 30559 20160
rect 30495 20100 30499 20156
rect 30499 20100 30555 20156
rect 30555 20100 30559 20156
rect 30495 20096 30559 20100
rect 30575 20156 30639 20160
rect 30575 20100 30579 20156
rect 30579 20100 30635 20156
rect 30635 20100 30639 20156
rect 30575 20096 30639 20100
rect 30655 20156 30719 20160
rect 30655 20100 30659 20156
rect 30659 20100 30715 20156
rect 30715 20100 30719 20156
rect 30655 20096 30719 20100
rect 30735 20156 30799 20160
rect 30735 20100 30739 20156
rect 30739 20100 30795 20156
rect 30795 20100 30799 20156
rect 30735 20096 30799 20100
rect 9392 19612 9456 19616
rect 9392 19556 9396 19612
rect 9396 19556 9452 19612
rect 9452 19556 9456 19612
rect 9392 19552 9456 19556
rect 9472 19612 9536 19616
rect 9472 19556 9476 19612
rect 9476 19556 9532 19612
rect 9532 19556 9536 19612
rect 9472 19552 9536 19556
rect 9552 19612 9616 19616
rect 9552 19556 9556 19612
rect 9556 19556 9612 19612
rect 9612 19556 9616 19612
rect 9552 19552 9616 19556
rect 9632 19612 9696 19616
rect 9632 19556 9636 19612
rect 9636 19556 9692 19612
rect 9692 19556 9696 19612
rect 9632 19552 9696 19556
rect 17833 19612 17897 19616
rect 17833 19556 17837 19612
rect 17837 19556 17893 19612
rect 17893 19556 17897 19612
rect 17833 19552 17897 19556
rect 17913 19612 17977 19616
rect 17913 19556 17917 19612
rect 17917 19556 17973 19612
rect 17973 19556 17977 19612
rect 17913 19552 17977 19556
rect 17993 19612 18057 19616
rect 17993 19556 17997 19612
rect 17997 19556 18053 19612
rect 18053 19556 18057 19612
rect 17993 19552 18057 19556
rect 18073 19612 18137 19616
rect 18073 19556 18077 19612
rect 18077 19556 18133 19612
rect 18133 19556 18137 19612
rect 18073 19552 18137 19556
rect 26274 19612 26338 19616
rect 26274 19556 26278 19612
rect 26278 19556 26334 19612
rect 26334 19556 26338 19612
rect 26274 19552 26338 19556
rect 26354 19612 26418 19616
rect 26354 19556 26358 19612
rect 26358 19556 26414 19612
rect 26414 19556 26418 19612
rect 26354 19552 26418 19556
rect 26434 19612 26498 19616
rect 26434 19556 26438 19612
rect 26438 19556 26494 19612
rect 26494 19556 26498 19612
rect 26434 19552 26498 19556
rect 26514 19612 26578 19616
rect 26514 19556 26518 19612
rect 26518 19556 26574 19612
rect 26574 19556 26578 19612
rect 26514 19552 26578 19556
rect 34715 19612 34779 19616
rect 34715 19556 34719 19612
rect 34719 19556 34775 19612
rect 34775 19556 34779 19612
rect 34715 19552 34779 19556
rect 34795 19612 34859 19616
rect 34795 19556 34799 19612
rect 34799 19556 34855 19612
rect 34855 19556 34859 19612
rect 34795 19552 34859 19556
rect 34875 19612 34939 19616
rect 34875 19556 34879 19612
rect 34879 19556 34935 19612
rect 34935 19556 34939 19612
rect 34875 19552 34939 19556
rect 34955 19612 35019 19616
rect 34955 19556 34959 19612
rect 34959 19556 35015 19612
rect 35015 19556 35019 19612
rect 34955 19552 35019 19556
rect 5172 19068 5236 19072
rect 5172 19012 5176 19068
rect 5176 19012 5232 19068
rect 5232 19012 5236 19068
rect 5172 19008 5236 19012
rect 5252 19068 5316 19072
rect 5252 19012 5256 19068
rect 5256 19012 5312 19068
rect 5312 19012 5316 19068
rect 5252 19008 5316 19012
rect 5332 19068 5396 19072
rect 5332 19012 5336 19068
rect 5336 19012 5392 19068
rect 5392 19012 5396 19068
rect 5332 19008 5396 19012
rect 5412 19068 5476 19072
rect 5412 19012 5416 19068
rect 5416 19012 5472 19068
rect 5472 19012 5476 19068
rect 5412 19008 5476 19012
rect 13613 19068 13677 19072
rect 13613 19012 13617 19068
rect 13617 19012 13673 19068
rect 13673 19012 13677 19068
rect 13613 19008 13677 19012
rect 13693 19068 13757 19072
rect 13693 19012 13697 19068
rect 13697 19012 13753 19068
rect 13753 19012 13757 19068
rect 13693 19008 13757 19012
rect 13773 19068 13837 19072
rect 13773 19012 13777 19068
rect 13777 19012 13833 19068
rect 13833 19012 13837 19068
rect 13773 19008 13837 19012
rect 13853 19068 13917 19072
rect 13853 19012 13857 19068
rect 13857 19012 13913 19068
rect 13913 19012 13917 19068
rect 13853 19008 13917 19012
rect 22054 19068 22118 19072
rect 22054 19012 22058 19068
rect 22058 19012 22114 19068
rect 22114 19012 22118 19068
rect 22054 19008 22118 19012
rect 22134 19068 22198 19072
rect 22134 19012 22138 19068
rect 22138 19012 22194 19068
rect 22194 19012 22198 19068
rect 22134 19008 22198 19012
rect 22214 19068 22278 19072
rect 22214 19012 22218 19068
rect 22218 19012 22274 19068
rect 22274 19012 22278 19068
rect 22214 19008 22278 19012
rect 22294 19068 22358 19072
rect 22294 19012 22298 19068
rect 22298 19012 22354 19068
rect 22354 19012 22358 19068
rect 22294 19008 22358 19012
rect 30495 19068 30559 19072
rect 30495 19012 30499 19068
rect 30499 19012 30555 19068
rect 30555 19012 30559 19068
rect 30495 19008 30559 19012
rect 30575 19068 30639 19072
rect 30575 19012 30579 19068
rect 30579 19012 30635 19068
rect 30635 19012 30639 19068
rect 30575 19008 30639 19012
rect 30655 19068 30719 19072
rect 30655 19012 30659 19068
rect 30659 19012 30715 19068
rect 30715 19012 30719 19068
rect 30655 19008 30719 19012
rect 30735 19068 30799 19072
rect 30735 19012 30739 19068
rect 30739 19012 30795 19068
rect 30795 19012 30799 19068
rect 30735 19008 30799 19012
rect 9392 18524 9456 18528
rect 9392 18468 9396 18524
rect 9396 18468 9452 18524
rect 9452 18468 9456 18524
rect 9392 18464 9456 18468
rect 9472 18524 9536 18528
rect 9472 18468 9476 18524
rect 9476 18468 9532 18524
rect 9532 18468 9536 18524
rect 9472 18464 9536 18468
rect 9552 18524 9616 18528
rect 9552 18468 9556 18524
rect 9556 18468 9612 18524
rect 9612 18468 9616 18524
rect 9552 18464 9616 18468
rect 9632 18524 9696 18528
rect 9632 18468 9636 18524
rect 9636 18468 9692 18524
rect 9692 18468 9696 18524
rect 9632 18464 9696 18468
rect 17833 18524 17897 18528
rect 17833 18468 17837 18524
rect 17837 18468 17893 18524
rect 17893 18468 17897 18524
rect 17833 18464 17897 18468
rect 17913 18524 17977 18528
rect 17913 18468 17917 18524
rect 17917 18468 17973 18524
rect 17973 18468 17977 18524
rect 17913 18464 17977 18468
rect 17993 18524 18057 18528
rect 17993 18468 17997 18524
rect 17997 18468 18053 18524
rect 18053 18468 18057 18524
rect 17993 18464 18057 18468
rect 18073 18524 18137 18528
rect 18073 18468 18077 18524
rect 18077 18468 18133 18524
rect 18133 18468 18137 18524
rect 18073 18464 18137 18468
rect 26274 18524 26338 18528
rect 26274 18468 26278 18524
rect 26278 18468 26334 18524
rect 26334 18468 26338 18524
rect 26274 18464 26338 18468
rect 26354 18524 26418 18528
rect 26354 18468 26358 18524
rect 26358 18468 26414 18524
rect 26414 18468 26418 18524
rect 26354 18464 26418 18468
rect 26434 18524 26498 18528
rect 26434 18468 26438 18524
rect 26438 18468 26494 18524
rect 26494 18468 26498 18524
rect 26434 18464 26498 18468
rect 26514 18524 26578 18528
rect 26514 18468 26518 18524
rect 26518 18468 26574 18524
rect 26574 18468 26578 18524
rect 26514 18464 26578 18468
rect 34715 18524 34779 18528
rect 34715 18468 34719 18524
rect 34719 18468 34775 18524
rect 34775 18468 34779 18524
rect 34715 18464 34779 18468
rect 34795 18524 34859 18528
rect 34795 18468 34799 18524
rect 34799 18468 34855 18524
rect 34855 18468 34859 18524
rect 34795 18464 34859 18468
rect 34875 18524 34939 18528
rect 34875 18468 34879 18524
rect 34879 18468 34935 18524
rect 34935 18468 34939 18524
rect 34875 18464 34939 18468
rect 34955 18524 35019 18528
rect 34955 18468 34959 18524
rect 34959 18468 35015 18524
rect 35015 18468 35019 18524
rect 34955 18464 35019 18468
rect 5172 17980 5236 17984
rect 5172 17924 5176 17980
rect 5176 17924 5232 17980
rect 5232 17924 5236 17980
rect 5172 17920 5236 17924
rect 5252 17980 5316 17984
rect 5252 17924 5256 17980
rect 5256 17924 5312 17980
rect 5312 17924 5316 17980
rect 5252 17920 5316 17924
rect 5332 17980 5396 17984
rect 5332 17924 5336 17980
rect 5336 17924 5392 17980
rect 5392 17924 5396 17980
rect 5332 17920 5396 17924
rect 5412 17980 5476 17984
rect 5412 17924 5416 17980
rect 5416 17924 5472 17980
rect 5472 17924 5476 17980
rect 5412 17920 5476 17924
rect 13613 17980 13677 17984
rect 13613 17924 13617 17980
rect 13617 17924 13673 17980
rect 13673 17924 13677 17980
rect 13613 17920 13677 17924
rect 13693 17980 13757 17984
rect 13693 17924 13697 17980
rect 13697 17924 13753 17980
rect 13753 17924 13757 17980
rect 13693 17920 13757 17924
rect 13773 17980 13837 17984
rect 13773 17924 13777 17980
rect 13777 17924 13833 17980
rect 13833 17924 13837 17980
rect 13773 17920 13837 17924
rect 13853 17980 13917 17984
rect 13853 17924 13857 17980
rect 13857 17924 13913 17980
rect 13913 17924 13917 17980
rect 13853 17920 13917 17924
rect 22054 17980 22118 17984
rect 22054 17924 22058 17980
rect 22058 17924 22114 17980
rect 22114 17924 22118 17980
rect 22054 17920 22118 17924
rect 22134 17980 22198 17984
rect 22134 17924 22138 17980
rect 22138 17924 22194 17980
rect 22194 17924 22198 17980
rect 22134 17920 22198 17924
rect 22214 17980 22278 17984
rect 22214 17924 22218 17980
rect 22218 17924 22274 17980
rect 22274 17924 22278 17980
rect 22214 17920 22278 17924
rect 22294 17980 22358 17984
rect 22294 17924 22298 17980
rect 22298 17924 22354 17980
rect 22354 17924 22358 17980
rect 22294 17920 22358 17924
rect 30495 17980 30559 17984
rect 30495 17924 30499 17980
rect 30499 17924 30555 17980
rect 30555 17924 30559 17980
rect 30495 17920 30559 17924
rect 30575 17980 30639 17984
rect 30575 17924 30579 17980
rect 30579 17924 30635 17980
rect 30635 17924 30639 17980
rect 30575 17920 30639 17924
rect 30655 17980 30719 17984
rect 30655 17924 30659 17980
rect 30659 17924 30715 17980
rect 30715 17924 30719 17980
rect 30655 17920 30719 17924
rect 30735 17980 30799 17984
rect 30735 17924 30739 17980
rect 30739 17924 30795 17980
rect 30795 17924 30799 17980
rect 30735 17920 30799 17924
rect 9392 17436 9456 17440
rect 9392 17380 9396 17436
rect 9396 17380 9452 17436
rect 9452 17380 9456 17436
rect 9392 17376 9456 17380
rect 9472 17436 9536 17440
rect 9472 17380 9476 17436
rect 9476 17380 9532 17436
rect 9532 17380 9536 17436
rect 9472 17376 9536 17380
rect 9552 17436 9616 17440
rect 9552 17380 9556 17436
rect 9556 17380 9612 17436
rect 9612 17380 9616 17436
rect 9552 17376 9616 17380
rect 9632 17436 9696 17440
rect 9632 17380 9636 17436
rect 9636 17380 9692 17436
rect 9692 17380 9696 17436
rect 9632 17376 9696 17380
rect 17833 17436 17897 17440
rect 17833 17380 17837 17436
rect 17837 17380 17893 17436
rect 17893 17380 17897 17436
rect 17833 17376 17897 17380
rect 17913 17436 17977 17440
rect 17913 17380 17917 17436
rect 17917 17380 17973 17436
rect 17973 17380 17977 17436
rect 17913 17376 17977 17380
rect 17993 17436 18057 17440
rect 17993 17380 17997 17436
rect 17997 17380 18053 17436
rect 18053 17380 18057 17436
rect 17993 17376 18057 17380
rect 18073 17436 18137 17440
rect 18073 17380 18077 17436
rect 18077 17380 18133 17436
rect 18133 17380 18137 17436
rect 18073 17376 18137 17380
rect 26274 17436 26338 17440
rect 26274 17380 26278 17436
rect 26278 17380 26334 17436
rect 26334 17380 26338 17436
rect 26274 17376 26338 17380
rect 26354 17436 26418 17440
rect 26354 17380 26358 17436
rect 26358 17380 26414 17436
rect 26414 17380 26418 17436
rect 26354 17376 26418 17380
rect 26434 17436 26498 17440
rect 26434 17380 26438 17436
rect 26438 17380 26494 17436
rect 26494 17380 26498 17436
rect 26434 17376 26498 17380
rect 26514 17436 26578 17440
rect 26514 17380 26518 17436
rect 26518 17380 26574 17436
rect 26574 17380 26578 17436
rect 26514 17376 26578 17380
rect 34715 17436 34779 17440
rect 34715 17380 34719 17436
rect 34719 17380 34775 17436
rect 34775 17380 34779 17436
rect 34715 17376 34779 17380
rect 34795 17436 34859 17440
rect 34795 17380 34799 17436
rect 34799 17380 34855 17436
rect 34855 17380 34859 17436
rect 34795 17376 34859 17380
rect 34875 17436 34939 17440
rect 34875 17380 34879 17436
rect 34879 17380 34935 17436
rect 34935 17380 34939 17436
rect 34875 17376 34939 17380
rect 34955 17436 35019 17440
rect 34955 17380 34959 17436
rect 34959 17380 35015 17436
rect 35015 17380 35019 17436
rect 34955 17376 35019 17380
rect 5172 16892 5236 16896
rect 5172 16836 5176 16892
rect 5176 16836 5232 16892
rect 5232 16836 5236 16892
rect 5172 16832 5236 16836
rect 5252 16892 5316 16896
rect 5252 16836 5256 16892
rect 5256 16836 5312 16892
rect 5312 16836 5316 16892
rect 5252 16832 5316 16836
rect 5332 16892 5396 16896
rect 5332 16836 5336 16892
rect 5336 16836 5392 16892
rect 5392 16836 5396 16892
rect 5332 16832 5396 16836
rect 5412 16892 5476 16896
rect 5412 16836 5416 16892
rect 5416 16836 5472 16892
rect 5472 16836 5476 16892
rect 5412 16832 5476 16836
rect 13613 16892 13677 16896
rect 13613 16836 13617 16892
rect 13617 16836 13673 16892
rect 13673 16836 13677 16892
rect 13613 16832 13677 16836
rect 13693 16892 13757 16896
rect 13693 16836 13697 16892
rect 13697 16836 13753 16892
rect 13753 16836 13757 16892
rect 13693 16832 13757 16836
rect 13773 16892 13837 16896
rect 13773 16836 13777 16892
rect 13777 16836 13833 16892
rect 13833 16836 13837 16892
rect 13773 16832 13837 16836
rect 13853 16892 13917 16896
rect 13853 16836 13857 16892
rect 13857 16836 13913 16892
rect 13913 16836 13917 16892
rect 13853 16832 13917 16836
rect 22054 16892 22118 16896
rect 22054 16836 22058 16892
rect 22058 16836 22114 16892
rect 22114 16836 22118 16892
rect 22054 16832 22118 16836
rect 22134 16892 22198 16896
rect 22134 16836 22138 16892
rect 22138 16836 22194 16892
rect 22194 16836 22198 16892
rect 22134 16832 22198 16836
rect 22214 16892 22278 16896
rect 22214 16836 22218 16892
rect 22218 16836 22274 16892
rect 22274 16836 22278 16892
rect 22214 16832 22278 16836
rect 22294 16892 22358 16896
rect 22294 16836 22298 16892
rect 22298 16836 22354 16892
rect 22354 16836 22358 16892
rect 22294 16832 22358 16836
rect 30495 16892 30559 16896
rect 30495 16836 30499 16892
rect 30499 16836 30555 16892
rect 30555 16836 30559 16892
rect 30495 16832 30559 16836
rect 30575 16892 30639 16896
rect 30575 16836 30579 16892
rect 30579 16836 30635 16892
rect 30635 16836 30639 16892
rect 30575 16832 30639 16836
rect 30655 16892 30719 16896
rect 30655 16836 30659 16892
rect 30659 16836 30715 16892
rect 30715 16836 30719 16892
rect 30655 16832 30719 16836
rect 30735 16892 30799 16896
rect 30735 16836 30739 16892
rect 30739 16836 30795 16892
rect 30795 16836 30799 16892
rect 30735 16832 30799 16836
rect 9392 16348 9456 16352
rect 9392 16292 9396 16348
rect 9396 16292 9452 16348
rect 9452 16292 9456 16348
rect 9392 16288 9456 16292
rect 9472 16348 9536 16352
rect 9472 16292 9476 16348
rect 9476 16292 9532 16348
rect 9532 16292 9536 16348
rect 9472 16288 9536 16292
rect 9552 16348 9616 16352
rect 9552 16292 9556 16348
rect 9556 16292 9612 16348
rect 9612 16292 9616 16348
rect 9552 16288 9616 16292
rect 9632 16348 9696 16352
rect 9632 16292 9636 16348
rect 9636 16292 9692 16348
rect 9692 16292 9696 16348
rect 9632 16288 9696 16292
rect 17833 16348 17897 16352
rect 17833 16292 17837 16348
rect 17837 16292 17893 16348
rect 17893 16292 17897 16348
rect 17833 16288 17897 16292
rect 17913 16348 17977 16352
rect 17913 16292 17917 16348
rect 17917 16292 17973 16348
rect 17973 16292 17977 16348
rect 17913 16288 17977 16292
rect 17993 16348 18057 16352
rect 17993 16292 17997 16348
rect 17997 16292 18053 16348
rect 18053 16292 18057 16348
rect 17993 16288 18057 16292
rect 18073 16348 18137 16352
rect 18073 16292 18077 16348
rect 18077 16292 18133 16348
rect 18133 16292 18137 16348
rect 18073 16288 18137 16292
rect 26274 16348 26338 16352
rect 26274 16292 26278 16348
rect 26278 16292 26334 16348
rect 26334 16292 26338 16348
rect 26274 16288 26338 16292
rect 26354 16348 26418 16352
rect 26354 16292 26358 16348
rect 26358 16292 26414 16348
rect 26414 16292 26418 16348
rect 26354 16288 26418 16292
rect 26434 16348 26498 16352
rect 26434 16292 26438 16348
rect 26438 16292 26494 16348
rect 26494 16292 26498 16348
rect 26434 16288 26498 16292
rect 26514 16348 26578 16352
rect 26514 16292 26518 16348
rect 26518 16292 26574 16348
rect 26574 16292 26578 16348
rect 26514 16288 26578 16292
rect 34715 16348 34779 16352
rect 34715 16292 34719 16348
rect 34719 16292 34775 16348
rect 34775 16292 34779 16348
rect 34715 16288 34779 16292
rect 34795 16348 34859 16352
rect 34795 16292 34799 16348
rect 34799 16292 34855 16348
rect 34855 16292 34859 16348
rect 34795 16288 34859 16292
rect 34875 16348 34939 16352
rect 34875 16292 34879 16348
rect 34879 16292 34935 16348
rect 34935 16292 34939 16348
rect 34875 16288 34939 16292
rect 34955 16348 35019 16352
rect 34955 16292 34959 16348
rect 34959 16292 35015 16348
rect 35015 16292 35019 16348
rect 34955 16288 35019 16292
rect 5172 15804 5236 15808
rect 5172 15748 5176 15804
rect 5176 15748 5232 15804
rect 5232 15748 5236 15804
rect 5172 15744 5236 15748
rect 5252 15804 5316 15808
rect 5252 15748 5256 15804
rect 5256 15748 5312 15804
rect 5312 15748 5316 15804
rect 5252 15744 5316 15748
rect 5332 15804 5396 15808
rect 5332 15748 5336 15804
rect 5336 15748 5392 15804
rect 5392 15748 5396 15804
rect 5332 15744 5396 15748
rect 5412 15804 5476 15808
rect 5412 15748 5416 15804
rect 5416 15748 5472 15804
rect 5472 15748 5476 15804
rect 5412 15744 5476 15748
rect 13613 15804 13677 15808
rect 13613 15748 13617 15804
rect 13617 15748 13673 15804
rect 13673 15748 13677 15804
rect 13613 15744 13677 15748
rect 13693 15804 13757 15808
rect 13693 15748 13697 15804
rect 13697 15748 13753 15804
rect 13753 15748 13757 15804
rect 13693 15744 13757 15748
rect 13773 15804 13837 15808
rect 13773 15748 13777 15804
rect 13777 15748 13833 15804
rect 13833 15748 13837 15804
rect 13773 15744 13837 15748
rect 13853 15804 13917 15808
rect 13853 15748 13857 15804
rect 13857 15748 13913 15804
rect 13913 15748 13917 15804
rect 13853 15744 13917 15748
rect 22054 15804 22118 15808
rect 22054 15748 22058 15804
rect 22058 15748 22114 15804
rect 22114 15748 22118 15804
rect 22054 15744 22118 15748
rect 22134 15804 22198 15808
rect 22134 15748 22138 15804
rect 22138 15748 22194 15804
rect 22194 15748 22198 15804
rect 22134 15744 22198 15748
rect 22214 15804 22278 15808
rect 22214 15748 22218 15804
rect 22218 15748 22274 15804
rect 22274 15748 22278 15804
rect 22214 15744 22278 15748
rect 22294 15804 22358 15808
rect 22294 15748 22298 15804
rect 22298 15748 22354 15804
rect 22354 15748 22358 15804
rect 22294 15744 22358 15748
rect 30495 15804 30559 15808
rect 30495 15748 30499 15804
rect 30499 15748 30555 15804
rect 30555 15748 30559 15804
rect 30495 15744 30559 15748
rect 30575 15804 30639 15808
rect 30575 15748 30579 15804
rect 30579 15748 30635 15804
rect 30635 15748 30639 15804
rect 30575 15744 30639 15748
rect 30655 15804 30719 15808
rect 30655 15748 30659 15804
rect 30659 15748 30715 15804
rect 30715 15748 30719 15804
rect 30655 15744 30719 15748
rect 30735 15804 30799 15808
rect 30735 15748 30739 15804
rect 30739 15748 30795 15804
rect 30795 15748 30799 15804
rect 30735 15744 30799 15748
rect 9392 15260 9456 15264
rect 9392 15204 9396 15260
rect 9396 15204 9452 15260
rect 9452 15204 9456 15260
rect 9392 15200 9456 15204
rect 9472 15260 9536 15264
rect 9472 15204 9476 15260
rect 9476 15204 9532 15260
rect 9532 15204 9536 15260
rect 9472 15200 9536 15204
rect 9552 15260 9616 15264
rect 9552 15204 9556 15260
rect 9556 15204 9612 15260
rect 9612 15204 9616 15260
rect 9552 15200 9616 15204
rect 9632 15260 9696 15264
rect 9632 15204 9636 15260
rect 9636 15204 9692 15260
rect 9692 15204 9696 15260
rect 9632 15200 9696 15204
rect 17833 15260 17897 15264
rect 17833 15204 17837 15260
rect 17837 15204 17893 15260
rect 17893 15204 17897 15260
rect 17833 15200 17897 15204
rect 17913 15260 17977 15264
rect 17913 15204 17917 15260
rect 17917 15204 17973 15260
rect 17973 15204 17977 15260
rect 17913 15200 17977 15204
rect 17993 15260 18057 15264
rect 17993 15204 17997 15260
rect 17997 15204 18053 15260
rect 18053 15204 18057 15260
rect 17993 15200 18057 15204
rect 18073 15260 18137 15264
rect 18073 15204 18077 15260
rect 18077 15204 18133 15260
rect 18133 15204 18137 15260
rect 18073 15200 18137 15204
rect 26274 15260 26338 15264
rect 26274 15204 26278 15260
rect 26278 15204 26334 15260
rect 26334 15204 26338 15260
rect 26274 15200 26338 15204
rect 26354 15260 26418 15264
rect 26354 15204 26358 15260
rect 26358 15204 26414 15260
rect 26414 15204 26418 15260
rect 26354 15200 26418 15204
rect 26434 15260 26498 15264
rect 26434 15204 26438 15260
rect 26438 15204 26494 15260
rect 26494 15204 26498 15260
rect 26434 15200 26498 15204
rect 26514 15260 26578 15264
rect 26514 15204 26518 15260
rect 26518 15204 26574 15260
rect 26574 15204 26578 15260
rect 26514 15200 26578 15204
rect 34715 15260 34779 15264
rect 34715 15204 34719 15260
rect 34719 15204 34775 15260
rect 34775 15204 34779 15260
rect 34715 15200 34779 15204
rect 34795 15260 34859 15264
rect 34795 15204 34799 15260
rect 34799 15204 34855 15260
rect 34855 15204 34859 15260
rect 34795 15200 34859 15204
rect 34875 15260 34939 15264
rect 34875 15204 34879 15260
rect 34879 15204 34935 15260
rect 34935 15204 34939 15260
rect 34875 15200 34939 15204
rect 34955 15260 35019 15264
rect 34955 15204 34959 15260
rect 34959 15204 35015 15260
rect 35015 15204 35019 15260
rect 34955 15200 35019 15204
rect 5172 14716 5236 14720
rect 5172 14660 5176 14716
rect 5176 14660 5232 14716
rect 5232 14660 5236 14716
rect 5172 14656 5236 14660
rect 5252 14716 5316 14720
rect 5252 14660 5256 14716
rect 5256 14660 5312 14716
rect 5312 14660 5316 14716
rect 5252 14656 5316 14660
rect 5332 14716 5396 14720
rect 5332 14660 5336 14716
rect 5336 14660 5392 14716
rect 5392 14660 5396 14716
rect 5332 14656 5396 14660
rect 5412 14716 5476 14720
rect 5412 14660 5416 14716
rect 5416 14660 5472 14716
rect 5472 14660 5476 14716
rect 5412 14656 5476 14660
rect 13613 14716 13677 14720
rect 13613 14660 13617 14716
rect 13617 14660 13673 14716
rect 13673 14660 13677 14716
rect 13613 14656 13677 14660
rect 13693 14716 13757 14720
rect 13693 14660 13697 14716
rect 13697 14660 13753 14716
rect 13753 14660 13757 14716
rect 13693 14656 13757 14660
rect 13773 14716 13837 14720
rect 13773 14660 13777 14716
rect 13777 14660 13833 14716
rect 13833 14660 13837 14716
rect 13773 14656 13837 14660
rect 13853 14716 13917 14720
rect 13853 14660 13857 14716
rect 13857 14660 13913 14716
rect 13913 14660 13917 14716
rect 13853 14656 13917 14660
rect 22054 14716 22118 14720
rect 22054 14660 22058 14716
rect 22058 14660 22114 14716
rect 22114 14660 22118 14716
rect 22054 14656 22118 14660
rect 22134 14716 22198 14720
rect 22134 14660 22138 14716
rect 22138 14660 22194 14716
rect 22194 14660 22198 14716
rect 22134 14656 22198 14660
rect 22214 14716 22278 14720
rect 22214 14660 22218 14716
rect 22218 14660 22274 14716
rect 22274 14660 22278 14716
rect 22214 14656 22278 14660
rect 22294 14716 22358 14720
rect 22294 14660 22298 14716
rect 22298 14660 22354 14716
rect 22354 14660 22358 14716
rect 22294 14656 22358 14660
rect 30495 14716 30559 14720
rect 30495 14660 30499 14716
rect 30499 14660 30555 14716
rect 30555 14660 30559 14716
rect 30495 14656 30559 14660
rect 30575 14716 30639 14720
rect 30575 14660 30579 14716
rect 30579 14660 30635 14716
rect 30635 14660 30639 14716
rect 30575 14656 30639 14660
rect 30655 14716 30719 14720
rect 30655 14660 30659 14716
rect 30659 14660 30715 14716
rect 30715 14660 30719 14716
rect 30655 14656 30719 14660
rect 30735 14716 30799 14720
rect 30735 14660 30739 14716
rect 30739 14660 30795 14716
rect 30795 14660 30799 14716
rect 30735 14656 30799 14660
rect 9392 14172 9456 14176
rect 9392 14116 9396 14172
rect 9396 14116 9452 14172
rect 9452 14116 9456 14172
rect 9392 14112 9456 14116
rect 9472 14172 9536 14176
rect 9472 14116 9476 14172
rect 9476 14116 9532 14172
rect 9532 14116 9536 14172
rect 9472 14112 9536 14116
rect 9552 14172 9616 14176
rect 9552 14116 9556 14172
rect 9556 14116 9612 14172
rect 9612 14116 9616 14172
rect 9552 14112 9616 14116
rect 9632 14172 9696 14176
rect 9632 14116 9636 14172
rect 9636 14116 9692 14172
rect 9692 14116 9696 14172
rect 9632 14112 9696 14116
rect 17833 14172 17897 14176
rect 17833 14116 17837 14172
rect 17837 14116 17893 14172
rect 17893 14116 17897 14172
rect 17833 14112 17897 14116
rect 17913 14172 17977 14176
rect 17913 14116 17917 14172
rect 17917 14116 17973 14172
rect 17973 14116 17977 14172
rect 17913 14112 17977 14116
rect 17993 14172 18057 14176
rect 17993 14116 17997 14172
rect 17997 14116 18053 14172
rect 18053 14116 18057 14172
rect 17993 14112 18057 14116
rect 18073 14172 18137 14176
rect 18073 14116 18077 14172
rect 18077 14116 18133 14172
rect 18133 14116 18137 14172
rect 18073 14112 18137 14116
rect 26274 14172 26338 14176
rect 26274 14116 26278 14172
rect 26278 14116 26334 14172
rect 26334 14116 26338 14172
rect 26274 14112 26338 14116
rect 26354 14172 26418 14176
rect 26354 14116 26358 14172
rect 26358 14116 26414 14172
rect 26414 14116 26418 14172
rect 26354 14112 26418 14116
rect 26434 14172 26498 14176
rect 26434 14116 26438 14172
rect 26438 14116 26494 14172
rect 26494 14116 26498 14172
rect 26434 14112 26498 14116
rect 26514 14172 26578 14176
rect 26514 14116 26518 14172
rect 26518 14116 26574 14172
rect 26574 14116 26578 14172
rect 26514 14112 26578 14116
rect 34715 14172 34779 14176
rect 34715 14116 34719 14172
rect 34719 14116 34775 14172
rect 34775 14116 34779 14172
rect 34715 14112 34779 14116
rect 34795 14172 34859 14176
rect 34795 14116 34799 14172
rect 34799 14116 34855 14172
rect 34855 14116 34859 14172
rect 34795 14112 34859 14116
rect 34875 14172 34939 14176
rect 34875 14116 34879 14172
rect 34879 14116 34935 14172
rect 34935 14116 34939 14172
rect 34875 14112 34939 14116
rect 34955 14172 35019 14176
rect 34955 14116 34959 14172
rect 34959 14116 35015 14172
rect 35015 14116 35019 14172
rect 34955 14112 35019 14116
rect 5172 13628 5236 13632
rect 5172 13572 5176 13628
rect 5176 13572 5232 13628
rect 5232 13572 5236 13628
rect 5172 13568 5236 13572
rect 5252 13628 5316 13632
rect 5252 13572 5256 13628
rect 5256 13572 5312 13628
rect 5312 13572 5316 13628
rect 5252 13568 5316 13572
rect 5332 13628 5396 13632
rect 5332 13572 5336 13628
rect 5336 13572 5392 13628
rect 5392 13572 5396 13628
rect 5332 13568 5396 13572
rect 5412 13628 5476 13632
rect 5412 13572 5416 13628
rect 5416 13572 5472 13628
rect 5472 13572 5476 13628
rect 5412 13568 5476 13572
rect 13613 13628 13677 13632
rect 13613 13572 13617 13628
rect 13617 13572 13673 13628
rect 13673 13572 13677 13628
rect 13613 13568 13677 13572
rect 13693 13628 13757 13632
rect 13693 13572 13697 13628
rect 13697 13572 13753 13628
rect 13753 13572 13757 13628
rect 13693 13568 13757 13572
rect 13773 13628 13837 13632
rect 13773 13572 13777 13628
rect 13777 13572 13833 13628
rect 13833 13572 13837 13628
rect 13773 13568 13837 13572
rect 13853 13628 13917 13632
rect 13853 13572 13857 13628
rect 13857 13572 13913 13628
rect 13913 13572 13917 13628
rect 13853 13568 13917 13572
rect 22054 13628 22118 13632
rect 22054 13572 22058 13628
rect 22058 13572 22114 13628
rect 22114 13572 22118 13628
rect 22054 13568 22118 13572
rect 22134 13628 22198 13632
rect 22134 13572 22138 13628
rect 22138 13572 22194 13628
rect 22194 13572 22198 13628
rect 22134 13568 22198 13572
rect 22214 13628 22278 13632
rect 22214 13572 22218 13628
rect 22218 13572 22274 13628
rect 22274 13572 22278 13628
rect 22214 13568 22278 13572
rect 22294 13628 22358 13632
rect 22294 13572 22298 13628
rect 22298 13572 22354 13628
rect 22354 13572 22358 13628
rect 22294 13568 22358 13572
rect 30495 13628 30559 13632
rect 30495 13572 30499 13628
rect 30499 13572 30555 13628
rect 30555 13572 30559 13628
rect 30495 13568 30559 13572
rect 30575 13628 30639 13632
rect 30575 13572 30579 13628
rect 30579 13572 30635 13628
rect 30635 13572 30639 13628
rect 30575 13568 30639 13572
rect 30655 13628 30719 13632
rect 30655 13572 30659 13628
rect 30659 13572 30715 13628
rect 30715 13572 30719 13628
rect 30655 13568 30719 13572
rect 30735 13628 30799 13632
rect 30735 13572 30739 13628
rect 30739 13572 30795 13628
rect 30795 13572 30799 13628
rect 30735 13568 30799 13572
rect 9392 13084 9456 13088
rect 9392 13028 9396 13084
rect 9396 13028 9452 13084
rect 9452 13028 9456 13084
rect 9392 13024 9456 13028
rect 9472 13084 9536 13088
rect 9472 13028 9476 13084
rect 9476 13028 9532 13084
rect 9532 13028 9536 13084
rect 9472 13024 9536 13028
rect 9552 13084 9616 13088
rect 9552 13028 9556 13084
rect 9556 13028 9612 13084
rect 9612 13028 9616 13084
rect 9552 13024 9616 13028
rect 9632 13084 9696 13088
rect 9632 13028 9636 13084
rect 9636 13028 9692 13084
rect 9692 13028 9696 13084
rect 9632 13024 9696 13028
rect 17833 13084 17897 13088
rect 17833 13028 17837 13084
rect 17837 13028 17893 13084
rect 17893 13028 17897 13084
rect 17833 13024 17897 13028
rect 17913 13084 17977 13088
rect 17913 13028 17917 13084
rect 17917 13028 17973 13084
rect 17973 13028 17977 13084
rect 17913 13024 17977 13028
rect 17993 13084 18057 13088
rect 17993 13028 17997 13084
rect 17997 13028 18053 13084
rect 18053 13028 18057 13084
rect 17993 13024 18057 13028
rect 18073 13084 18137 13088
rect 18073 13028 18077 13084
rect 18077 13028 18133 13084
rect 18133 13028 18137 13084
rect 18073 13024 18137 13028
rect 26274 13084 26338 13088
rect 26274 13028 26278 13084
rect 26278 13028 26334 13084
rect 26334 13028 26338 13084
rect 26274 13024 26338 13028
rect 26354 13084 26418 13088
rect 26354 13028 26358 13084
rect 26358 13028 26414 13084
rect 26414 13028 26418 13084
rect 26354 13024 26418 13028
rect 26434 13084 26498 13088
rect 26434 13028 26438 13084
rect 26438 13028 26494 13084
rect 26494 13028 26498 13084
rect 26434 13024 26498 13028
rect 26514 13084 26578 13088
rect 26514 13028 26518 13084
rect 26518 13028 26574 13084
rect 26574 13028 26578 13084
rect 26514 13024 26578 13028
rect 34715 13084 34779 13088
rect 34715 13028 34719 13084
rect 34719 13028 34775 13084
rect 34775 13028 34779 13084
rect 34715 13024 34779 13028
rect 34795 13084 34859 13088
rect 34795 13028 34799 13084
rect 34799 13028 34855 13084
rect 34855 13028 34859 13084
rect 34795 13024 34859 13028
rect 34875 13084 34939 13088
rect 34875 13028 34879 13084
rect 34879 13028 34935 13084
rect 34935 13028 34939 13084
rect 34875 13024 34939 13028
rect 34955 13084 35019 13088
rect 34955 13028 34959 13084
rect 34959 13028 35015 13084
rect 35015 13028 35019 13084
rect 34955 13024 35019 13028
rect 5172 12540 5236 12544
rect 5172 12484 5176 12540
rect 5176 12484 5232 12540
rect 5232 12484 5236 12540
rect 5172 12480 5236 12484
rect 5252 12540 5316 12544
rect 5252 12484 5256 12540
rect 5256 12484 5312 12540
rect 5312 12484 5316 12540
rect 5252 12480 5316 12484
rect 5332 12540 5396 12544
rect 5332 12484 5336 12540
rect 5336 12484 5392 12540
rect 5392 12484 5396 12540
rect 5332 12480 5396 12484
rect 5412 12540 5476 12544
rect 5412 12484 5416 12540
rect 5416 12484 5472 12540
rect 5472 12484 5476 12540
rect 5412 12480 5476 12484
rect 13613 12540 13677 12544
rect 13613 12484 13617 12540
rect 13617 12484 13673 12540
rect 13673 12484 13677 12540
rect 13613 12480 13677 12484
rect 13693 12540 13757 12544
rect 13693 12484 13697 12540
rect 13697 12484 13753 12540
rect 13753 12484 13757 12540
rect 13693 12480 13757 12484
rect 13773 12540 13837 12544
rect 13773 12484 13777 12540
rect 13777 12484 13833 12540
rect 13833 12484 13837 12540
rect 13773 12480 13837 12484
rect 13853 12540 13917 12544
rect 13853 12484 13857 12540
rect 13857 12484 13913 12540
rect 13913 12484 13917 12540
rect 13853 12480 13917 12484
rect 22054 12540 22118 12544
rect 22054 12484 22058 12540
rect 22058 12484 22114 12540
rect 22114 12484 22118 12540
rect 22054 12480 22118 12484
rect 22134 12540 22198 12544
rect 22134 12484 22138 12540
rect 22138 12484 22194 12540
rect 22194 12484 22198 12540
rect 22134 12480 22198 12484
rect 22214 12540 22278 12544
rect 22214 12484 22218 12540
rect 22218 12484 22274 12540
rect 22274 12484 22278 12540
rect 22214 12480 22278 12484
rect 22294 12540 22358 12544
rect 22294 12484 22298 12540
rect 22298 12484 22354 12540
rect 22354 12484 22358 12540
rect 22294 12480 22358 12484
rect 30495 12540 30559 12544
rect 30495 12484 30499 12540
rect 30499 12484 30555 12540
rect 30555 12484 30559 12540
rect 30495 12480 30559 12484
rect 30575 12540 30639 12544
rect 30575 12484 30579 12540
rect 30579 12484 30635 12540
rect 30635 12484 30639 12540
rect 30575 12480 30639 12484
rect 30655 12540 30719 12544
rect 30655 12484 30659 12540
rect 30659 12484 30715 12540
rect 30715 12484 30719 12540
rect 30655 12480 30719 12484
rect 30735 12540 30799 12544
rect 30735 12484 30739 12540
rect 30739 12484 30795 12540
rect 30795 12484 30799 12540
rect 30735 12480 30799 12484
rect 9392 11996 9456 12000
rect 9392 11940 9396 11996
rect 9396 11940 9452 11996
rect 9452 11940 9456 11996
rect 9392 11936 9456 11940
rect 9472 11996 9536 12000
rect 9472 11940 9476 11996
rect 9476 11940 9532 11996
rect 9532 11940 9536 11996
rect 9472 11936 9536 11940
rect 9552 11996 9616 12000
rect 9552 11940 9556 11996
rect 9556 11940 9612 11996
rect 9612 11940 9616 11996
rect 9552 11936 9616 11940
rect 9632 11996 9696 12000
rect 9632 11940 9636 11996
rect 9636 11940 9692 11996
rect 9692 11940 9696 11996
rect 9632 11936 9696 11940
rect 17833 11996 17897 12000
rect 17833 11940 17837 11996
rect 17837 11940 17893 11996
rect 17893 11940 17897 11996
rect 17833 11936 17897 11940
rect 17913 11996 17977 12000
rect 17913 11940 17917 11996
rect 17917 11940 17973 11996
rect 17973 11940 17977 11996
rect 17913 11936 17977 11940
rect 17993 11996 18057 12000
rect 17993 11940 17997 11996
rect 17997 11940 18053 11996
rect 18053 11940 18057 11996
rect 17993 11936 18057 11940
rect 18073 11996 18137 12000
rect 18073 11940 18077 11996
rect 18077 11940 18133 11996
rect 18133 11940 18137 11996
rect 18073 11936 18137 11940
rect 26274 11996 26338 12000
rect 26274 11940 26278 11996
rect 26278 11940 26334 11996
rect 26334 11940 26338 11996
rect 26274 11936 26338 11940
rect 26354 11996 26418 12000
rect 26354 11940 26358 11996
rect 26358 11940 26414 11996
rect 26414 11940 26418 11996
rect 26354 11936 26418 11940
rect 26434 11996 26498 12000
rect 26434 11940 26438 11996
rect 26438 11940 26494 11996
rect 26494 11940 26498 11996
rect 26434 11936 26498 11940
rect 26514 11996 26578 12000
rect 26514 11940 26518 11996
rect 26518 11940 26574 11996
rect 26574 11940 26578 11996
rect 26514 11936 26578 11940
rect 34715 11996 34779 12000
rect 34715 11940 34719 11996
rect 34719 11940 34775 11996
rect 34775 11940 34779 11996
rect 34715 11936 34779 11940
rect 34795 11996 34859 12000
rect 34795 11940 34799 11996
rect 34799 11940 34855 11996
rect 34855 11940 34859 11996
rect 34795 11936 34859 11940
rect 34875 11996 34939 12000
rect 34875 11940 34879 11996
rect 34879 11940 34935 11996
rect 34935 11940 34939 11996
rect 34875 11936 34939 11940
rect 34955 11996 35019 12000
rect 34955 11940 34959 11996
rect 34959 11940 35015 11996
rect 35015 11940 35019 11996
rect 34955 11936 35019 11940
rect 5172 11452 5236 11456
rect 5172 11396 5176 11452
rect 5176 11396 5232 11452
rect 5232 11396 5236 11452
rect 5172 11392 5236 11396
rect 5252 11452 5316 11456
rect 5252 11396 5256 11452
rect 5256 11396 5312 11452
rect 5312 11396 5316 11452
rect 5252 11392 5316 11396
rect 5332 11452 5396 11456
rect 5332 11396 5336 11452
rect 5336 11396 5392 11452
rect 5392 11396 5396 11452
rect 5332 11392 5396 11396
rect 5412 11452 5476 11456
rect 5412 11396 5416 11452
rect 5416 11396 5472 11452
rect 5472 11396 5476 11452
rect 5412 11392 5476 11396
rect 13613 11452 13677 11456
rect 13613 11396 13617 11452
rect 13617 11396 13673 11452
rect 13673 11396 13677 11452
rect 13613 11392 13677 11396
rect 13693 11452 13757 11456
rect 13693 11396 13697 11452
rect 13697 11396 13753 11452
rect 13753 11396 13757 11452
rect 13693 11392 13757 11396
rect 13773 11452 13837 11456
rect 13773 11396 13777 11452
rect 13777 11396 13833 11452
rect 13833 11396 13837 11452
rect 13773 11392 13837 11396
rect 13853 11452 13917 11456
rect 13853 11396 13857 11452
rect 13857 11396 13913 11452
rect 13913 11396 13917 11452
rect 13853 11392 13917 11396
rect 22054 11452 22118 11456
rect 22054 11396 22058 11452
rect 22058 11396 22114 11452
rect 22114 11396 22118 11452
rect 22054 11392 22118 11396
rect 22134 11452 22198 11456
rect 22134 11396 22138 11452
rect 22138 11396 22194 11452
rect 22194 11396 22198 11452
rect 22134 11392 22198 11396
rect 22214 11452 22278 11456
rect 22214 11396 22218 11452
rect 22218 11396 22274 11452
rect 22274 11396 22278 11452
rect 22214 11392 22278 11396
rect 22294 11452 22358 11456
rect 22294 11396 22298 11452
rect 22298 11396 22354 11452
rect 22354 11396 22358 11452
rect 22294 11392 22358 11396
rect 30495 11452 30559 11456
rect 30495 11396 30499 11452
rect 30499 11396 30555 11452
rect 30555 11396 30559 11452
rect 30495 11392 30559 11396
rect 30575 11452 30639 11456
rect 30575 11396 30579 11452
rect 30579 11396 30635 11452
rect 30635 11396 30639 11452
rect 30575 11392 30639 11396
rect 30655 11452 30719 11456
rect 30655 11396 30659 11452
rect 30659 11396 30715 11452
rect 30715 11396 30719 11452
rect 30655 11392 30719 11396
rect 30735 11452 30799 11456
rect 30735 11396 30739 11452
rect 30739 11396 30795 11452
rect 30795 11396 30799 11452
rect 30735 11392 30799 11396
rect 9392 10908 9456 10912
rect 9392 10852 9396 10908
rect 9396 10852 9452 10908
rect 9452 10852 9456 10908
rect 9392 10848 9456 10852
rect 9472 10908 9536 10912
rect 9472 10852 9476 10908
rect 9476 10852 9532 10908
rect 9532 10852 9536 10908
rect 9472 10848 9536 10852
rect 9552 10908 9616 10912
rect 9552 10852 9556 10908
rect 9556 10852 9612 10908
rect 9612 10852 9616 10908
rect 9552 10848 9616 10852
rect 9632 10908 9696 10912
rect 9632 10852 9636 10908
rect 9636 10852 9692 10908
rect 9692 10852 9696 10908
rect 9632 10848 9696 10852
rect 17833 10908 17897 10912
rect 17833 10852 17837 10908
rect 17837 10852 17893 10908
rect 17893 10852 17897 10908
rect 17833 10848 17897 10852
rect 17913 10908 17977 10912
rect 17913 10852 17917 10908
rect 17917 10852 17973 10908
rect 17973 10852 17977 10908
rect 17913 10848 17977 10852
rect 17993 10908 18057 10912
rect 17993 10852 17997 10908
rect 17997 10852 18053 10908
rect 18053 10852 18057 10908
rect 17993 10848 18057 10852
rect 18073 10908 18137 10912
rect 18073 10852 18077 10908
rect 18077 10852 18133 10908
rect 18133 10852 18137 10908
rect 18073 10848 18137 10852
rect 26274 10908 26338 10912
rect 26274 10852 26278 10908
rect 26278 10852 26334 10908
rect 26334 10852 26338 10908
rect 26274 10848 26338 10852
rect 26354 10908 26418 10912
rect 26354 10852 26358 10908
rect 26358 10852 26414 10908
rect 26414 10852 26418 10908
rect 26354 10848 26418 10852
rect 26434 10908 26498 10912
rect 26434 10852 26438 10908
rect 26438 10852 26494 10908
rect 26494 10852 26498 10908
rect 26434 10848 26498 10852
rect 26514 10908 26578 10912
rect 26514 10852 26518 10908
rect 26518 10852 26574 10908
rect 26574 10852 26578 10908
rect 26514 10848 26578 10852
rect 34715 10908 34779 10912
rect 34715 10852 34719 10908
rect 34719 10852 34775 10908
rect 34775 10852 34779 10908
rect 34715 10848 34779 10852
rect 34795 10908 34859 10912
rect 34795 10852 34799 10908
rect 34799 10852 34855 10908
rect 34855 10852 34859 10908
rect 34795 10848 34859 10852
rect 34875 10908 34939 10912
rect 34875 10852 34879 10908
rect 34879 10852 34935 10908
rect 34935 10852 34939 10908
rect 34875 10848 34939 10852
rect 34955 10908 35019 10912
rect 34955 10852 34959 10908
rect 34959 10852 35015 10908
rect 35015 10852 35019 10908
rect 34955 10848 35019 10852
rect 5172 10364 5236 10368
rect 5172 10308 5176 10364
rect 5176 10308 5232 10364
rect 5232 10308 5236 10364
rect 5172 10304 5236 10308
rect 5252 10364 5316 10368
rect 5252 10308 5256 10364
rect 5256 10308 5312 10364
rect 5312 10308 5316 10364
rect 5252 10304 5316 10308
rect 5332 10364 5396 10368
rect 5332 10308 5336 10364
rect 5336 10308 5392 10364
rect 5392 10308 5396 10364
rect 5332 10304 5396 10308
rect 5412 10364 5476 10368
rect 5412 10308 5416 10364
rect 5416 10308 5472 10364
rect 5472 10308 5476 10364
rect 5412 10304 5476 10308
rect 13613 10364 13677 10368
rect 13613 10308 13617 10364
rect 13617 10308 13673 10364
rect 13673 10308 13677 10364
rect 13613 10304 13677 10308
rect 13693 10364 13757 10368
rect 13693 10308 13697 10364
rect 13697 10308 13753 10364
rect 13753 10308 13757 10364
rect 13693 10304 13757 10308
rect 13773 10364 13837 10368
rect 13773 10308 13777 10364
rect 13777 10308 13833 10364
rect 13833 10308 13837 10364
rect 13773 10304 13837 10308
rect 13853 10364 13917 10368
rect 13853 10308 13857 10364
rect 13857 10308 13913 10364
rect 13913 10308 13917 10364
rect 13853 10304 13917 10308
rect 22054 10364 22118 10368
rect 22054 10308 22058 10364
rect 22058 10308 22114 10364
rect 22114 10308 22118 10364
rect 22054 10304 22118 10308
rect 22134 10364 22198 10368
rect 22134 10308 22138 10364
rect 22138 10308 22194 10364
rect 22194 10308 22198 10364
rect 22134 10304 22198 10308
rect 22214 10364 22278 10368
rect 22214 10308 22218 10364
rect 22218 10308 22274 10364
rect 22274 10308 22278 10364
rect 22214 10304 22278 10308
rect 22294 10364 22358 10368
rect 22294 10308 22298 10364
rect 22298 10308 22354 10364
rect 22354 10308 22358 10364
rect 22294 10304 22358 10308
rect 30495 10364 30559 10368
rect 30495 10308 30499 10364
rect 30499 10308 30555 10364
rect 30555 10308 30559 10364
rect 30495 10304 30559 10308
rect 30575 10364 30639 10368
rect 30575 10308 30579 10364
rect 30579 10308 30635 10364
rect 30635 10308 30639 10364
rect 30575 10304 30639 10308
rect 30655 10364 30719 10368
rect 30655 10308 30659 10364
rect 30659 10308 30715 10364
rect 30715 10308 30719 10364
rect 30655 10304 30719 10308
rect 30735 10364 30799 10368
rect 30735 10308 30739 10364
rect 30739 10308 30795 10364
rect 30795 10308 30799 10364
rect 30735 10304 30799 10308
rect 9392 9820 9456 9824
rect 9392 9764 9396 9820
rect 9396 9764 9452 9820
rect 9452 9764 9456 9820
rect 9392 9760 9456 9764
rect 9472 9820 9536 9824
rect 9472 9764 9476 9820
rect 9476 9764 9532 9820
rect 9532 9764 9536 9820
rect 9472 9760 9536 9764
rect 9552 9820 9616 9824
rect 9552 9764 9556 9820
rect 9556 9764 9612 9820
rect 9612 9764 9616 9820
rect 9552 9760 9616 9764
rect 9632 9820 9696 9824
rect 9632 9764 9636 9820
rect 9636 9764 9692 9820
rect 9692 9764 9696 9820
rect 9632 9760 9696 9764
rect 17833 9820 17897 9824
rect 17833 9764 17837 9820
rect 17837 9764 17893 9820
rect 17893 9764 17897 9820
rect 17833 9760 17897 9764
rect 17913 9820 17977 9824
rect 17913 9764 17917 9820
rect 17917 9764 17973 9820
rect 17973 9764 17977 9820
rect 17913 9760 17977 9764
rect 17993 9820 18057 9824
rect 17993 9764 17997 9820
rect 17997 9764 18053 9820
rect 18053 9764 18057 9820
rect 17993 9760 18057 9764
rect 18073 9820 18137 9824
rect 18073 9764 18077 9820
rect 18077 9764 18133 9820
rect 18133 9764 18137 9820
rect 18073 9760 18137 9764
rect 26274 9820 26338 9824
rect 26274 9764 26278 9820
rect 26278 9764 26334 9820
rect 26334 9764 26338 9820
rect 26274 9760 26338 9764
rect 26354 9820 26418 9824
rect 26354 9764 26358 9820
rect 26358 9764 26414 9820
rect 26414 9764 26418 9820
rect 26354 9760 26418 9764
rect 26434 9820 26498 9824
rect 26434 9764 26438 9820
rect 26438 9764 26494 9820
rect 26494 9764 26498 9820
rect 26434 9760 26498 9764
rect 26514 9820 26578 9824
rect 26514 9764 26518 9820
rect 26518 9764 26574 9820
rect 26574 9764 26578 9820
rect 26514 9760 26578 9764
rect 34715 9820 34779 9824
rect 34715 9764 34719 9820
rect 34719 9764 34775 9820
rect 34775 9764 34779 9820
rect 34715 9760 34779 9764
rect 34795 9820 34859 9824
rect 34795 9764 34799 9820
rect 34799 9764 34855 9820
rect 34855 9764 34859 9820
rect 34795 9760 34859 9764
rect 34875 9820 34939 9824
rect 34875 9764 34879 9820
rect 34879 9764 34935 9820
rect 34935 9764 34939 9820
rect 34875 9760 34939 9764
rect 34955 9820 35019 9824
rect 34955 9764 34959 9820
rect 34959 9764 35015 9820
rect 35015 9764 35019 9820
rect 34955 9760 35019 9764
rect 5172 9276 5236 9280
rect 5172 9220 5176 9276
rect 5176 9220 5232 9276
rect 5232 9220 5236 9276
rect 5172 9216 5236 9220
rect 5252 9276 5316 9280
rect 5252 9220 5256 9276
rect 5256 9220 5312 9276
rect 5312 9220 5316 9276
rect 5252 9216 5316 9220
rect 5332 9276 5396 9280
rect 5332 9220 5336 9276
rect 5336 9220 5392 9276
rect 5392 9220 5396 9276
rect 5332 9216 5396 9220
rect 5412 9276 5476 9280
rect 5412 9220 5416 9276
rect 5416 9220 5472 9276
rect 5472 9220 5476 9276
rect 5412 9216 5476 9220
rect 13613 9276 13677 9280
rect 13613 9220 13617 9276
rect 13617 9220 13673 9276
rect 13673 9220 13677 9276
rect 13613 9216 13677 9220
rect 13693 9276 13757 9280
rect 13693 9220 13697 9276
rect 13697 9220 13753 9276
rect 13753 9220 13757 9276
rect 13693 9216 13757 9220
rect 13773 9276 13837 9280
rect 13773 9220 13777 9276
rect 13777 9220 13833 9276
rect 13833 9220 13837 9276
rect 13773 9216 13837 9220
rect 13853 9276 13917 9280
rect 13853 9220 13857 9276
rect 13857 9220 13913 9276
rect 13913 9220 13917 9276
rect 13853 9216 13917 9220
rect 22054 9276 22118 9280
rect 22054 9220 22058 9276
rect 22058 9220 22114 9276
rect 22114 9220 22118 9276
rect 22054 9216 22118 9220
rect 22134 9276 22198 9280
rect 22134 9220 22138 9276
rect 22138 9220 22194 9276
rect 22194 9220 22198 9276
rect 22134 9216 22198 9220
rect 22214 9276 22278 9280
rect 22214 9220 22218 9276
rect 22218 9220 22274 9276
rect 22274 9220 22278 9276
rect 22214 9216 22278 9220
rect 22294 9276 22358 9280
rect 22294 9220 22298 9276
rect 22298 9220 22354 9276
rect 22354 9220 22358 9276
rect 22294 9216 22358 9220
rect 30495 9276 30559 9280
rect 30495 9220 30499 9276
rect 30499 9220 30555 9276
rect 30555 9220 30559 9276
rect 30495 9216 30559 9220
rect 30575 9276 30639 9280
rect 30575 9220 30579 9276
rect 30579 9220 30635 9276
rect 30635 9220 30639 9276
rect 30575 9216 30639 9220
rect 30655 9276 30719 9280
rect 30655 9220 30659 9276
rect 30659 9220 30715 9276
rect 30715 9220 30719 9276
rect 30655 9216 30719 9220
rect 30735 9276 30799 9280
rect 30735 9220 30739 9276
rect 30739 9220 30795 9276
rect 30795 9220 30799 9276
rect 30735 9216 30799 9220
rect 9392 8732 9456 8736
rect 9392 8676 9396 8732
rect 9396 8676 9452 8732
rect 9452 8676 9456 8732
rect 9392 8672 9456 8676
rect 9472 8732 9536 8736
rect 9472 8676 9476 8732
rect 9476 8676 9532 8732
rect 9532 8676 9536 8732
rect 9472 8672 9536 8676
rect 9552 8732 9616 8736
rect 9552 8676 9556 8732
rect 9556 8676 9612 8732
rect 9612 8676 9616 8732
rect 9552 8672 9616 8676
rect 9632 8732 9696 8736
rect 9632 8676 9636 8732
rect 9636 8676 9692 8732
rect 9692 8676 9696 8732
rect 9632 8672 9696 8676
rect 17833 8732 17897 8736
rect 17833 8676 17837 8732
rect 17837 8676 17893 8732
rect 17893 8676 17897 8732
rect 17833 8672 17897 8676
rect 17913 8732 17977 8736
rect 17913 8676 17917 8732
rect 17917 8676 17973 8732
rect 17973 8676 17977 8732
rect 17913 8672 17977 8676
rect 17993 8732 18057 8736
rect 17993 8676 17997 8732
rect 17997 8676 18053 8732
rect 18053 8676 18057 8732
rect 17993 8672 18057 8676
rect 18073 8732 18137 8736
rect 18073 8676 18077 8732
rect 18077 8676 18133 8732
rect 18133 8676 18137 8732
rect 18073 8672 18137 8676
rect 26274 8732 26338 8736
rect 26274 8676 26278 8732
rect 26278 8676 26334 8732
rect 26334 8676 26338 8732
rect 26274 8672 26338 8676
rect 26354 8732 26418 8736
rect 26354 8676 26358 8732
rect 26358 8676 26414 8732
rect 26414 8676 26418 8732
rect 26354 8672 26418 8676
rect 26434 8732 26498 8736
rect 26434 8676 26438 8732
rect 26438 8676 26494 8732
rect 26494 8676 26498 8732
rect 26434 8672 26498 8676
rect 26514 8732 26578 8736
rect 26514 8676 26518 8732
rect 26518 8676 26574 8732
rect 26574 8676 26578 8732
rect 26514 8672 26578 8676
rect 34715 8732 34779 8736
rect 34715 8676 34719 8732
rect 34719 8676 34775 8732
rect 34775 8676 34779 8732
rect 34715 8672 34779 8676
rect 34795 8732 34859 8736
rect 34795 8676 34799 8732
rect 34799 8676 34855 8732
rect 34855 8676 34859 8732
rect 34795 8672 34859 8676
rect 34875 8732 34939 8736
rect 34875 8676 34879 8732
rect 34879 8676 34935 8732
rect 34935 8676 34939 8732
rect 34875 8672 34939 8676
rect 34955 8732 35019 8736
rect 34955 8676 34959 8732
rect 34959 8676 35015 8732
rect 35015 8676 35019 8732
rect 34955 8672 35019 8676
rect 5172 8188 5236 8192
rect 5172 8132 5176 8188
rect 5176 8132 5232 8188
rect 5232 8132 5236 8188
rect 5172 8128 5236 8132
rect 5252 8188 5316 8192
rect 5252 8132 5256 8188
rect 5256 8132 5312 8188
rect 5312 8132 5316 8188
rect 5252 8128 5316 8132
rect 5332 8188 5396 8192
rect 5332 8132 5336 8188
rect 5336 8132 5392 8188
rect 5392 8132 5396 8188
rect 5332 8128 5396 8132
rect 5412 8188 5476 8192
rect 5412 8132 5416 8188
rect 5416 8132 5472 8188
rect 5472 8132 5476 8188
rect 5412 8128 5476 8132
rect 13613 8188 13677 8192
rect 13613 8132 13617 8188
rect 13617 8132 13673 8188
rect 13673 8132 13677 8188
rect 13613 8128 13677 8132
rect 13693 8188 13757 8192
rect 13693 8132 13697 8188
rect 13697 8132 13753 8188
rect 13753 8132 13757 8188
rect 13693 8128 13757 8132
rect 13773 8188 13837 8192
rect 13773 8132 13777 8188
rect 13777 8132 13833 8188
rect 13833 8132 13837 8188
rect 13773 8128 13837 8132
rect 13853 8188 13917 8192
rect 13853 8132 13857 8188
rect 13857 8132 13913 8188
rect 13913 8132 13917 8188
rect 13853 8128 13917 8132
rect 22054 8188 22118 8192
rect 22054 8132 22058 8188
rect 22058 8132 22114 8188
rect 22114 8132 22118 8188
rect 22054 8128 22118 8132
rect 22134 8188 22198 8192
rect 22134 8132 22138 8188
rect 22138 8132 22194 8188
rect 22194 8132 22198 8188
rect 22134 8128 22198 8132
rect 22214 8188 22278 8192
rect 22214 8132 22218 8188
rect 22218 8132 22274 8188
rect 22274 8132 22278 8188
rect 22214 8128 22278 8132
rect 22294 8188 22358 8192
rect 22294 8132 22298 8188
rect 22298 8132 22354 8188
rect 22354 8132 22358 8188
rect 22294 8128 22358 8132
rect 30495 8188 30559 8192
rect 30495 8132 30499 8188
rect 30499 8132 30555 8188
rect 30555 8132 30559 8188
rect 30495 8128 30559 8132
rect 30575 8188 30639 8192
rect 30575 8132 30579 8188
rect 30579 8132 30635 8188
rect 30635 8132 30639 8188
rect 30575 8128 30639 8132
rect 30655 8188 30719 8192
rect 30655 8132 30659 8188
rect 30659 8132 30715 8188
rect 30715 8132 30719 8188
rect 30655 8128 30719 8132
rect 30735 8188 30799 8192
rect 30735 8132 30739 8188
rect 30739 8132 30795 8188
rect 30795 8132 30799 8188
rect 30735 8128 30799 8132
rect 9392 7644 9456 7648
rect 9392 7588 9396 7644
rect 9396 7588 9452 7644
rect 9452 7588 9456 7644
rect 9392 7584 9456 7588
rect 9472 7644 9536 7648
rect 9472 7588 9476 7644
rect 9476 7588 9532 7644
rect 9532 7588 9536 7644
rect 9472 7584 9536 7588
rect 9552 7644 9616 7648
rect 9552 7588 9556 7644
rect 9556 7588 9612 7644
rect 9612 7588 9616 7644
rect 9552 7584 9616 7588
rect 9632 7644 9696 7648
rect 9632 7588 9636 7644
rect 9636 7588 9692 7644
rect 9692 7588 9696 7644
rect 9632 7584 9696 7588
rect 17833 7644 17897 7648
rect 17833 7588 17837 7644
rect 17837 7588 17893 7644
rect 17893 7588 17897 7644
rect 17833 7584 17897 7588
rect 17913 7644 17977 7648
rect 17913 7588 17917 7644
rect 17917 7588 17973 7644
rect 17973 7588 17977 7644
rect 17913 7584 17977 7588
rect 17993 7644 18057 7648
rect 17993 7588 17997 7644
rect 17997 7588 18053 7644
rect 18053 7588 18057 7644
rect 17993 7584 18057 7588
rect 18073 7644 18137 7648
rect 18073 7588 18077 7644
rect 18077 7588 18133 7644
rect 18133 7588 18137 7644
rect 18073 7584 18137 7588
rect 26274 7644 26338 7648
rect 26274 7588 26278 7644
rect 26278 7588 26334 7644
rect 26334 7588 26338 7644
rect 26274 7584 26338 7588
rect 26354 7644 26418 7648
rect 26354 7588 26358 7644
rect 26358 7588 26414 7644
rect 26414 7588 26418 7644
rect 26354 7584 26418 7588
rect 26434 7644 26498 7648
rect 26434 7588 26438 7644
rect 26438 7588 26494 7644
rect 26494 7588 26498 7644
rect 26434 7584 26498 7588
rect 26514 7644 26578 7648
rect 26514 7588 26518 7644
rect 26518 7588 26574 7644
rect 26574 7588 26578 7644
rect 26514 7584 26578 7588
rect 34715 7644 34779 7648
rect 34715 7588 34719 7644
rect 34719 7588 34775 7644
rect 34775 7588 34779 7644
rect 34715 7584 34779 7588
rect 34795 7644 34859 7648
rect 34795 7588 34799 7644
rect 34799 7588 34855 7644
rect 34855 7588 34859 7644
rect 34795 7584 34859 7588
rect 34875 7644 34939 7648
rect 34875 7588 34879 7644
rect 34879 7588 34935 7644
rect 34935 7588 34939 7644
rect 34875 7584 34939 7588
rect 34955 7644 35019 7648
rect 34955 7588 34959 7644
rect 34959 7588 35015 7644
rect 35015 7588 35019 7644
rect 34955 7584 35019 7588
rect 5172 7100 5236 7104
rect 5172 7044 5176 7100
rect 5176 7044 5232 7100
rect 5232 7044 5236 7100
rect 5172 7040 5236 7044
rect 5252 7100 5316 7104
rect 5252 7044 5256 7100
rect 5256 7044 5312 7100
rect 5312 7044 5316 7100
rect 5252 7040 5316 7044
rect 5332 7100 5396 7104
rect 5332 7044 5336 7100
rect 5336 7044 5392 7100
rect 5392 7044 5396 7100
rect 5332 7040 5396 7044
rect 5412 7100 5476 7104
rect 5412 7044 5416 7100
rect 5416 7044 5472 7100
rect 5472 7044 5476 7100
rect 5412 7040 5476 7044
rect 13613 7100 13677 7104
rect 13613 7044 13617 7100
rect 13617 7044 13673 7100
rect 13673 7044 13677 7100
rect 13613 7040 13677 7044
rect 13693 7100 13757 7104
rect 13693 7044 13697 7100
rect 13697 7044 13753 7100
rect 13753 7044 13757 7100
rect 13693 7040 13757 7044
rect 13773 7100 13837 7104
rect 13773 7044 13777 7100
rect 13777 7044 13833 7100
rect 13833 7044 13837 7100
rect 13773 7040 13837 7044
rect 13853 7100 13917 7104
rect 13853 7044 13857 7100
rect 13857 7044 13913 7100
rect 13913 7044 13917 7100
rect 13853 7040 13917 7044
rect 22054 7100 22118 7104
rect 22054 7044 22058 7100
rect 22058 7044 22114 7100
rect 22114 7044 22118 7100
rect 22054 7040 22118 7044
rect 22134 7100 22198 7104
rect 22134 7044 22138 7100
rect 22138 7044 22194 7100
rect 22194 7044 22198 7100
rect 22134 7040 22198 7044
rect 22214 7100 22278 7104
rect 22214 7044 22218 7100
rect 22218 7044 22274 7100
rect 22274 7044 22278 7100
rect 22214 7040 22278 7044
rect 22294 7100 22358 7104
rect 22294 7044 22298 7100
rect 22298 7044 22354 7100
rect 22354 7044 22358 7100
rect 22294 7040 22358 7044
rect 30495 7100 30559 7104
rect 30495 7044 30499 7100
rect 30499 7044 30555 7100
rect 30555 7044 30559 7100
rect 30495 7040 30559 7044
rect 30575 7100 30639 7104
rect 30575 7044 30579 7100
rect 30579 7044 30635 7100
rect 30635 7044 30639 7100
rect 30575 7040 30639 7044
rect 30655 7100 30719 7104
rect 30655 7044 30659 7100
rect 30659 7044 30715 7100
rect 30715 7044 30719 7100
rect 30655 7040 30719 7044
rect 30735 7100 30799 7104
rect 30735 7044 30739 7100
rect 30739 7044 30795 7100
rect 30795 7044 30799 7100
rect 30735 7040 30799 7044
rect 9392 6556 9456 6560
rect 9392 6500 9396 6556
rect 9396 6500 9452 6556
rect 9452 6500 9456 6556
rect 9392 6496 9456 6500
rect 9472 6556 9536 6560
rect 9472 6500 9476 6556
rect 9476 6500 9532 6556
rect 9532 6500 9536 6556
rect 9472 6496 9536 6500
rect 9552 6556 9616 6560
rect 9552 6500 9556 6556
rect 9556 6500 9612 6556
rect 9612 6500 9616 6556
rect 9552 6496 9616 6500
rect 9632 6556 9696 6560
rect 9632 6500 9636 6556
rect 9636 6500 9692 6556
rect 9692 6500 9696 6556
rect 9632 6496 9696 6500
rect 17833 6556 17897 6560
rect 17833 6500 17837 6556
rect 17837 6500 17893 6556
rect 17893 6500 17897 6556
rect 17833 6496 17897 6500
rect 17913 6556 17977 6560
rect 17913 6500 17917 6556
rect 17917 6500 17973 6556
rect 17973 6500 17977 6556
rect 17913 6496 17977 6500
rect 17993 6556 18057 6560
rect 17993 6500 17997 6556
rect 17997 6500 18053 6556
rect 18053 6500 18057 6556
rect 17993 6496 18057 6500
rect 18073 6556 18137 6560
rect 18073 6500 18077 6556
rect 18077 6500 18133 6556
rect 18133 6500 18137 6556
rect 18073 6496 18137 6500
rect 26274 6556 26338 6560
rect 26274 6500 26278 6556
rect 26278 6500 26334 6556
rect 26334 6500 26338 6556
rect 26274 6496 26338 6500
rect 26354 6556 26418 6560
rect 26354 6500 26358 6556
rect 26358 6500 26414 6556
rect 26414 6500 26418 6556
rect 26354 6496 26418 6500
rect 26434 6556 26498 6560
rect 26434 6500 26438 6556
rect 26438 6500 26494 6556
rect 26494 6500 26498 6556
rect 26434 6496 26498 6500
rect 26514 6556 26578 6560
rect 26514 6500 26518 6556
rect 26518 6500 26574 6556
rect 26574 6500 26578 6556
rect 26514 6496 26578 6500
rect 34715 6556 34779 6560
rect 34715 6500 34719 6556
rect 34719 6500 34775 6556
rect 34775 6500 34779 6556
rect 34715 6496 34779 6500
rect 34795 6556 34859 6560
rect 34795 6500 34799 6556
rect 34799 6500 34855 6556
rect 34855 6500 34859 6556
rect 34795 6496 34859 6500
rect 34875 6556 34939 6560
rect 34875 6500 34879 6556
rect 34879 6500 34935 6556
rect 34935 6500 34939 6556
rect 34875 6496 34939 6500
rect 34955 6556 35019 6560
rect 34955 6500 34959 6556
rect 34959 6500 35015 6556
rect 35015 6500 35019 6556
rect 34955 6496 35019 6500
rect 5172 6012 5236 6016
rect 5172 5956 5176 6012
rect 5176 5956 5232 6012
rect 5232 5956 5236 6012
rect 5172 5952 5236 5956
rect 5252 6012 5316 6016
rect 5252 5956 5256 6012
rect 5256 5956 5312 6012
rect 5312 5956 5316 6012
rect 5252 5952 5316 5956
rect 5332 6012 5396 6016
rect 5332 5956 5336 6012
rect 5336 5956 5392 6012
rect 5392 5956 5396 6012
rect 5332 5952 5396 5956
rect 5412 6012 5476 6016
rect 5412 5956 5416 6012
rect 5416 5956 5472 6012
rect 5472 5956 5476 6012
rect 5412 5952 5476 5956
rect 13613 6012 13677 6016
rect 13613 5956 13617 6012
rect 13617 5956 13673 6012
rect 13673 5956 13677 6012
rect 13613 5952 13677 5956
rect 13693 6012 13757 6016
rect 13693 5956 13697 6012
rect 13697 5956 13753 6012
rect 13753 5956 13757 6012
rect 13693 5952 13757 5956
rect 13773 6012 13837 6016
rect 13773 5956 13777 6012
rect 13777 5956 13833 6012
rect 13833 5956 13837 6012
rect 13773 5952 13837 5956
rect 13853 6012 13917 6016
rect 13853 5956 13857 6012
rect 13857 5956 13913 6012
rect 13913 5956 13917 6012
rect 13853 5952 13917 5956
rect 22054 6012 22118 6016
rect 22054 5956 22058 6012
rect 22058 5956 22114 6012
rect 22114 5956 22118 6012
rect 22054 5952 22118 5956
rect 22134 6012 22198 6016
rect 22134 5956 22138 6012
rect 22138 5956 22194 6012
rect 22194 5956 22198 6012
rect 22134 5952 22198 5956
rect 22214 6012 22278 6016
rect 22214 5956 22218 6012
rect 22218 5956 22274 6012
rect 22274 5956 22278 6012
rect 22214 5952 22278 5956
rect 22294 6012 22358 6016
rect 22294 5956 22298 6012
rect 22298 5956 22354 6012
rect 22354 5956 22358 6012
rect 22294 5952 22358 5956
rect 30495 6012 30559 6016
rect 30495 5956 30499 6012
rect 30499 5956 30555 6012
rect 30555 5956 30559 6012
rect 30495 5952 30559 5956
rect 30575 6012 30639 6016
rect 30575 5956 30579 6012
rect 30579 5956 30635 6012
rect 30635 5956 30639 6012
rect 30575 5952 30639 5956
rect 30655 6012 30719 6016
rect 30655 5956 30659 6012
rect 30659 5956 30715 6012
rect 30715 5956 30719 6012
rect 30655 5952 30719 5956
rect 30735 6012 30799 6016
rect 30735 5956 30739 6012
rect 30739 5956 30795 6012
rect 30795 5956 30799 6012
rect 30735 5952 30799 5956
rect 9392 5468 9456 5472
rect 9392 5412 9396 5468
rect 9396 5412 9452 5468
rect 9452 5412 9456 5468
rect 9392 5408 9456 5412
rect 9472 5468 9536 5472
rect 9472 5412 9476 5468
rect 9476 5412 9532 5468
rect 9532 5412 9536 5468
rect 9472 5408 9536 5412
rect 9552 5468 9616 5472
rect 9552 5412 9556 5468
rect 9556 5412 9612 5468
rect 9612 5412 9616 5468
rect 9552 5408 9616 5412
rect 9632 5468 9696 5472
rect 9632 5412 9636 5468
rect 9636 5412 9692 5468
rect 9692 5412 9696 5468
rect 9632 5408 9696 5412
rect 17833 5468 17897 5472
rect 17833 5412 17837 5468
rect 17837 5412 17893 5468
rect 17893 5412 17897 5468
rect 17833 5408 17897 5412
rect 17913 5468 17977 5472
rect 17913 5412 17917 5468
rect 17917 5412 17973 5468
rect 17973 5412 17977 5468
rect 17913 5408 17977 5412
rect 17993 5468 18057 5472
rect 17993 5412 17997 5468
rect 17997 5412 18053 5468
rect 18053 5412 18057 5468
rect 17993 5408 18057 5412
rect 18073 5468 18137 5472
rect 18073 5412 18077 5468
rect 18077 5412 18133 5468
rect 18133 5412 18137 5468
rect 18073 5408 18137 5412
rect 26274 5468 26338 5472
rect 26274 5412 26278 5468
rect 26278 5412 26334 5468
rect 26334 5412 26338 5468
rect 26274 5408 26338 5412
rect 26354 5468 26418 5472
rect 26354 5412 26358 5468
rect 26358 5412 26414 5468
rect 26414 5412 26418 5468
rect 26354 5408 26418 5412
rect 26434 5468 26498 5472
rect 26434 5412 26438 5468
rect 26438 5412 26494 5468
rect 26494 5412 26498 5468
rect 26434 5408 26498 5412
rect 26514 5468 26578 5472
rect 26514 5412 26518 5468
rect 26518 5412 26574 5468
rect 26574 5412 26578 5468
rect 26514 5408 26578 5412
rect 34715 5468 34779 5472
rect 34715 5412 34719 5468
rect 34719 5412 34775 5468
rect 34775 5412 34779 5468
rect 34715 5408 34779 5412
rect 34795 5468 34859 5472
rect 34795 5412 34799 5468
rect 34799 5412 34855 5468
rect 34855 5412 34859 5468
rect 34795 5408 34859 5412
rect 34875 5468 34939 5472
rect 34875 5412 34879 5468
rect 34879 5412 34935 5468
rect 34935 5412 34939 5468
rect 34875 5408 34939 5412
rect 34955 5468 35019 5472
rect 34955 5412 34959 5468
rect 34959 5412 35015 5468
rect 35015 5412 35019 5468
rect 34955 5408 35019 5412
rect 5172 4924 5236 4928
rect 5172 4868 5176 4924
rect 5176 4868 5232 4924
rect 5232 4868 5236 4924
rect 5172 4864 5236 4868
rect 5252 4924 5316 4928
rect 5252 4868 5256 4924
rect 5256 4868 5312 4924
rect 5312 4868 5316 4924
rect 5252 4864 5316 4868
rect 5332 4924 5396 4928
rect 5332 4868 5336 4924
rect 5336 4868 5392 4924
rect 5392 4868 5396 4924
rect 5332 4864 5396 4868
rect 5412 4924 5476 4928
rect 5412 4868 5416 4924
rect 5416 4868 5472 4924
rect 5472 4868 5476 4924
rect 5412 4864 5476 4868
rect 13613 4924 13677 4928
rect 13613 4868 13617 4924
rect 13617 4868 13673 4924
rect 13673 4868 13677 4924
rect 13613 4864 13677 4868
rect 13693 4924 13757 4928
rect 13693 4868 13697 4924
rect 13697 4868 13753 4924
rect 13753 4868 13757 4924
rect 13693 4864 13757 4868
rect 13773 4924 13837 4928
rect 13773 4868 13777 4924
rect 13777 4868 13833 4924
rect 13833 4868 13837 4924
rect 13773 4864 13837 4868
rect 13853 4924 13917 4928
rect 13853 4868 13857 4924
rect 13857 4868 13913 4924
rect 13913 4868 13917 4924
rect 13853 4864 13917 4868
rect 22054 4924 22118 4928
rect 22054 4868 22058 4924
rect 22058 4868 22114 4924
rect 22114 4868 22118 4924
rect 22054 4864 22118 4868
rect 22134 4924 22198 4928
rect 22134 4868 22138 4924
rect 22138 4868 22194 4924
rect 22194 4868 22198 4924
rect 22134 4864 22198 4868
rect 22214 4924 22278 4928
rect 22214 4868 22218 4924
rect 22218 4868 22274 4924
rect 22274 4868 22278 4924
rect 22214 4864 22278 4868
rect 22294 4924 22358 4928
rect 22294 4868 22298 4924
rect 22298 4868 22354 4924
rect 22354 4868 22358 4924
rect 22294 4864 22358 4868
rect 30495 4924 30559 4928
rect 30495 4868 30499 4924
rect 30499 4868 30555 4924
rect 30555 4868 30559 4924
rect 30495 4864 30559 4868
rect 30575 4924 30639 4928
rect 30575 4868 30579 4924
rect 30579 4868 30635 4924
rect 30635 4868 30639 4924
rect 30575 4864 30639 4868
rect 30655 4924 30719 4928
rect 30655 4868 30659 4924
rect 30659 4868 30715 4924
rect 30715 4868 30719 4924
rect 30655 4864 30719 4868
rect 30735 4924 30799 4928
rect 30735 4868 30739 4924
rect 30739 4868 30795 4924
rect 30795 4868 30799 4924
rect 30735 4864 30799 4868
rect 9392 4380 9456 4384
rect 9392 4324 9396 4380
rect 9396 4324 9452 4380
rect 9452 4324 9456 4380
rect 9392 4320 9456 4324
rect 9472 4380 9536 4384
rect 9472 4324 9476 4380
rect 9476 4324 9532 4380
rect 9532 4324 9536 4380
rect 9472 4320 9536 4324
rect 9552 4380 9616 4384
rect 9552 4324 9556 4380
rect 9556 4324 9612 4380
rect 9612 4324 9616 4380
rect 9552 4320 9616 4324
rect 9632 4380 9696 4384
rect 9632 4324 9636 4380
rect 9636 4324 9692 4380
rect 9692 4324 9696 4380
rect 9632 4320 9696 4324
rect 17833 4380 17897 4384
rect 17833 4324 17837 4380
rect 17837 4324 17893 4380
rect 17893 4324 17897 4380
rect 17833 4320 17897 4324
rect 17913 4380 17977 4384
rect 17913 4324 17917 4380
rect 17917 4324 17973 4380
rect 17973 4324 17977 4380
rect 17913 4320 17977 4324
rect 17993 4380 18057 4384
rect 17993 4324 17997 4380
rect 17997 4324 18053 4380
rect 18053 4324 18057 4380
rect 17993 4320 18057 4324
rect 18073 4380 18137 4384
rect 18073 4324 18077 4380
rect 18077 4324 18133 4380
rect 18133 4324 18137 4380
rect 18073 4320 18137 4324
rect 26274 4380 26338 4384
rect 26274 4324 26278 4380
rect 26278 4324 26334 4380
rect 26334 4324 26338 4380
rect 26274 4320 26338 4324
rect 26354 4380 26418 4384
rect 26354 4324 26358 4380
rect 26358 4324 26414 4380
rect 26414 4324 26418 4380
rect 26354 4320 26418 4324
rect 26434 4380 26498 4384
rect 26434 4324 26438 4380
rect 26438 4324 26494 4380
rect 26494 4324 26498 4380
rect 26434 4320 26498 4324
rect 26514 4380 26578 4384
rect 26514 4324 26518 4380
rect 26518 4324 26574 4380
rect 26574 4324 26578 4380
rect 26514 4320 26578 4324
rect 34715 4380 34779 4384
rect 34715 4324 34719 4380
rect 34719 4324 34775 4380
rect 34775 4324 34779 4380
rect 34715 4320 34779 4324
rect 34795 4380 34859 4384
rect 34795 4324 34799 4380
rect 34799 4324 34855 4380
rect 34855 4324 34859 4380
rect 34795 4320 34859 4324
rect 34875 4380 34939 4384
rect 34875 4324 34879 4380
rect 34879 4324 34935 4380
rect 34935 4324 34939 4380
rect 34875 4320 34939 4324
rect 34955 4380 35019 4384
rect 34955 4324 34959 4380
rect 34959 4324 35015 4380
rect 35015 4324 35019 4380
rect 34955 4320 35019 4324
rect 5172 3836 5236 3840
rect 5172 3780 5176 3836
rect 5176 3780 5232 3836
rect 5232 3780 5236 3836
rect 5172 3776 5236 3780
rect 5252 3836 5316 3840
rect 5252 3780 5256 3836
rect 5256 3780 5312 3836
rect 5312 3780 5316 3836
rect 5252 3776 5316 3780
rect 5332 3836 5396 3840
rect 5332 3780 5336 3836
rect 5336 3780 5392 3836
rect 5392 3780 5396 3836
rect 5332 3776 5396 3780
rect 5412 3836 5476 3840
rect 5412 3780 5416 3836
rect 5416 3780 5472 3836
rect 5472 3780 5476 3836
rect 5412 3776 5476 3780
rect 13613 3836 13677 3840
rect 13613 3780 13617 3836
rect 13617 3780 13673 3836
rect 13673 3780 13677 3836
rect 13613 3776 13677 3780
rect 13693 3836 13757 3840
rect 13693 3780 13697 3836
rect 13697 3780 13753 3836
rect 13753 3780 13757 3836
rect 13693 3776 13757 3780
rect 13773 3836 13837 3840
rect 13773 3780 13777 3836
rect 13777 3780 13833 3836
rect 13833 3780 13837 3836
rect 13773 3776 13837 3780
rect 13853 3836 13917 3840
rect 13853 3780 13857 3836
rect 13857 3780 13913 3836
rect 13913 3780 13917 3836
rect 13853 3776 13917 3780
rect 22054 3836 22118 3840
rect 22054 3780 22058 3836
rect 22058 3780 22114 3836
rect 22114 3780 22118 3836
rect 22054 3776 22118 3780
rect 22134 3836 22198 3840
rect 22134 3780 22138 3836
rect 22138 3780 22194 3836
rect 22194 3780 22198 3836
rect 22134 3776 22198 3780
rect 22214 3836 22278 3840
rect 22214 3780 22218 3836
rect 22218 3780 22274 3836
rect 22274 3780 22278 3836
rect 22214 3776 22278 3780
rect 22294 3836 22358 3840
rect 22294 3780 22298 3836
rect 22298 3780 22354 3836
rect 22354 3780 22358 3836
rect 22294 3776 22358 3780
rect 30495 3836 30559 3840
rect 30495 3780 30499 3836
rect 30499 3780 30555 3836
rect 30555 3780 30559 3836
rect 30495 3776 30559 3780
rect 30575 3836 30639 3840
rect 30575 3780 30579 3836
rect 30579 3780 30635 3836
rect 30635 3780 30639 3836
rect 30575 3776 30639 3780
rect 30655 3836 30719 3840
rect 30655 3780 30659 3836
rect 30659 3780 30715 3836
rect 30715 3780 30719 3836
rect 30655 3776 30719 3780
rect 30735 3836 30799 3840
rect 30735 3780 30739 3836
rect 30739 3780 30795 3836
rect 30795 3780 30799 3836
rect 30735 3776 30799 3780
rect 9392 3292 9456 3296
rect 9392 3236 9396 3292
rect 9396 3236 9452 3292
rect 9452 3236 9456 3292
rect 9392 3232 9456 3236
rect 9472 3292 9536 3296
rect 9472 3236 9476 3292
rect 9476 3236 9532 3292
rect 9532 3236 9536 3292
rect 9472 3232 9536 3236
rect 9552 3292 9616 3296
rect 9552 3236 9556 3292
rect 9556 3236 9612 3292
rect 9612 3236 9616 3292
rect 9552 3232 9616 3236
rect 9632 3292 9696 3296
rect 9632 3236 9636 3292
rect 9636 3236 9692 3292
rect 9692 3236 9696 3292
rect 9632 3232 9696 3236
rect 17833 3292 17897 3296
rect 17833 3236 17837 3292
rect 17837 3236 17893 3292
rect 17893 3236 17897 3292
rect 17833 3232 17897 3236
rect 17913 3292 17977 3296
rect 17913 3236 17917 3292
rect 17917 3236 17973 3292
rect 17973 3236 17977 3292
rect 17913 3232 17977 3236
rect 17993 3292 18057 3296
rect 17993 3236 17997 3292
rect 17997 3236 18053 3292
rect 18053 3236 18057 3292
rect 17993 3232 18057 3236
rect 18073 3292 18137 3296
rect 18073 3236 18077 3292
rect 18077 3236 18133 3292
rect 18133 3236 18137 3292
rect 18073 3232 18137 3236
rect 26274 3292 26338 3296
rect 26274 3236 26278 3292
rect 26278 3236 26334 3292
rect 26334 3236 26338 3292
rect 26274 3232 26338 3236
rect 26354 3292 26418 3296
rect 26354 3236 26358 3292
rect 26358 3236 26414 3292
rect 26414 3236 26418 3292
rect 26354 3232 26418 3236
rect 26434 3292 26498 3296
rect 26434 3236 26438 3292
rect 26438 3236 26494 3292
rect 26494 3236 26498 3292
rect 26434 3232 26498 3236
rect 26514 3292 26578 3296
rect 26514 3236 26518 3292
rect 26518 3236 26574 3292
rect 26574 3236 26578 3292
rect 26514 3232 26578 3236
rect 34715 3292 34779 3296
rect 34715 3236 34719 3292
rect 34719 3236 34775 3292
rect 34775 3236 34779 3292
rect 34715 3232 34779 3236
rect 34795 3292 34859 3296
rect 34795 3236 34799 3292
rect 34799 3236 34855 3292
rect 34855 3236 34859 3292
rect 34795 3232 34859 3236
rect 34875 3292 34939 3296
rect 34875 3236 34879 3292
rect 34879 3236 34935 3292
rect 34935 3236 34939 3292
rect 34875 3232 34939 3236
rect 34955 3292 35019 3296
rect 34955 3236 34959 3292
rect 34959 3236 35015 3292
rect 35015 3236 35019 3292
rect 34955 3232 35019 3236
rect 5172 2748 5236 2752
rect 5172 2692 5176 2748
rect 5176 2692 5232 2748
rect 5232 2692 5236 2748
rect 5172 2688 5236 2692
rect 5252 2748 5316 2752
rect 5252 2692 5256 2748
rect 5256 2692 5312 2748
rect 5312 2692 5316 2748
rect 5252 2688 5316 2692
rect 5332 2748 5396 2752
rect 5332 2692 5336 2748
rect 5336 2692 5392 2748
rect 5392 2692 5396 2748
rect 5332 2688 5396 2692
rect 5412 2748 5476 2752
rect 5412 2692 5416 2748
rect 5416 2692 5472 2748
rect 5472 2692 5476 2748
rect 5412 2688 5476 2692
rect 13613 2748 13677 2752
rect 13613 2692 13617 2748
rect 13617 2692 13673 2748
rect 13673 2692 13677 2748
rect 13613 2688 13677 2692
rect 13693 2748 13757 2752
rect 13693 2692 13697 2748
rect 13697 2692 13753 2748
rect 13753 2692 13757 2748
rect 13693 2688 13757 2692
rect 13773 2748 13837 2752
rect 13773 2692 13777 2748
rect 13777 2692 13833 2748
rect 13833 2692 13837 2748
rect 13773 2688 13837 2692
rect 13853 2748 13917 2752
rect 13853 2692 13857 2748
rect 13857 2692 13913 2748
rect 13913 2692 13917 2748
rect 13853 2688 13917 2692
rect 22054 2748 22118 2752
rect 22054 2692 22058 2748
rect 22058 2692 22114 2748
rect 22114 2692 22118 2748
rect 22054 2688 22118 2692
rect 22134 2748 22198 2752
rect 22134 2692 22138 2748
rect 22138 2692 22194 2748
rect 22194 2692 22198 2748
rect 22134 2688 22198 2692
rect 22214 2748 22278 2752
rect 22214 2692 22218 2748
rect 22218 2692 22274 2748
rect 22274 2692 22278 2748
rect 22214 2688 22278 2692
rect 22294 2748 22358 2752
rect 22294 2692 22298 2748
rect 22298 2692 22354 2748
rect 22354 2692 22358 2748
rect 22294 2688 22358 2692
rect 30495 2748 30559 2752
rect 30495 2692 30499 2748
rect 30499 2692 30555 2748
rect 30555 2692 30559 2748
rect 30495 2688 30559 2692
rect 30575 2748 30639 2752
rect 30575 2692 30579 2748
rect 30579 2692 30635 2748
rect 30635 2692 30639 2748
rect 30575 2688 30639 2692
rect 30655 2748 30719 2752
rect 30655 2692 30659 2748
rect 30659 2692 30715 2748
rect 30715 2692 30719 2748
rect 30655 2688 30719 2692
rect 30735 2748 30799 2752
rect 30735 2692 30739 2748
rect 30739 2692 30795 2748
rect 30795 2692 30799 2748
rect 30735 2688 30799 2692
rect 9392 2204 9456 2208
rect 9392 2148 9396 2204
rect 9396 2148 9452 2204
rect 9452 2148 9456 2204
rect 9392 2144 9456 2148
rect 9472 2204 9536 2208
rect 9472 2148 9476 2204
rect 9476 2148 9532 2204
rect 9532 2148 9536 2204
rect 9472 2144 9536 2148
rect 9552 2204 9616 2208
rect 9552 2148 9556 2204
rect 9556 2148 9612 2204
rect 9612 2148 9616 2204
rect 9552 2144 9616 2148
rect 9632 2204 9696 2208
rect 9632 2148 9636 2204
rect 9636 2148 9692 2204
rect 9692 2148 9696 2204
rect 9632 2144 9696 2148
rect 17833 2204 17897 2208
rect 17833 2148 17837 2204
rect 17837 2148 17893 2204
rect 17893 2148 17897 2204
rect 17833 2144 17897 2148
rect 17913 2204 17977 2208
rect 17913 2148 17917 2204
rect 17917 2148 17973 2204
rect 17973 2148 17977 2204
rect 17913 2144 17977 2148
rect 17993 2204 18057 2208
rect 17993 2148 17997 2204
rect 17997 2148 18053 2204
rect 18053 2148 18057 2204
rect 17993 2144 18057 2148
rect 18073 2204 18137 2208
rect 18073 2148 18077 2204
rect 18077 2148 18133 2204
rect 18133 2148 18137 2204
rect 18073 2144 18137 2148
rect 26274 2204 26338 2208
rect 26274 2148 26278 2204
rect 26278 2148 26334 2204
rect 26334 2148 26338 2204
rect 26274 2144 26338 2148
rect 26354 2204 26418 2208
rect 26354 2148 26358 2204
rect 26358 2148 26414 2204
rect 26414 2148 26418 2204
rect 26354 2144 26418 2148
rect 26434 2204 26498 2208
rect 26434 2148 26438 2204
rect 26438 2148 26494 2204
rect 26494 2148 26498 2204
rect 26434 2144 26498 2148
rect 26514 2204 26578 2208
rect 26514 2148 26518 2204
rect 26518 2148 26574 2204
rect 26574 2148 26578 2204
rect 26514 2144 26578 2148
rect 34715 2204 34779 2208
rect 34715 2148 34719 2204
rect 34719 2148 34775 2204
rect 34775 2148 34779 2204
rect 34715 2144 34779 2148
rect 34795 2204 34859 2208
rect 34795 2148 34799 2204
rect 34799 2148 34855 2204
rect 34855 2148 34859 2204
rect 34795 2144 34859 2148
rect 34875 2204 34939 2208
rect 34875 2148 34879 2204
rect 34879 2148 34935 2204
rect 34935 2148 34939 2204
rect 34875 2144 34939 2148
rect 34955 2204 35019 2208
rect 34955 2148 34959 2204
rect 34959 2148 35015 2204
rect 35015 2148 35019 2204
rect 34955 2144 35019 2148
<< metal4 >>
rect 5164 33216 5484 33776
rect 5164 33152 5172 33216
rect 5236 33152 5252 33216
rect 5316 33152 5332 33216
rect 5396 33152 5412 33216
rect 5476 33152 5484 33216
rect 5164 32128 5484 33152
rect 5164 32064 5172 32128
rect 5236 32064 5252 32128
rect 5316 32064 5332 32128
rect 5396 32064 5412 32128
rect 5476 32064 5484 32128
rect 5164 31040 5484 32064
rect 5164 30976 5172 31040
rect 5236 30976 5252 31040
rect 5316 30976 5332 31040
rect 5396 30976 5412 31040
rect 5476 30976 5484 31040
rect 5164 29952 5484 30976
rect 5164 29888 5172 29952
rect 5236 29888 5252 29952
rect 5316 29888 5332 29952
rect 5396 29888 5412 29952
rect 5476 29888 5484 29952
rect 5164 28864 5484 29888
rect 5164 28800 5172 28864
rect 5236 28800 5252 28864
rect 5316 28800 5332 28864
rect 5396 28800 5412 28864
rect 5476 28800 5484 28864
rect 5164 27776 5484 28800
rect 5164 27712 5172 27776
rect 5236 27712 5252 27776
rect 5316 27712 5332 27776
rect 5396 27712 5412 27776
rect 5476 27712 5484 27776
rect 5164 26688 5484 27712
rect 5164 26624 5172 26688
rect 5236 26624 5252 26688
rect 5316 26624 5332 26688
rect 5396 26624 5412 26688
rect 5476 26624 5484 26688
rect 5164 25600 5484 26624
rect 5164 25536 5172 25600
rect 5236 25536 5252 25600
rect 5316 25536 5332 25600
rect 5396 25536 5412 25600
rect 5476 25536 5484 25600
rect 5164 24512 5484 25536
rect 5164 24448 5172 24512
rect 5236 24448 5252 24512
rect 5316 24448 5332 24512
rect 5396 24448 5412 24512
rect 5476 24448 5484 24512
rect 5164 23424 5484 24448
rect 5164 23360 5172 23424
rect 5236 23360 5252 23424
rect 5316 23360 5332 23424
rect 5396 23360 5412 23424
rect 5476 23360 5484 23424
rect 5164 22336 5484 23360
rect 5164 22272 5172 22336
rect 5236 22272 5252 22336
rect 5316 22272 5332 22336
rect 5396 22272 5412 22336
rect 5476 22272 5484 22336
rect 5164 21248 5484 22272
rect 5164 21184 5172 21248
rect 5236 21184 5252 21248
rect 5316 21184 5332 21248
rect 5396 21184 5412 21248
rect 5476 21184 5484 21248
rect 5164 20160 5484 21184
rect 5164 20096 5172 20160
rect 5236 20096 5252 20160
rect 5316 20096 5332 20160
rect 5396 20096 5412 20160
rect 5476 20096 5484 20160
rect 5164 19072 5484 20096
rect 5164 19008 5172 19072
rect 5236 19008 5252 19072
rect 5316 19008 5332 19072
rect 5396 19008 5412 19072
rect 5476 19008 5484 19072
rect 5164 17984 5484 19008
rect 5164 17920 5172 17984
rect 5236 17920 5252 17984
rect 5316 17920 5332 17984
rect 5396 17920 5412 17984
rect 5476 17920 5484 17984
rect 5164 16896 5484 17920
rect 5164 16832 5172 16896
rect 5236 16832 5252 16896
rect 5316 16832 5332 16896
rect 5396 16832 5412 16896
rect 5476 16832 5484 16896
rect 5164 15808 5484 16832
rect 5164 15744 5172 15808
rect 5236 15744 5252 15808
rect 5316 15744 5332 15808
rect 5396 15744 5412 15808
rect 5476 15744 5484 15808
rect 5164 14720 5484 15744
rect 5164 14656 5172 14720
rect 5236 14656 5252 14720
rect 5316 14656 5332 14720
rect 5396 14656 5412 14720
rect 5476 14656 5484 14720
rect 5164 13632 5484 14656
rect 5164 13568 5172 13632
rect 5236 13568 5252 13632
rect 5316 13568 5332 13632
rect 5396 13568 5412 13632
rect 5476 13568 5484 13632
rect 5164 12544 5484 13568
rect 5164 12480 5172 12544
rect 5236 12480 5252 12544
rect 5316 12480 5332 12544
rect 5396 12480 5412 12544
rect 5476 12480 5484 12544
rect 5164 11456 5484 12480
rect 5164 11392 5172 11456
rect 5236 11392 5252 11456
rect 5316 11392 5332 11456
rect 5396 11392 5412 11456
rect 5476 11392 5484 11456
rect 5164 10368 5484 11392
rect 5164 10304 5172 10368
rect 5236 10304 5252 10368
rect 5316 10304 5332 10368
rect 5396 10304 5412 10368
rect 5476 10304 5484 10368
rect 5164 9280 5484 10304
rect 5164 9216 5172 9280
rect 5236 9216 5252 9280
rect 5316 9216 5332 9280
rect 5396 9216 5412 9280
rect 5476 9216 5484 9280
rect 5164 8192 5484 9216
rect 5164 8128 5172 8192
rect 5236 8128 5252 8192
rect 5316 8128 5332 8192
rect 5396 8128 5412 8192
rect 5476 8128 5484 8192
rect 5164 7104 5484 8128
rect 5164 7040 5172 7104
rect 5236 7040 5252 7104
rect 5316 7040 5332 7104
rect 5396 7040 5412 7104
rect 5476 7040 5484 7104
rect 5164 6016 5484 7040
rect 5164 5952 5172 6016
rect 5236 5952 5252 6016
rect 5316 5952 5332 6016
rect 5396 5952 5412 6016
rect 5476 5952 5484 6016
rect 5164 4928 5484 5952
rect 5164 4864 5172 4928
rect 5236 4864 5252 4928
rect 5316 4864 5332 4928
rect 5396 4864 5412 4928
rect 5476 4864 5484 4928
rect 5164 3840 5484 4864
rect 5164 3776 5172 3840
rect 5236 3776 5252 3840
rect 5316 3776 5332 3840
rect 5396 3776 5412 3840
rect 5476 3776 5484 3840
rect 5164 2752 5484 3776
rect 5164 2688 5172 2752
rect 5236 2688 5252 2752
rect 5316 2688 5332 2752
rect 5396 2688 5412 2752
rect 5476 2688 5484 2752
rect 5164 2128 5484 2688
rect 9384 33760 9704 33776
rect 9384 33696 9392 33760
rect 9456 33696 9472 33760
rect 9536 33696 9552 33760
rect 9616 33696 9632 33760
rect 9696 33696 9704 33760
rect 9384 32672 9704 33696
rect 9384 32608 9392 32672
rect 9456 32608 9472 32672
rect 9536 32608 9552 32672
rect 9616 32608 9632 32672
rect 9696 32608 9704 32672
rect 9384 31584 9704 32608
rect 9384 31520 9392 31584
rect 9456 31520 9472 31584
rect 9536 31520 9552 31584
rect 9616 31520 9632 31584
rect 9696 31520 9704 31584
rect 9384 30496 9704 31520
rect 9384 30432 9392 30496
rect 9456 30432 9472 30496
rect 9536 30432 9552 30496
rect 9616 30432 9632 30496
rect 9696 30432 9704 30496
rect 9384 29408 9704 30432
rect 9384 29344 9392 29408
rect 9456 29344 9472 29408
rect 9536 29344 9552 29408
rect 9616 29344 9632 29408
rect 9696 29344 9704 29408
rect 9384 28320 9704 29344
rect 9384 28256 9392 28320
rect 9456 28256 9472 28320
rect 9536 28256 9552 28320
rect 9616 28256 9632 28320
rect 9696 28256 9704 28320
rect 9384 27232 9704 28256
rect 9384 27168 9392 27232
rect 9456 27168 9472 27232
rect 9536 27168 9552 27232
rect 9616 27168 9632 27232
rect 9696 27168 9704 27232
rect 9384 26144 9704 27168
rect 9384 26080 9392 26144
rect 9456 26080 9472 26144
rect 9536 26080 9552 26144
rect 9616 26080 9632 26144
rect 9696 26080 9704 26144
rect 9384 25056 9704 26080
rect 9384 24992 9392 25056
rect 9456 24992 9472 25056
rect 9536 24992 9552 25056
rect 9616 24992 9632 25056
rect 9696 24992 9704 25056
rect 9384 23968 9704 24992
rect 9384 23904 9392 23968
rect 9456 23904 9472 23968
rect 9536 23904 9552 23968
rect 9616 23904 9632 23968
rect 9696 23904 9704 23968
rect 9384 22880 9704 23904
rect 9384 22816 9392 22880
rect 9456 22816 9472 22880
rect 9536 22816 9552 22880
rect 9616 22816 9632 22880
rect 9696 22816 9704 22880
rect 9384 21792 9704 22816
rect 9384 21728 9392 21792
rect 9456 21728 9472 21792
rect 9536 21728 9552 21792
rect 9616 21728 9632 21792
rect 9696 21728 9704 21792
rect 9384 20704 9704 21728
rect 9384 20640 9392 20704
rect 9456 20640 9472 20704
rect 9536 20640 9552 20704
rect 9616 20640 9632 20704
rect 9696 20640 9704 20704
rect 9384 19616 9704 20640
rect 9384 19552 9392 19616
rect 9456 19552 9472 19616
rect 9536 19552 9552 19616
rect 9616 19552 9632 19616
rect 9696 19552 9704 19616
rect 9384 18528 9704 19552
rect 9384 18464 9392 18528
rect 9456 18464 9472 18528
rect 9536 18464 9552 18528
rect 9616 18464 9632 18528
rect 9696 18464 9704 18528
rect 9384 17440 9704 18464
rect 9384 17376 9392 17440
rect 9456 17376 9472 17440
rect 9536 17376 9552 17440
rect 9616 17376 9632 17440
rect 9696 17376 9704 17440
rect 9384 16352 9704 17376
rect 9384 16288 9392 16352
rect 9456 16288 9472 16352
rect 9536 16288 9552 16352
rect 9616 16288 9632 16352
rect 9696 16288 9704 16352
rect 9384 15264 9704 16288
rect 9384 15200 9392 15264
rect 9456 15200 9472 15264
rect 9536 15200 9552 15264
rect 9616 15200 9632 15264
rect 9696 15200 9704 15264
rect 9384 14176 9704 15200
rect 9384 14112 9392 14176
rect 9456 14112 9472 14176
rect 9536 14112 9552 14176
rect 9616 14112 9632 14176
rect 9696 14112 9704 14176
rect 9384 13088 9704 14112
rect 9384 13024 9392 13088
rect 9456 13024 9472 13088
rect 9536 13024 9552 13088
rect 9616 13024 9632 13088
rect 9696 13024 9704 13088
rect 9384 12000 9704 13024
rect 9384 11936 9392 12000
rect 9456 11936 9472 12000
rect 9536 11936 9552 12000
rect 9616 11936 9632 12000
rect 9696 11936 9704 12000
rect 9384 10912 9704 11936
rect 9384 10848 9392 10912
rect 9456 10848 9472 10912
rect 9536 10848 9552 10912
rect 9616 10848 9632 10912
rect 9696 10848 9704 10912
rect 9384 9824 9704 10848
rect 9384 9760 9392 9824
rect 9456 9760 9472 9824
rect 9536 9760 9552 9824
rect 9616 9760 9632 9824
rect 9696 9760 9704 9824
rect 9384 8736 9704 9760
rect 9384 8672 9392 8736
rect 9456 8672 9472 8736
rect 9536 8672 9552 8736
rect 9616 8672 9632 8736
rect 9696 8672 9704 8736
rect 9384 7648 9704 8672
rect 9384 7584 9392 7648
rect 9456 7584 9472 7648
rect 9536 7584 9552 7648
rect 9616 7584 9632 7648
rect 9696 7584 9704 7648
rect 9384 6560 9704 7584
rect 9384 6496 9392 6560
rect 9456 6496 9472 6560
rect 9536 6496 9552 6560
rect 9616 6496 9632 6560
rect 9696 6496 9704 6560
rect 9384 5472 9704 6496
rect 9384 5408 9392 5472
rect 9456 5408 9472 5472
rect 9536 5408 9552 5472
rect 9616 5408 9632 5472
rect 9696 5408 9704 5472
rect 9384 4384 9704 5408
rect 9384 4320 9392 4384
rect 9456 4320 9472 4384
rect 9536 4320 9552 4384
rect 9616 4320 9632 4384
rect 9696 4320 9704 4384
rect 9384 3296 9704 4320
rect 9384 3232 9392 3296
rect 9456 3232 9472 3296
rect 9536 3232 9552 3296
rect 9616 3232 9632 3296
rect 9696 3232 9704 3296
rect 9384 2208 9704 3232
rect 9384 2144 9392 2208
rect 9456 2144 9472 2208
rect 9536 2144 9552 2208
rect 9616 2144 9632 2208
rect 9696 2144 9704 2208
rect 9384 2128 9704 2144
rect 13605 33216 13925 33776
rect 13605 33152 13613 33216
rect 13677 33152 13693 33216
rect 13757 33152 13773 33216
rect 13837 33152 13853 33216
rect 13917 33152 13925 33216
rect 13605 32128 13925 33152
rect 13605 32064 13613 32128
rect 13677 32064 13693 32128
rect 13757 32064 13773 32128
rect 13837 32064 13853 32128
rect 13917 32064 13925 32128
rect 13605 31040 13925 32064
rect 13605 30976 13613 31040
rect 13677 30976 13693 31040
rect 13757 30976 13773 31040
rect 13837 30976 13853 31040
rect 13917 30976 13925 31040
rect 13605 29952 13925 30976
rect 13605 29888 13613 29952
rect 13677 29888 13693 29952
rect 13757 29888 13773 29952
rect 13837 29888 13853 29952
rect 13917 29888 13925 29952
rect 13605 28864 13925 29888
rect 13605 28800 13613 28864
rect 13677 28800 13693 28864
rect 13757 28800 13773 28864
rect 13837 28800 13853 28864
rect 13917 28800 13925 28864
rect 13605 27776 13925 28800
rect 13605 27712 13613 27776
rect 13677 27712 13693 27776
rect 13757 27712 13773 27776
rect 13837 27712 13853 27776
rect 13917 27712 13925 27776
rect 13605 26688 13925 27712
rect 13605 26624 13613 26688
rect 13677 26624 13693 26688
rect 13757 26624 13773 26688
rect 13837 26624 13853 26688
rect 13917 26624 13925 26688
rect 13605 25600 13925 26624
rect 13605 25536 13613 25600
rect 13677 25536 13693 25600
rect 13757 25536 13773 25600
rect 13837 25536 13853 25600
rect 13917 25536 13925 25600
rect 13605 24512 13925 25536
rect 13605 24448 13613 24512
rect 13677 24448 13693 24512
rect 13757 24448 13773 24512
rect 13837 24448 13853 24512
rect 13917 24448 13925 24512
rect 13605 23424 13925 24448
rect 13605 23360 13613 23424
rect 13677 23360 13693 23424
rect 13757 23360 13773 23424
rect 13837 23360 13853 23424
rect 13917 23360 13925 23424
rect 13605 22336 13925 23360
rect 13605 22272 13613 22336
rect 13677 22272 13693 22336
rect 13757 22272 13773 22336
rect 13837 22272 13853 22336
rect 13917 22272 13925 22336
rect 13605 21248 13925 22272
rect 13605 21184 13613 21248
rect 13677 21184 13693 21248
rect 13757 21184 13773 21248
rect 13837 21184 13853 21248
rect 13917 21184 13925 21248
rect 13605 20160 13925 21184
rect 13605 20096 13613 20160
rect 13677 20096 13693 20160
rect 13757 20096 13773 20160
rect 13837 20096 13853 20160
rect 13917 20096 13925 20160
rect 13605 19072 13925 20096
rect 13605 19008 13613 19072
rect 13677 19008 13693 19072
rect 13757 19008 13773 19072
rect 13837 19008 13853 19072
rect 13917 19008 13925 19072
rect 13605 17984 13925 19008
rect 13605 17920 13613 17984
rect 13677 17920 13693 17984
rect 13757 17920 13773 17984
rect 13837 17920 13853 17984
rect 13917 17920 13925 17984
rect 13605 16896 13925 17920
rect 13605 16832 13613 16896
rect 13677 16832 13693 16896
rect 13757 16832 13773 16896
rect 13837 16832 13853 16896
rect 13917 16832 13925 16896
rect 13605 15808 13925 16832
rect 13605 15744 13613 15808
rect 13677 15744 13693 15808
rect 13757 15744 13773 15808
rect 13837 15744 13853 15808
rect 13917 15744 13925 15808
rect 13605 14720 13925 15744
rect 13605 14656 13613 14720
rect 13677 14656 13693 14720
rect 13757 14656 13773 14720
rect 13837 14656 13853 14720
rect 13917 14656 13925 14720
rect 13605 13632 13925 14656
rect 13605 13568 13613 13632
rect 13677 13568 13693 13632
rect 13757 13568 13773 13632
rect 13837 13568 13853 13632
rect 13917 13568 13925 13632
rect 13605 12544 13925 13568
rect 13605 12480 13613 12544
rect 13677 12480 13693 12544
rect 13757 12480 13773 12544
rect 13837 12480 13853 12544
rect 13917 12480 13925 12544
rect 13605 11456 13925 12480
rect 13605 11392 13613 11456
rect 13677 11392 13693 11456
rect 13757 11392 13773 11456
rect 13837 11392 13853 11456
rect 13917 11392 13925 11456
rect 13605 10368 13925 11392
rect 13605 10304 13613 10368
rect 13677 10304 13693 10368
rect 13757 10304 13773 10368
rect 13837 10304 13853 10368
rect 13917 10304 13925 10368
rect 13605 9280 13925 10304
rect 13605 9216 13613 9280
rect 13677 9216 13693 9280
rect 13757 9216 13773 9280
rect 13837 9216 13853 9280
rect 13917 9216 13925 9280
rect 13605 8192 13925 9216
rect 13605 8128 13613 8192
rect 13677 8128 13693 8192
rect 13757 8128 13773 8192
rect 13837 8128 13853 8192
rect 13917 8128 13925 8192
rect 13605 7104 13925 8128
rect 13605 7040 13613 7104
rect 13677 7040 13693 7104
rect 13757 7040 13773 7104
rect 13837 7040 13853 7104
rect 13917 7040 13925 7104
rect 13605 6016 13925 7040
rect 13605 5952 13613 6016
rect 13677 5952 13693 6016
rect 13757 5952 13773 6016
rect 13837 5952 13853 6016
rect 13917 5952 13925 6016
rect 13605 4928 13925 5952
rect 13605 4864 13613 4928
rect 13677 4864 13693 4928
rect 13757 4864 13773 4928
rect 13837 4864 13853 4928
rect 13917 4864 13925 4928
rect 13605 3840 13925 4864
rect 13605 3776 13613 3840
rect 13677 3776 13693 3840
rect 13757 3776 13773 3840
rect 13837 3776 13853 3840
rect 13917 3776 13925 3840
rect 13605 2752 13925 3776
rect 13605 2688 13613 2752
rect 13677 2688 13693 2752
rect 13757 2688 13773 2752
rect 13837 2688 13853 2752
rect 13917 2688 13925 2752
rect 13605 2128 13925 2688
rect 17825 33760 18145 33776
rect 17825 33696 17833 33760
rect 17897 33696 17913 33760
rect 17977 33696 17993 33760
rect 18057 33696 18073 33760
rect 18137 33696 18145 33760
rect 17825 32672 18145 33696
rect 17825 32608 17833 32672
rect 17897 32608 17913 32672
rect 17977 32608 17993 32672
rect 18057 32608 18073 32672
rect 18137 32608 18145 32672
rect 17825 31584 18145 32608
rect 17825 31520 17833 31584
rect 17897 31520 17913 31584
rect 17977 31520 17993 31584
rect 18057 31520 18073 31584
rect 18137 31520 18145 31584
rect 17825 30496 18145 31520
rect 17825 30432 17833 30496
rect 17897 30432 17913 30496
rect 17977 30432 17993 30496
rect 18057 30432 18073 30496
rect 18137 30432 18145 30496
rect 17825 29408 18145 30432
rect 17825 29344 17833 29408
rect 17897 29344 17913 29408
rect 17977 29344 17993 29408
rect 18057 29344 18073 29408
rect 18137 29344 18145 29408
rect 17825 28320 18145 29344
rect 17825 28256 17833 28320
rect 17897 28256 17913 28320
rect 17977 28256 17993 28320
rect 18057 28256 18073 28320
rect 18137 28256 18145 28320
rect 17825 27232 18145 28256
rect 17825 27168 17833 27232
rect 17897 27168 17913 27232
rect 17977 27168 17993 27232
rect 18057 27168 18073 27232
rect 18137 27168 18145 27232
rect 17825 26144 18145 27168
rect 17825 26080 17833 26144
rect 17897 26080 17913 26144
rect 17977 26080 17993 26144
rect 18057 26080 18073 26144
rect 18137 26080 18145 26144
rect 17825 25056 18145 26080
rect 17825 24992 17833 25056
rect 17897 24992 17913 25056
rect 17977 24992 17993 25056
rect 18057 24992 18073 25056
rect 18137 24992 18145 25056
rect 17825 23968 18145 24992
rect 17825 23904 17833 23968
rect 17897 23904 17913 23968
rect 17977 23904 17993 23968
rect 18057 23904 18073 23968
rect 18137 23904 18145 23968
rect 17825 22880 18145 23904
rect 17825 22816 17833 22880
rect 17897 22816 17913 22880
rect 17977 22816 17993 22880
rect 18057 22816 18073 22880
rect 18137 22816 18145 22880
rect 17825 21792 18145 22816
rect 17825 21728 17833 21792
rect 17897 21728 17913 21792
rect 17977 21728 17993 21792
rect 18057 21728 18073 21792
rect 18137 21728 18145 21792
rect 17825 20704 18145 21728
rect 17825 20640 17833 20704
rect 17897 20640 17913 20704
rect 17977 20640 17993 20704
rect 18057 20640 18073 20704
rect 18137 20640 18145 20704
rect 17825 19616 18145 20640
rect 17825 19552 17833 19616
rect 17897 19552 17913 19616
rect 17977 19552 17993 19616
rect 18057 19552 18073 19616
rect 18137 19552 18145 19616
rect 17825 18528 18145 19552
rect 17825 18464 17833 18528
rect 17897 18464 17913 18528
rect 17977 18464 17993 18528
rect 18057 18464 18073 18528
rect 18137 18464 18145 18528
rect 17825 17440 18145 18464
rect 17825 17376 17833 17440
rect 17897 17376 17913 17440
rect 17977 17376 17993 17440
rect 18057 17376 18073 17440
rect 18137 17376 18145 17440
rect 17825 16352 18145 17376
rect 17825 16288 17833 16352
rect 17897 16288 17913 16352
rect 17977 16288 17993 16352
rect 18057 16288 18073 16352
rect 18137 16288 18145 16352
rect 17825 15264 18145 16288
rect 17825 15200 17833 15264
rect 17897 15200 17913 15264
rect 17977 15200 17993 15264
rect 18057 15200 18073 15264
rect 18137 15200 18145 15264
rect 17825 14176 18145 15200
rect 17825 14112 17833 14176
rect 17897 14112 17913 14176
rect 17977 14112 17993 14176
rect 18057 14112 18073 14176
rect 18137 14112 18145 14176
rect 17825 13088 18145 14112
rect 17825 13024 17833 13088
rect 17897 13024 17913 13088
rect 17977 13024 17993 13088
rect 18057 13024 18073 13088
rect 18137 13024 18145 13088
rect 17825 12000 18145 13024
rect 17825 11936 17833 12000
rect 17897 11936 17913 12000
rect 17977 11936 17993 12000
rect 18057 11936 18073 12000
rect 18137 11936 18145 12000
rect 17825 10912 18145 11936
rect 17825 10848 17833 10912
rect 17897 10848 17913 10912
rect 17977 10848 17993 10912
rect 18057 10848 18073 10912
rect 18137 10848 18145 10912
rect 17825 9824 18145 10848
rect 17825 9760 17833 9824
rect 17897 9760 17913 9824
rect 17977 9760 17993 9824
rect 18057 9760 18073 9824
rect 18137 9760 18145 9824
rect 17825 8736 18145 9760
rect 17825 8672 17833 8736
rect 17897 8672 17913 8736
rect 17977 8672 17993 8736
rect 18057 8672 18073 8736
rect 18137 8672 18145 8736
rect 17825 7648 18145 8672
rect 17825 7584 17833 7648
rect 17897 7584 17913 7648
rect 17977 7584 17993 7648
rect 18057 7584 18073 7648
rect 18137 7584 18145 7648
rect 17825 6560 18145 7584
rect 17825 6496 17833 6560
rect 17897 6496 17913 6560
rect 17977 6496 17993 6560
rect 18057 6496 18073 6560
rect 18137 6496 18145 6560
rect 17825 5472 18145 6496
rect 17825 5408 17833 5472
rect 17897 5408 17913 5472
rect 17977 5408 17993 5472
rect 18057 5408 18073 5472
rect 18137 5408 18145 5472
rect 17825 4384 18145 5408
rect 17825 4320 17833 4384
rect 17897 4320 17913 4384
rect 17977 4320 17993 4384
rect 18057 4320 18073 4384
rect 18137 4320 18145 4384
rect 17825 3296 18145 4320
rect 17825 3232 17833 3296
rect 17897 3232 17913 3296
rect 17977 3232 17993 3296
rect 18057 3232 18073 3296
rect 18137 3232 18145 3296
rect 17825 2208 18145 3232
rect 17825 2144 17833 2208
rect 17897 2144 17913 2208
rect 17977 2144 17993 2208
rect 18057 2144 18073 2208
rect 18137 2144 18145 2208
rect 17825 2128 18145 2144
rect 22046 33216 22366 33776
rect 22046 33152 22054 33216
rect 22118 33152 22134 33216
rect 22198 33152 22214 33216
rect 22278 33152 22294 33216
rect 22358 33152 22366 33216
rect 22046 32128 22366 33152
rect 22046 32064 22054 32128
rect 22118 32064 22134 32128
rect 22198 32064 22214 32128
rect 22278 32064 22294 32128
rect 22358 32064 22366 32128
rect 22046 31040 22366 32064
rect 22046 30976 22054 31040
rect 22118 30976 22134 31040
rect 22198 30976 22214 31040
rect 22278 30976 22294 31040
rect 22358 30976 22366 31040
rect 22046 29952 22366 30976
rect 22046 29888 22054 29952
rect 22118 29888 22134 29952
rect 22198 29888 22214 29952
rect 22278 29888 22294 29952
rect 22358 29888 22366 29952
rect 22046 28864 22366 29888
rect 22046 28800 22054 28864
rect 22118 28800 22134 28864
rect 22198 28800 22214 28864
rect 22278 28800 22294 28864
rect 22358 28800 22366 28864
rect 22046 27776 22366 28800
rect 22046 27712 22054 27776
rect 22118 27712 22134 27776
rect 22198 27712 22214 27776
rect 22278 27712 22294 27776
rect 22358 27712 22366 27776
rect 22046 26688 22366 27712
rect 22046 26624 22054 26688
rect 22118 26624 22134 26688
rect 22198 26624 22214 26688
rect 22278 26624 22294 26688
rect 22358 26624 22366 26688
rect 22046 25600 22366 26624
rect 22046 25536 22054 25600
rect 22118 25536 22134 25600
rect 22198 25536 22214 25600
rect 22278 25536 22294 25600
rect 22358 25536 22366 25600
rect 22046 24512 22366 25536
rect 22046 24448 22054 24512
rect 22118 24448 22134 24512
rect 22198 24448 22214 24512
rect 22278 24448 22294 24512
rect 22358 24448 22366 24512
rect 22046 23424 22366 24448
rect 22046 23360 22054 23424
rect 22118 23360 22134 23424
rect 22198 23360 22214 23424
rect 22278 23360 22294 23424
rect 22358 23360 22366 23424
rect 22046 22336 22366 23360
rect 22046 22272 22054 22336
rect 22118 22272 22134 22336
rect 22198 22272 22214 22336
rect 22278 22272 22294 22336
rect 22358 22272 22366 22336
rect 22046 21248 22366 22272
rect 22046 21184 22054 21248
rect 22118 21184 22134 21248
rect 22198 21184 22214 21248
rect 22278 21184 22294 21248
rect 22358 21184 22366 21248
rect 22046 20160 22366 21184
rect 22046 20096 22054 20160
rect 22118 20096 22134 20160
rect 22198 20096 22214 20160
rect 22278 20096 22294 20160
rect 22358 20096 22366 20160
rect 22046 19072 22366 20096
rect 22046 19008 22054 19072
rect 22118 19008 22134 19072
rect 22198 19008 22214 19072
rect 22278 19008 22294 19072
rect 22358 19008 22366 19072
rect 22046 17984 22366 19008
rect 22046 17920 22054 17984
rect 22118 17920 22134 17984
rect 22198 17920 22214 17984
rect 22278 17920 22294 17984
rect 22358 17920 22366 17984
rect 22046 16896 22366 17920
rect 22046 16832 22054 16896
rect 22118 16832 22134 16896
rect 22198 16832 22214 16896
rect 22278 16832 22294 16896
rect 22358 16832 22366 16896
rect 22046 15808 22366 16832
rect 22046 15744 22054 15808
rect 22118 15744 22134 15808
rect 22198 15744 22214 15808
rect 22278 15744 22294 15808
rect 22358 15744 22366 15808
rect 22046 14720 22366 15744
rect 22046 14656 22054 14720
rect 22118 14656 22134 14720
rect 22198 14656 22214 14720
rect 22278 14656 22294 14720
rect 22358 14656 22366 14720
rect 22046 13632 22366 14656
rect 22046 13568 22054 13632
rect 22118 13568 22134 13632
rect 22198 13568 22214 13632
rect 22278 13568 22294 13632
rect 22358 13568 22366 13632
rect 22046 12544 22366 13568
rect 22046 12480 22054 12544
rect 22118 12480 22134 12544
rect 22198 12480 22214 12544
rect 22278 12480 22294 12544
rect 22358 12480 22366 12544
rect 22046 11456 22366 12480
rect 22046 11392 22054 11456
rect 22118 11392 22134 11456
rect 22198 11392 22214 11456
rect 22278 11392 22294 11456
rect 22358 11392 22366 11456
rect 22046 10368 22366 11392
rect 22046 10304 22054 10368
rect 22118 10304 22134 10368
rect 22198 10304 22214 10368
rect 22278 10304 22294 10368
rect 22358 10304 22366 10368
rect 22046 9280 22366 10304
rect 22046 9216 22054 9280
rect 22118 9216 22134 9280
rect 22198 9216 22214 9280
rect 22278 9216 22294 9280
rect 22358 9216 22366 9280
rect 22046 8192 22366 9216
rect 22046 8128 22054 8192
rect 22118 8128 22134 8192
rect 22198 8128 22214 8192
rect 22278 8128 22294 8192
rect 22358 8128 22366 8192
rect 22046 7104 22366 8128
rect 22046 7040 22054 7104
rect 22118 7040 22134 7104
rect 22198 7040 22214 7104
rect 22278 7040 22294 7104
rect 22358 7040 22366 7104
rect 22046 6016 22366 7040
rect 22046 5952 22054 6016
rect 22118 5952 22134 6016
rect 22198 5952 22214 6016
rect 22278 5952 22294 6016
rect 22358 5952 22366 6016
rect 22046 4928 22366 5952
rect 22046 4864 22054 4928
rect 22118 4864 22134 4928
rect 22198 4864 22214 4928
rect 22278 4864 22294 4928
rect 22358 4864 22366 4928
rect 22046 3840 22366 4864
rect 22046 3776 22054 3840
rect 22118 3776 22134 3840
rect 22198 3776 22214 3840
rect 22278 3776 22294 3840
rect 22358 3776 22366 3840
rect 22046 2752 22366 3776
rect 22046 2688 22054 2752
rect 22118 2688 22134 2752
rect 22198 2688 22214 2752
rect 22278 2688 22294 2752
rect 22358 2688 22366 2752
rect 22046 2128 22366 2688
rect 26266 33760 26586 33776
rect 26266 33696 26274 33760
rect 26338 33696 26354 33760
rect 26418 33696 26434 33760
rect 26498 33696 26514 33760
rect 26578 33696 26586 33760
rect 26266 32672 26586 33696
rect 26266 32608 26274 32672
rect 26338 32608 26354 32672
rect 26418 32608 26434 32672
rect 26498 32608 26514 32672
rect 26578 32608 26586 32672
rect 26266 31584 26586 32608
rect 26266 31520 26274 31584
rect 26338 31520 26354 31584
rect 26418 31520 26434 31584
rect 26498 31520 26514 31584
rect 26578 31520 26586 31584
rect 26266 30496 26586 31520
rect 26266 30432 26274 30496
rect 26338 30432 26354 30496
rect 26418 30432 26434 30496
rect 26498 30432 26514 30496
rect 26578 30432 26586 30496
rect 26266 29408 26586 30432
rect 26266 29344 26274 29408
rect 26338 29344 26354 29408
rect 26418 29344 26434 29408
rect 26498 29344 26514 29408
rect 26578 29344 26586 29408
rect 26266 28320 26586 29344
rect 26266 28256 26274 28320
rect 26338 28256 26354 28320
rect 26418 28256 26434 28320
rect 26498 28256 26514 28320
rect 26578 28256 26586 28320
rect 26266 27232 26586 28256
rect 26266 27168 26274 27232
rect 26338 27168 26354 27232
rect 26418 27168 26434 27232
rect 26498 27168 26514 27232
rect 26578 27168 26586 27232
rect 26266 26144 26586 27168
rect 26266 26080 26274 26144
rect 26338 26080 26354 26144
rect 26418 26080 26434 26144
rect 26498 26080 26514 26144
rect 26578 26080 26586 26144
rect 26266 25056 26586 26080
rect 26266 24992 26274 25056
rect 26338 24992 26354 25056
rect 26418 24992 26434 25056
rect 26498 24992 26514 25056
rect 26578 24992 26586 25056
rect 26266 23968 26586 24992
rect 26266 23904 26274 23968
rect 26338 23904 26354 23968
rect 26418 23904 26434 23968
rect 26498 23904 26514 23968
rect 26578 23904 26586 23968
rect 26266 22880 26586 23904
rect 26266 22816 26274 22880
rect 26338 22816 26354 22880
rect 26418 22816 26434 22880
rect 26498 22816 26514 22880
rect 26578 22816 26586 22880
rect 26266 21792 26586 22816
rect 26266 21728 26274 21792
rect 26338 21728 26354 21792
rect 26418 21728 26434 21792
rect 26498 21728 26514 21792
rect 26578 21728 26586 21792
rect 26266 20704 26586 21728
rect 26266 20640 26274 20704
rect 26338 20640 26354 20704
rect 26418 20640 26434 20704
rect 26498 20640 26514 20704
rect 26578 20640 26586 20704
rect 26266 19616 26586 20640
rect 26266 19552 26274 19616
rect 26338 19552 26354 19616
rect 26418 19552 26434 19616
rect 26498 19552 26514 19616
rect 26578 19552 26586 19616
rect 26266 18528 26586 19552
rect 26266 18464 26274 18528
rect 26338 18464 26354 18528
rect 26418 18464 26434 18528
rect 26498 18464 26514 18528
rect 26578 18464 26586 18528
rect 26266 17440 26586 18464
rect 26266 17376 26274 17440
rect 26338 17376 26354 17440
rect 26418 17376 26434 17440
rect 26498 17376 26514 17440
rect 26578 17376 26586 17440
rect 26266 16352 26586 17376
rect 26266 16288 26274 16352
rect 26338 16288 26354 16352
rect 26418 16288 26434 16352
rect 26498 16288 26514 16352
rect 26578 16288 26586 16352
rect 26266 15264 26586 16288
rect 26266 15200 26274 15264
rect 26338 15200 26354 15264
rect 26418 15200 26434 15264
rect 26498 15200 26514 15264
rect 26578 15200 26586 15264
rect 26266 14176 26586 15200
rect 26266 14112 26274 14176
rect 26338 14112 26354 14176
rect 26418 14112 26434 14176
rect 26498 14112 26514 14176
rect 26578 14112 26586 14176
rect 26266 13088 26586 14112
rect 26266 13024 26274 13088
rect 26338 13024 26354 13088
rect 26418 13024 26434 13088
rect 26498 13024 26514 13088
rect 26578 13024 26586 13088
rect 26266 12000 26586 13024
rect 26266 11936 26274 12000
rect 26338 11936 26354 12000
rect 26418 11936 26434 12000
rect 26498 11936 26514 12000
rect 26578 11936 26586 12000
rect 26266 10912 26586 11936
rect 26266 10848 26274 10912
rect 26338 10848 26354 10912
rect 26418 10848 26434 10912
rect 26498 10848 26514 10912
rect 26578 10848 26586 10912
rect 26266 9824 26586 10848
rect 26266 9760 26274 9824
rect 26338 9760 26354 9824
rect 26418 9760 26434 9824
rect 26498 9760 26514 9824
rect 26578 9760 26586 9824
rect 26266 8736 26586 9760
rect 26266 8672 26274 8736
rect 26338 8672 26354 8736
rect 26418 8672 26434 8736
rect 26498 8672 26514 8736
rect 26578 8672 26586 8736
rect 26266 7648 26586 8672
rect 26266 7584 26274 7648
rect 26338 7584 26354 7648
rect 26418 7584 26434 7648
rect 26498 7584 26514 7648
rect 26578 7584 26586 7648
rect 26266 6560 26586 7584
rect 26266 6496 26274 6560
rect 26338 6496 26354 6560
rect 26418 6496 26434 6560
rect 26498 6496 26514 6560
rect 26578 6496 26586 6560
rect 26266 5472 26586 6496
rect 26266 5408 26274 5472
rect 26338 5408 26354 5472
rect 26418 5408 26434 5472
rect 26498 5408 26514 5472
rect 26578 5408 26586 5472
rect 26266 4384 26586 5408
rect 26266 4320 26274 4384
rect 26338 4320 26354 4384
rect 26418 4320 26434 4384
rect 26498 4320 26514 4384
rect 26578 4320 26586 4384
rect 26266 3296 26586 4320
rect 26266 3232 26274 3296
rect 26338 3232 26354 3296
rect 26418 3232 26434 3296
rect 26498 3232 26514 3296
rect 26578 3232 26586 3296
rect 26266 2208 26586 3232
rect 26266 2144 26274 2208
rect 26338 2144 26354 2208
rect 26418 2144 26434 2208
rect 26498 2144 26514 2208
rect 26578 2144 26586 2208
rect 26266 2128 26586 2144
rect 30487 33216 30807 33776
rect 30487 33152 30495 33216
rect 30559 33152 30575 33216
rect 30639 33152 30655 33216
rect 30719 33152 30735 33216
rect 30799 33152 30807 33216
rect 30487 32128 30807 33152
rect 30487 32064 30495 32128
rect 30559 32064 30575 32128
rect 30639 32064 30655 32128
rect 30719 32064 30735 32128
rect 30799 32064 30807 32128
rect 30487 31040 30807 32064
rect 30487 30976 30495 31040
rect 30559 30976 30575 31040
rect 30639 30976 30655 31040
rect 30719 30976 30735 31040
rect 30799 30976 30807 31040
rect 30487 29952 30807 30976
rect 30487 29888 30495 29952
rect 30559 29888 30575 29952
rect 30639 29888 30655 29952
rect 30719 29888 30735 29952
rect 30799 29888 30807 29952
rect 30487 28864 30807 29888
rect 30487 28800 30495 28864
rect 30559 28800 30575 28864
rect 30639 28800 30655 28864
rect 30719 28800 30735 28864
rect 30799 28800 30807 28864
rect 30487 27776 30807 28800
rect 30487 27712 30495 27776
rect 30559 27712 30575 27776
rect 30639 27712 30655 27776
rect 30719 27712 30735 27776
rect 30799 27712 30807 27776
rect 30487 26688 30807 27712
rect 30487 26624 30495 26688
rect 30559 26624 30575 26688
rect 30639 26624 30655 26688
rect 30719 26624 30735 26688
rect 30799 26624 30807 26688
rect 30487 25600 30807 26624
rect 30487 25536 30495 25600
rect 30559 25536 30575 25600
rect 30639 25536 30655 25600
rect 30719 25536 30735 25600
rect 30799 25536 30807 25600
rect 30487 24512 30807 25536
rect 30487 24448 30495 24512
rect 30559 24448 30575 24512
rect 30639 24448 30655 24512
rect 30719 24448 30735 24512
rect 30799 24448 30807 24512
rect 30487 23424 30807 24448
rect 30487 23360 30495 23424
rect 30559 23360 30575 23424
rect 30639 23360 30655 23424
rect 30719 23360 30735 23424
rect 30799 23360 30807 23424
rect 30487 22336 30807 23360
rect 30487 22272 30495 22336
rect 30559 22272 30575 22336
rect 30639 22272 30655 22336
rect 30719 22272 30735 22336
rect 30799 22272 30807 22336
rect 30487 21248 30807 22272
rect 30487 21184 30495 21248
rect 30559 21184 30575 21248
rect 30639 21184 30655 21248
rect 30719 21184 30735 21248
rect 30799 21184 30807 21248
rect 30487 20160 30807 21184
rect 30487 20096 30495 20160
rect 30559 20096 30575 20160
rect 30639 20096 30655 20160
rect 30719 20096 30735 20160
rect 30799 20096 30807 20160
rect 30487 19072 30807 20096
rect 30487 19008 30495 19072
rect 30559 19008 30575 19072
rect 30639 19008 30655 19072
rect 30719 19008 30735 19072
rect 30799 19008 30807 19072
rect 30487 17984 30807 19008
rect 30487 17920 30495 17984
rect 30559 17920 30575 17984
rect 30639 17920 30655 17984
rect 30719 17920 30735 17984
rect 30799 17920 30807 17984
rect 30487 16896 30807 17920
rect 30487 16832 30495 16896
rect 30559 16832 30575 16896
rect 30639 16832 30655 16896
rect 30719 16832 30735 16896
rect 30799 16832 30807 16896
rect 30487 15808 30807 16832
rect 30487 15744 30495 15808
rect 30559 15744 30575 15808
rect 30639 15744 30655 15808
rect 30719 15744 30735 15808
rect 30799 15744 30807 15808
rect 30487 14720 30807 15744
rect 30487 14656 30495 14720
rect 30559 14656 30575 14720
rect 30639 14656 30655 14720
rect 30719 14656 30735 14720
rect 30799 14656 30807 14720
rect 30487 13632 30807 14656
rect 30487 13568 30495 13632
rect 30559 13568 30575 13632
rect 30639 13568 30655 13632
rect 30719 13568 30735 13632
rect 30799 13568 30807 13632
rect 30487 12544 30807 13568
rect 30487 12480 30495 12544
rect 30559 12480 30575 12544
rect 30639 12480 30655 12544
rect 30719 12480 30735 12544
rect 30799 12480 30807 12544
rect 30487 11456 30807 12480
rect 30487 11392 30495 11456
rect 30559 11392 30575 11456
rect 30639 11392 30655 11456
rect 30719 11392 30735 11456
rect 30799 11392 30807 11456
rect 30487 10368 30807 11392
rect 30487 10304 30495 10368
rect 30559 10304 30575 10368
rect 30639 10304 30655 10368
rect 30719 10304 30735 10368
rect 30799 10304 30807 10368
rect 30487 9280 30807 10304
rect 30487 9216 30495 9280
rect 30559 9216 30575 9280
rect 30639 9216 30655 9280
rect 30719 9216 30735 9280
rect 30799 9216 30807 9280
rect 30487 8192 30807 9216
rect 30487 8128 30495 8192
rect 30559 8128 30575 8192
rect 30639 8128 30655 8192
rect 30719 8128 30735 8192
rect 30799 8128 30807 8192
rect 30487 7104 30807 8128
rect 30487 7040 30495 7104
rect 30559 7040 30575 7104
rect 30639 7040 30655 7104
rect 30719 7040 30735 7104
rect 30799 7040 30807 7104
rect 30487 6016 30807 7040
rect 30487 5952 30495 6016
rect 30559 5952 30575 6016
rect 30639 5952 30655 6016
rect 30719 5952 30735 6016
rect 30799 5952 30807 6016
rect 30487 4928 30807 5952
rect 30487 4864 30495 4928
rect 30559 4864 30575 4928
rect 30639 4864 30655 4928
rect 30719 4864 30735 4928
rect 30799 4864 30807 4928
rect 30487 3840 30807 4864
rect 30487 3776 30495 3840
rect 30559 3776 30575 3840
rect 30639 3776 30655 3840
rect 30719 3776 30735 3840
rect 30799 3776 30807 3840
rect 30487 2752 30807 3776
rect 30487 2688 30495 2752
rect 30559 2688 30575 2752
rect 30639 2688 30655 2752
rect 30719 2688 30735 2752
rect 30799 2688 30807 2752
rect 30487 2128 30807 2688
rect 34707 33760 35027 33776
rect 34707 33696 34715 33760
rect 34779 33696 34795 33760
rect 34859 33696 34875 33760
rect 34939 33696 34955 33760
rect 35019 33696 35027 33760
rect 34707 32672 35027 33696
rect 34707 32608 34715 32672
rect 34779 32608 34795 32672
rect 34859 32608 34875 32672
rect 34939 32608 34955 32672
rect 35019 32608 35027 32672
rect 34707 31584 35027 32608
rect 34707 31520 34715 31584
rect 34779 31520 34795 31584
rect 34859 31520 34875 31584
rect 34939 31520 34955 31584
rect 35019 31520 35027 31584
rect 34707 30496 35027 31520
rect 34707 30432 34715 30496
rect 34779 30432 34795 30496
rect 34859 30432 34875 30496
rect 34939 30432 34955 30496
rect 35019 30432 35027 30496
rect 34707 29408 35027 30432
rect 34707 29344 34715 29408
rect 34779 29344 34795 29408
rect 34859 29344 34875 29408
rect 34939 29344 34955 29408
rect 35019 29344 35027 29408
rect 34707 28320 35027 29344
rect 34707 28256 34715 28320
rect 34779 28256 34795 28320
rect 34859 28256 34875 28320
rect 34939 28256 34955 28320
rect 35019 28256 35027 28320
rect 34707 27232 35027 28256
rect 34707 27168 34715 27232
rect 34779 27168 34795 27232
rect 34859 27168 34875 27232
rect 34939 27168 34955 27232
rect 35019 27168 35027 27232
rect 34707 26144 35027 27168
rect 34707 26080 34715 26144
rect 34779 26080 34795 26144
rect 34859 26080 34875 26144
rect 34939 26080 34955 26144
rect 35019 26080 35027 26144
rect 34707 25056 35027 26080
rect 34707 24992 34715 25056
rect 34779 24992 34795 25056
rect 34859 24992 34875 25056
rect 34939 24992 34955 25056
rect 35019 24992 35027 25056
rect 34707 23968 35027 24992
rect 34707 23904 34715 23968
rect 34779 23904 34795 23968
rect 34859 23904 34875 23968
rect 34939 23904 34955 23968
rect 35019 23904 35027 23968
rect 34707 22880 35027 23904
rect 34707 22816 34715 22880
rect 34779 22816 34795 22880
rect 34859 22816 34875 22880
rect 34939 22816 34955 22880
rect 35019 22816 35027 22880
rect 34707 21792 35027 22816
rect 34707 21728 34715 21792
rect 34779 21728 34795 21792
rect 34859 21728 34875 21792
rect 34939 21728 34955 21792
rect 35019 21728 35027 21792
rect 34707 20704 35027 21728
rect 34707 20640 34715 20704
rect 34779 20640 34795 20704
rect 34859 20640 34875 20704
rect 34939 20640 34955 20704
rect 35019 20640 35027 20704
rect 34707 19616 35027 20640
rect 34707 19552 34715 19616
rect 34779 19552 34795 19616
rect 34859 19552 34875 19616
rect 34939 19552 34955 19616
rect 35019 19552 35027 19616
rect 34707 18528 35027 19552
rect 34707 18464 34715 18528
rect 34779 18464 34795 18528
rect 34859 18464 34875 18528
rect 34939 18464 34955 18528
rect 35019 18464 35027 18528
rect 34707 17440 35027 18464
rect 34707 17376 34715 17440
rect 34779 17376 34795 17440
rect 34859 17376 34875 17440
rect 34939 17376 34955 17440
rect 35019 17376 35027 17440
rect 34707 16352 35027 17376
rect 34707 16288 34715 16352
rect 34779 16288 34795 16352
rect 34859 16288 34875 16352
rect 34939 16288 34955 16352
rect 35019 16288 35027 16352
rect 34707 15264 35027 16288
rect 34707 15200 34715 15264
rect 34779 15200 34795 15264
rect 34859 15200 34875 15264
rect 34939 15200 34955 15264
rect 35019 15200 35027 15264
rect 34707 14176 35027 15200
rect 34707 14112 34715 14176
rect 34779 14112 34795 14176
rect 34859 14112 34875 14176
rect 34939 14112 34955 14176
rect 35019 14112 35027 14176
rect 34707 13088 35027 14112
rect 34707 13024 34715 13088
rect 34779 13024 34795 13088
rect 34859 13024 34875 13088
rect 34939 13024 34955 13088
rect 35019 13024 35027 13088
rect 34707 12000 35027 13024
rect 34707 11936 34715 12000
rect 34779 11936 34795 12000
rect 34859 11936 34875 12000
rect 34939 11936 34955 12000
rect 35019 11936 35027 12000
rect 34707 10912 35027 11936
rect 34707 10848 34715 10912
rect 34779 10848 34795 10912
rect 34859 10848 34875 10912
rect 34939 10848 34955 10912
rect 35019 10848 35027 10912
rect 34707 9824 35027 10848
rect 34707 9760 34715 9824
rect 34779 9760 34795 9824
rect 34859 9760 34875 9824
rect 34939 9760 34955 9824
rect 35019 9760 35027 9824
rect 34707 8736 35027 9760
rect 34707 8672 34715 8736
rect 34779 8672 34795 8736
rect 34859 8672 34875 8736
rect 34939 8672 34955 8736
rect 35019 8672 35027 8736
rect 34707 7648 35027 8672
rect 34707 7584 34715 7648
rect 34779 7584 34795 7648
rect 34859 7584 34875 7648
rect 34939 7584 34955 7648
rect 35019 7584 35027 7648
rect 34707 6560 35027 7584
rect 34707 6496 34715 6560
rect 34779 6496 34795 6560
rect 34859 6496 34875 6560
rect 34939 6496 34955 6560
rect 35019 6496 35027 6560
rect 34707 5472 35027 6496
rect 34707 5408 34715 5472
rect 34779 5408 34795 5472
rect 34859 5408 34875 5472
rect 34939 5408 34955 5472
rect 35019 5408 35027 5472
rect 34707 4384 35027 5408
rect 34707 4320 34715 4384
rect 34779 4320 34795 4384
rect 34859 4320 34875 4384
rect 34939 4320 34955 4384
rect 35019 4320 35027 4384
rect 34707 3296 35027 4320
rect 34707 3232 34715 3296
rect 34779 3232 34795 3296
rect 34859 3232 34875 3296
rect 34939 3232 34955 3296
rect 35019 3232 35027 3296
rect 34707 2208 35027 3232
rect 34707 2144 34715 2208
rect 34779 2144 34795 2208
rect 34859 2144 34875 2208
rect 34939 2144 34955 2208
rect 35019 2144 35027 2208
rect 34707 2128 35027 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37
timestamp 1666464484
transform 1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43
timestamp 1666464484
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp 1666464484
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1666464484
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1666464484
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp 1666464484
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1666464484
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1666464484
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1666464484
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1666464484
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1666464484
transform 1 0 14812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_155
timestamp 1666464484
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1666464484
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_177
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1666464484
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1666464484
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_205
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_211
timestamp 1666464484
transform 1 0 20516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1666464484
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_233
timestamp 1666464484
transform 1 0 22540 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_239
timestamp 1666464484
transform 1 0 23092 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1666464484
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_261
timestamp 1666464484
transform 1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_267
timestamp 1666464484
transform 1 0 25668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1666464484
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_289
timestamp 1666464484
transform 1 0 27692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_295
timestamp 1666464484
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302
timestamp 1666464484
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_314
timestamp 1666464484
transform 1 0 29992 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_322
timestamp 1666464484
transform 1 0 30728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1666464484
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1666464484
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_342
timestamp 1666464484
transform 1 0 32568 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_350
timestamp 1666464484
transform 1 0 33304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_355
timestamp 1666464484
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1666464484
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1666464484
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_126
timestamp 1666464484
transform 1 0 12696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1666464484
transform 1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_156
timestamp 1666464484
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1666464484
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_203
timestamp 1666464484
transform 1 0 19780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1666464484
transform 1 0 20516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1666464484
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1666464484
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1666464484
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1666464484
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1666464484
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_361
timestamp 1666464484
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1666464484
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_159
timestamp 1666464484
transform 1 0 15732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1666464484
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_185
timestamp 1666464484
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1666464484
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_215
timestamp 1666464484
transform 1 0 20884 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1666464484
transform 1 0 21988 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1666464484
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 1666464484
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1666464484
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1666464484
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_296
timestamp 1666464484
transform 1 0 28336 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1666464484
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1666464484
transform 1 0 8924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1666464484
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1666464484
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_138
timestamp 1666464484
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_174
timestamp 1666464484
transform 1 0 17112 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_196
timestamp 1666464484
transform 1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1666464484
transform 1 0 19872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_243
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_251
timestamp 1666464484
transform 1 0 24196 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_268
timestamp 1666464484
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_299
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_311
timestamp 1666464484
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_323
timestamp 1666464484
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1666464484
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1666464484
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp 1666464484
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_107
timestamp 1666464484
transform 1 0 10948 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1666464484
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_124
timestamp 1666464484
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1666464484
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_147
timestamp 1666464484
transform 1 0 14628 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_155
timestamp 1666464484
transform 1 0 15364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_166
timestamp 1666464484
transform 1 0 16376 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp 1666464484
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1666464484
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1666464484
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_212
timestamp 1666464484
transform 1 0 20608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_220
timestamp 1666464484
transform 1 0 21344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_224
timestamp 1666464484
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_231
timestamp 1666464484
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1666464484
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_261
timestamp 1666464484
transform 1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_285
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_297
timestamp 1666464484
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1666464484
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1666464484
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1666464484
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1666464484
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_36
timestamp 1666464484
transform 1 0 4416 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1666464484
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1666464484
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1666464484
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1666464484
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1666464484
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_139
timestamp 1666464484
transform 1 0 13892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_154
timestamp 1666464484
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1666464484
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_185
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1666464484
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1666464484
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1666464484
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1666464484
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1666464484
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1666464484
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1666464484
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1666464484
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp 1666464484
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_55
timestamp 1666464484
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_67
timestamp 1666464484
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1666464484
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_271
timestamp 1666464484
transform 1 0 26036 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_283
timestamp 1666464484
transform 1 0 27140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_295
timestamp 1666464484
transform 1 0 28244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_299
timestamp 1666464484
transform 1 0 28612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666464484
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1666464484
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1666464484
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1666464484
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1666464484
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 1666464484
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_68
timestamp 1666464484
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_80
timestamp 1666464484
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1666464484
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1666464484
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_134
timestamp 1666464484
transform 1 0 13432 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_146
timestamp 1666464484
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 1666464484
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1666464484
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_260
timestamp 1666464484
transform 1 0 25024 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_272
timestamp 1666464484
transform 1 0 26128 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_313
timestamp 1666464484
transform 1 0 29900 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_325
timestamp 1666464484
transform 1 0 31004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1666464484
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1666464484
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1666464484
transform 1 0 6900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1666464484
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp 1666464484
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1666464484
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_173
timestamp 1666464484
transform 1 0 17020 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1666464484
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1666464484
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_235
timestamp 1666464484
transform 1 0 22724 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_243
timestamp 1666464484
transform 1 0 23460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_271
timestamp 1666464484
transform 1 0 26036 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_283
timestamp 1666464484
transform 1 0 27140 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666464484
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_331
timestamp 1666464484
transform 1 0 31556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_343
timestamp 1666464484
transform 1 0 32660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1666464484
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1666464484
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_18
timestamp 1666464484
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_30
timestamp 1666464484
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1666464484
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1666464484
transform 1 0 8372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1666464484
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1666464484
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1666464484
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1666464484
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1666464484
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_233
timestamp 1666464484
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp 1666464484
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1666464484
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1666464484
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1666464484
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1666464484
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1666464484
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1666464484
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1666464484
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_61
timestamp 1666464484
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_69
timestamp 1666464484
transform 1 0 7452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1666464484
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1666464484
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_99
timestamp 1666464484
transform 1 0 10212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_111
timestamp 1666464484
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 1666464484
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1666464484
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1666464484
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1666464484
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1666464484
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1666464484
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_275
timestamp 1666464484
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_287
timestamp 1666464484
transform 1 0 27508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1666464484
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1666464484
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1666464484
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1666464484
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1666464484
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1666464484
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1666464484
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1666464484
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1666464484
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1666464484
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1666464484
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_233
timestamp 1666464484
transform 1 0 22540 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_241
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1666464484
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1666464484
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_315
timestamp 1666464484
transform 1 0 30084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_325
timestamp 1666464484
transform 1 0 31004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1666464484
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_355
timestamp 1666464484
transform 1 0 33764 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp 1666464484
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1666464484
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_49
timestamp 1666464484
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_61
timestamp 1666464484
transform 1 0 6716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1666464484
transform 1 0 7820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1666464484
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1666464484
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1666464484
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1666464484
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_203
timestamp 1666464484
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_220
timestamp 1666464484
transform 1 0 21344 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1666464484
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1666464484
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_261
timestamp 1666464484
transform 1 0 25116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_273
timestamp 1666464484
transform 1 0 26220 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_285
timestamp 1666464484
transform 1 0 27324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_297
timestamp 1666464484
transform 1 0 28428 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1666464484
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_317
timestamp 1666464484
transform 1 0 30268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_329
timestamp 1666464484
transform 1 0 31372 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_337
timestamp 1666464484
transform 1 0 32108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_355
timestamp 1666464484
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1666464484
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1666464484
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1666464484
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1666464484
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1666464484
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_82
timestamp 1666464484
transform 1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_94
timestamp 1666464484
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1666464484
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_131
timestamp 1666464484
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_143
timestamp 1666464484
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1666464484
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_183
timestamp 1666464484
transform 1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1666464484
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_198
timestamp 1666464484
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_206
timestamp 1666464484
transform 1 0 20056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_216
timestamp 1666464484
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_290
timestamp 1666464484
transform 1 0 27784 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_302
timestamp 1666464484
transform 1 0 28888 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_314
timestamp 1666464484
transform 1 0 29992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_326
timestamp 1666464484
transform 1 0 31096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1666464484
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_359
timestamp 1666464484
transform 1 0 34132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_363
timestamp 1666464484
transform 1 0 34500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1666464484
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1666464484
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1666464484
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_36
timestamp 1666464484
transform 1 0 4416 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1666464484
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_62
timestamp 1666464484
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1666464484
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_126
timestamp 1666464484
transform 1 0 12696 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_220
timestamp 1666464484
transform 1 0 21344 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1666464484
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1666464484
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_271
timestamp 1666464484
transform 1 0 26036 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_283
timestamp 1666464484
transform 1 0 27140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1666464484
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_318
timestamp 1666464484
transform 1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_326
timestamp 1666464484
transform 1 0 31096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_347
timestamp 1666464484
transform 1 0 33028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_19
timestamp 1666464484
transform 1 0 2852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_34
timestamp 1666464484
transform 1 0 4232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_46
timestamp 1666464484
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1666464484
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1666464484
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_100
timestamp 1666464484
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1666464484
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_140
timestamp 1666464484
transform 1 0 13984 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_152
timestamp 1666464484
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1666464484
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_206
timestamp 1666464484
transform 1 0 20056 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1666464484
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 1666464484
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_262
timestamp 1666464484
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1666464484
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1666464484
transform 1 0 28244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1666464484
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_355
timestamp 1666464484
transform 1 0 33764 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_363
timestamp 1666464484
transform 1 0 34500 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_36
timestamp 1666464484
transform 1 0 4416 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_64
timestamp 1666464484
transform 1 0 6992 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1666464484
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_116
timestamp 1666464484
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1666464484
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1666464484
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1666464484
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1666464484
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_212
timestamp 1666464484
transform 1 0 20608 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_222
timestamp 1666464484
transform 1 0 21528 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_234
timestamp 1666464484
transform 1 0 22632 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_242
timestamp 1666464484
transform 1 0 23368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1666464484
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_265
timestamp 1666464484
transform 1 0 25484 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_291
timestamp 1666464484
transform 1 0 27876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1666464484
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_317
timestamp 1666464484
transform 1 0 30268 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_329
timestamp 1666464484
transform 1 0 31372 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1666464484
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1666464484
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_141
timestamp 1666464484
transform 1 0 14076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_151
timestamp 1666464484
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1666464484
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1666464484
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_189
timestamp 1666464484
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1666464484
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1666464484
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_238
timestamp 1666464484
transform 1 0 23000 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_246
timestamp 1666464484
transform 1 0 23736 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1666464484
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_285
timestamp 1666464484
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_302
timestamp 1666464484
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_314
timestamp 1666464484
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1666464484
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_345
timestamp 1666464484
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_357
timestamp 1666464484
transform 1 0 33948 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_363
timestamp 1666464484
transform 1 0 34500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_19
timestamp 1666464484
transform 1 0 2852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1666464484
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1666464484
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1666464484
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_172
timestamp 1666464484
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_205
timestamp 1666464484
transform 1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1666464484
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1666464484
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_261
timestamp 1666464484
transform 1 0 25116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_273
timestamp 1666464484
transform 1 0 26220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_285
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_291
timestamp 1666464484
transform 1 0 27876 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1666464484
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1666464484
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1666464484
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 1666464484
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1666464484
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1666464484
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_94
timestamp 1666464484
transform 1 0 9752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1666464484
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1666464484
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1666464484
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1666464484
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1666464484
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1666464484
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1666464484
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_238
timestamp 1666464484
transform 1 0 23000 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_250
timestamp 1666464484
transform 1 0 24104 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_262
timestamp 1666464484
transform 1 0 25208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1666464484
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_292
timestamp 1666464484
transform 1 0 27968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_302
timestamp 1666464484
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_312
timestamp 1666464484
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_324
timestamp 1666464484
transform 1 0 30912 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_345
timestamp 1666464484
transform 1 0 32844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_357
timestamp 1666464484
transform 1 0 33948 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_363
timestamp 1666464484
transform 1 0 34500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1666464484
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1666464484
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 1666464484
transform 1 0 5152 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_50
timestamp 1666464484
transform 1 0 5704 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_62
timestamp 1666464484
transform 1 0 6808 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_74
timestamp 1666464484
transform 1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_108
timestamp 1666464484
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1666464484
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1666464484
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1666464484
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_171
timestamp 1666464484
transform 1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1666464484
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1666464484
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_205
timestamp 1666464484
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_228
timestamp 1666464484
transform 1 0 22080 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1666464484
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1666464484
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1666464484
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1666464484
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_321
timestamp 1666464484
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1666464484
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1666464484
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_18
timestamp 1666464484
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp 1666464484
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1666464484
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_65
timestamp 1666464484
transform 1 0 7084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_77
timestamp 1666464484
transform 1 0 8188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1666464484
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_96
timestamp 1666464484
transform 1 0 9936 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1666464484
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_146
timestamp 1666464484
transform 1 0 14536 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_154
timestamp 1666464484
transform 1 0 15272 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_180
timestamp 1666464484
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1666464484
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1666464484
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_234
timestamp 1666464484
transform 1 0 22632 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_246
timestamp 1666464484
transform 1 0 23736 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_254
timestamp 1666464484
transform 1 0 24472 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1666464484
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1666464484
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_299
timestamp 1666464484
transform 1 0 28612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1666464484
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_316
timestamp 1666464484
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1666464484
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_358
timestamp 1666464484
transform 1 0 34040 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1666464484
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1666464484
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1666464484
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_96
timestamp 1666464484
transform 1 0 9936 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1666464484
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_120
timestamp 1666464484
transform 1 0 12144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1666464484
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_190
timestamp 1666464484
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_205
timestamp 1666464484
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1666464484
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1666464484
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1666464484
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1666464484
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1666464484
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_330
timestamp 1666464484
transform 1 0 31464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1666464484
transform 1 0 33580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1666464484
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_34
timestamp 1666464484
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1666464484
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1666464484
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1666464484
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1666464484
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_178
timestamp 1666464484
transform 1 0 17480 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_206
timestamp 1666464484
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_216
timestamp 1666464484
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_233
timestamp 1666464484
transform 1 0 22540 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1666464484
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_265
timestamp 1666464484
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1666464484
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1666464484
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1666464484
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_309
timestamp 1666464484
transform 1 0 29532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1666464484
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1666464484
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1666464484
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_359
timestamp 1666464484
transform 1 0 34132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_363
timestamp 1666464484
transform 1 0 34500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1666464484
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_48
timestamp 1666464484
transform 1 0 5520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_64
timestamp 1666464484
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1666464484
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1666464484
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_132
timestamp 1666464484
transform 1 0 13248 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1666464484
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_155
timestamp 1666464484
transform 1 0 15364 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_159
timestamp 1666464484
transform 1 0 15732 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_169
timestamp 1666464484
transform 1 0 16652 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_187
timestamp 1666464484
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1666464484
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1666464484
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1666464484
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_281
timestamp 1666464484
transform 1 0 26956 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_289
timestamp 1666464484
transform 1 0 27692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1666464484
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_321
timestamp 1666464484
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_347
timestamp 1666464484
transform 1 0 33028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_45
timestamp 1666464484
transform 1 0 5244 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1666464484
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_62
timestamp 1666464484
transform 1 0 6808 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_75
timestamp 1666464484
transform 1 0 8004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_86
timestamp 1666464484
transform 1 0 9016 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_94
timestamp 1666464484
transform 1 0 9752 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1666464484
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_136
timestamp 1666464484
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1666464484
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_182
timestamp 1666464484
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1666464484
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1666464484
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_235
timestamp 1666464484
transform 1 0 22724 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_241
timestamp 1666464484
transform 1 0 23276 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_262
timestamp 1666464484
transform 1 0 25208 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_270
timestamp 1666464484
transform 1 0 25944 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1666464484
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_293
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_303
timestamp 1666464484
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_310
timestamp 1666464484
transform 1 0 29624 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_322
timestamp 1666464484
transform 1 0 30728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1666464484
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_356
timestamp 1666464484
transform 1 0 33856 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1666464484
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_36
timestamp 1666464484
transform 1 0 4416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_54
timestamp 1666464484
transform 1 0 6072 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1666464484
transform 1 0 6624 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1666464484
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1666464484
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_100
timestamp 1666464484
transform 1 0 10304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_112
timestamp 1666464484
transform 1 0 11408 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1666464484
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1666464484
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_150
timestamp 1666464484
transform 1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1666464484
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_183
timestamp 1666464484
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1666464484
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_223
timestamp 1666464484
transform 1 0 21620 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_235
timestamp 1666464484
transform 1 0 22724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1666464484
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1666464484
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_281
timestamp 1666464484
transform 1 0 26956 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1666464484
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_319
timestamp 1666464484
transform 1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1666464484
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1666464484
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_343
timestamp 1666464484
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1666464484
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666464484
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_37
timestamp 1666464484
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1666464484
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1666464484
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_78
timestamp 1666464484
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_98
timestamp 1666464484
transform 1 0 10120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_136
timestamp 1666464484
transform 1 0 13616 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_148
timestamp 1666464484
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1666464484
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1666464484
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_182
timestamp 1666464484
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_206
timestamp 1666464484
transform 1 0 20056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1666464484
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_237
timestamp 1666464484
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_256
timestamp 1666464484
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_268
timestamp 1666464484
transform 1 0 25760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1666464484
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_302
timestamp 1666464484
transform 1 0 28888 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_310
timestamp 1666464484
transform 1 0 29624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_314
timestamp 1666464484
transform 1 0 29992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_318
timestamp 1666464484
transform 1 0 30360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_326
timestamp 1666464484
transform 1 0 31096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1666464484
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_344
timestamp 1666464484
transform 1 0 32752 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_351
timestamp 1666464484
transform 1 0 33396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_363
timestamp 1666464484
transform 1 0 34500 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1666464484
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_60
timestamp 1666464484
transform 1 0 6624 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_72
timestamp 1666464484
transform 1 0 7728 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1666464484
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1666464484
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1666464484
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_187
timestamp 1666464484
transform 1 0 18308 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1666464484
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_225
timestamp 1666464484
transform 1 0 21804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_237
timestamp 1666464484
transform 1 0 22908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_261
timestamp 1666464484
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_273
timestamp 1666464484
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_285
timestamp 1666464484
transform 1 0 27324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1666464484
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_321
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_327
timestamp 1666464484
transform 1 0 31188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_336
timestamp 1666464484
transform 1 0 32016 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_345
timestamp 1666464484
transform 1 0 32844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1666464484
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1666464484
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_78
timestamp 1666464484
transform 1 0 8280 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_90
timestamp 1666464484
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_101
timestamp 1666464484
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1666464484
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1666464484
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1666464484
transform 1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1666464484
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_237
timestamp 1666464484
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1666464484
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1666464484
transform 1 0 28152 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_315
timestamp 1666464484
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1666464484
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666464484
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_346
timestamp 1666464484
transform 1 0 32936 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_358
timestamp 1666464484
transform 1 0 34040 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_362
timestamp 1666464484
transform 1 0 34408 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_21
timestamp 1666464484
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1666464484
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1666464484
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_104
timestamp 1666464484
transform 1 0 10672 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1666464484
transform 1 0 11776 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_123
timestamp 1666464484
transform 1 0 12420 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1666464484
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_150
timestamp 1666464484
transform 1 0 14904 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_170
timestamp 1666464484
transform 1 0 16744 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_182
timestamp 1666464484
transform 1 0 17848 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_215
timestamp 1666464484
transform 1 0 20884 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_227
timestamp 1666464484
transform 1 0 21988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_239
timestamp 1666464484
transform 1 0 23092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_243
timestamp 1666464484
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_261
timestamp 1666464484
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_276
timestamp 1666464484
transform 1 0 26496 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_284
timestamp 1666464484
transform 1 0 27232 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1666464484
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1666464484
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_316
timestamp 1666464484
transform 1 0 30176 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_328
timestamp 1666464484
transform 1 0 31280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1666464484
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_349
timestamp 1666464484
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1666464484
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_32
timestamp 1666464484
transform 1 0 4048 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1666464484
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1666464484
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1666464484
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1666464484
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1666464484
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1666464484
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_127
timestamp 1666464484
transform 1 0 12788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_139
timestamp 1666464484
transform 1 0 13892 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_147
timestamp 1666464484
transform 1 0 14628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_177
timestamp 1666464484
transform 1 0 17388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1666464484
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_210
timestamp 1666464484
transform 1 0 20424 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1666464484
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_237
timestamp 1666464484
transform 1 0 22908 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_258
timestamp 1666464484
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1666464484
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_287
timestamp 1666464484
transform 1 0 27508 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_295
timestamp 1666464484
transform 1 0 28244 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_310
timestamp 1666464484
transform 1 0 29624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_322
timestamp 1666464484
transform 1 0 30728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_331
timestamp 1666464484
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_346
timestamp 1666464484
transform 1 0 32936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_358
timestamp 1666464484
transform 1 0 34040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1666464484
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1666464484
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_39
timestamp 1666464484
transform 1 0 4692 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_47
timestamp 1666464484
transform 1 0 5428 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1666464484
transform 1 0 6532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1666464484
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1666464484
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_91
timestamp 1666464484
transform 1 0 9476 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1666464484
transform 1 0 10212 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_118
timestamp 1666464484
transform 1 0 11960 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_130
timestamp 1666464484
transform 1 0 13064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1666464484
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1666464484
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1666464484
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_185
timestamp 1666464484
transform 1 0 18124 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_207
timestamp 1666464484
transform 1 0 20148 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1666464484
transform 1 0 20700 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_234
timestamp 1666464484
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1666464484
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1666464484
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1666464484
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666464484
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1666464484
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_333
timestamp 1666464484
transform 1 0 31740 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1666464484
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1666464484
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_19
timestamp 1666464484
transform 1 0 2852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1666464484
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_74
timestamp 1666464484
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_82
timestamp 1666464484
transform 1 0 8648 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1666464484
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1666464484
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1666464484
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_154
timestamp 1666464484
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1666464484
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_201
timestamp 1666464484
transform 1 0 19596 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1666464484
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1666464484
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_237
timestamp 1666464484
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_260
timestamp 1666464484
transform 1 0 25024 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1666464484
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1666464484
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1666464484
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1666464484
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1666464484
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_348
timestamp 1666464484
transform 1 0 33120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_360
timestamp 1666464484
transform 1 0 34224 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1666464484
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_72
timestamp 1666464484
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_105
timestamp 1666464484
transform 1 0 10764 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_117
timestamp 1666464484
transform 1 0 11868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1666464484
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1666464484
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_149
timestamp 1666464484
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1666464484
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1666464484
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1666464484
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_208
timestamp 1666464484
transform 1 0 20240 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_234
timestamp 1666464484
transform 1 0 22632 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_242
timestamp 1666464484
transform 1 0 23368 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_261
timestamp 1666464484
transform 1 0 25116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_273
timestamp 1666464484
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_285
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1666464484
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_321
timestamp 1666464484
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_327
timestamp 1666464484
transform 1 0 31188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1666464484
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_342
timestamp 1666464484
transform 1 0 32568 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_349
timestamp 1666464484
transform 1 0 33212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1666464484
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1666464484
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_34
timestamp 1666464484
transform 1 0 4232 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_46
timestamp 1666464484
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1666464484
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_120
timestamp 1666464484
transform 1 0 12144 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_132
timestamp 1666464484
transform 1 0 13248 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_144
timestamp 1666464484
transform 1 0 14352 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_148
timestamp 1666464484
transform 1 0 14720 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1666464484
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1666464484
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1666464484
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_232
timestamp 1666464484
transform 1 0 22448 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_259
timestamp 1666464484
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_271
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1666464484
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_309
timestamp 1666464484
transform 1 0 29532 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_315
timestamp 1666464484
transform 1 0 30084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_320
timestamp 1666464484
transform 1 0 30544 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_328
timestamp 1666464484
transform 1 0 31280 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1666464484
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1666464484
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_61
timestamp 1666464484
transform 1 0 6716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_68
timestamp 1666464484
transform 1 0 7360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_76
timestamp 1666464484
transform 1 0 8096 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1666464484
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1666464484
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1666464484
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_188
timestamp 1666464484
transform 1 0 18400 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1666464484
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1666464484
transform 1 0 20240 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1666464484
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1666464484
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_263
timestamp 1666464484
transform 1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_274
timestamp 1666464484
transform 1 0 26312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_291
timestamp 1666464484
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_300
timestamp 1666464484
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_318
timestamp 1666464484
transform 1 0 30360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1666464484
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_332
timestamp 1666464484
transform 1 0 31648 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1666464484
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_347
timestamp 1666464484
transform 1 0 33028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1666464484
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1666464484
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_35
timestamp 1666464484
transform 1 0 4324 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_43
timestamp 1666464484
transform 1 0 5060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_65
timestamp 1666464484
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_72
timestamp 1666464484
transform 1 0 7728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1666464484
transform 1 0 9752 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1666464484
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1666464484
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_122
timestamp 1666464484
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_140
timestamp 1666464484
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_148
timestamp 1666464484
transform 1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_158
timestamp 1666464484
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1666464484
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_175
timestamp 1666464484
transform 1 0 17204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1666464484
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_191
timestamp 1666464484
transform 1 0 18676 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_210
timestamp 1666464484
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_230
timestamp 1666464484
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_242
timestamp 1666464484
transform 1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_248
timestamp 1666464484
transform 1 0 23920 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_254
timestamp 1666464484
transform 1 0 24472 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1666464484
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1666464484
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_307
timestamp 1666464484
transform 1 0 29348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_316
timestamp 1666464484
transform 1 0 30176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_322
timestamp 1666464484
transform 1 0 30728 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1666464484
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1666464484
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_359
timestamp 1666464484
transform 1 0 34132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_363
timestamp 1666464484
transform 1 0 34500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_21
timestamp 1666464484
transform 1 0 3036 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1666464484
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_36
timestamp 1666464484
transform 1 0 4416 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_48
timestamp 1666464484
transform 1 0 5520 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_60
timestamp 1666464484
transform 1 0 6624 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_71
timestamp 1666464484
transform 1 0 7636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1666464484
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_91
timestamp 1666464484
transform 1 0 9476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_120
timestamp 1666464484
transform 1 0 12144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1666464484
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1666464484
transform 1 0 14812 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1666464484
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_168
timestamp 1666464484
transform 1 0 16560 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1666464484
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_204
timestamp 1666464484
transform 1 0 19872 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_232
timestamp 1666464484
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1666464484
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_264
timestamp 1666464484
transform 1 0 25392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_276
timestamp 1666464484
transform 1 0 26496 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_284
timestamp 1666464484
transform 1 0 27232 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_296
timestamp 1666464484
transform 1 0 28336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_321
timestamp 1666464484
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_338
timestamp 1666464484
transform 1 0 32200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_349
timestamp 1666464484
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1666464484
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1666464484
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1666464484
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1666464484
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_100
timestamp 1666464484
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_135
timestamp 1666464484
transform 1 0 13524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_141
timestamp 1666464484
transform 1 0 14076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1666464484
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_157
timestamp 1666464484
transform 1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1666464484
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_185
timestamp 1666464484
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1666464484
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1666464484
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_236
timestamp 1666464484
transform 1 0 22816 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_248
timestamp 1666464484
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_260
timestamp 1666464484
transform 1 0 25024 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_266
timestamp 1666464484
transform 1 0 25576 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1666464484
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1666464484
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_319
timestamp 1666464484
transform 1 0 30452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1666464484
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666464484
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1666464484
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_14
timestamp 1666464484
transform 1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1666464484
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1666464484
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_51
timestamp 1666464484
transform 1 0 5796 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_59
timestamp 1666464484
transform 1 0 6532 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1666464484
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_120
timestamp 1666464484
transform 1 0 12144 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1666464484
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_150
timestamp 1666464484
transform 1 0 14904 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_161
timestamp 1666464484
transform 1 0 15916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_176
timestamp 1666464484
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_186
timestamp 1666464484
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_217
timestamp 1666464484
transform 1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1666464484
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1666464484
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_261
timestamp 1666464484
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1666464484
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_317
timestamp 1666464484
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_326
timestamp 1666464484
transform 1 0 31096 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_338
timestamp 1666464484
transform 1 0 32200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_350
timestamp 1666464484
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1666464484
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1666464484
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_32
timestamp 1666464484
transform 1 0 4048 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1666464484
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1666464484
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_75
timestamp 1666464484
transform 1 0 8004 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_87
timestamp 1666464484
transform 1 0 9108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1666464484
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_157
timestamp 1666464484
transform 1 0 15548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1666464484
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_201
timestamp 1666464484
transform 1 0 19596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_213
timestamp 1666464484
transform 1 0 20700 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_246
timestamp 1666464484
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_258
timestamp 1666464484
transform 1 0 24840 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_265
timestamp 1666464484
transform 1 0 25484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1666464484
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1666464484
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_313
timestamp 1666464484
transform 1 0 29900 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_331
timestamp 1666464484
transform 1 0 31556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1666464484
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_36
timestamp 1666464484
transform 1 0 4416 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_48
timestamp 1666464484
transform 1 0 5520 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_60
timestamp 1666464484
transform 1 0 6624 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_64
timestamp 1666464484
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1666464484
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_127
timestamp 1666464484
transform 1 0 12788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_158
timestamp 1666464484
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1666464484
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_178
timestamp 1666464484
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1666464484
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1666464484
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1666464484
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_261
timestamp 1666464484
transform 1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_269
timestamp 1666464484
transform 1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_278
timestamp 1666464484
transform 1 0 26680 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_287
timestamp 1666464484
transform 1 0 27508 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_293
timestamp 1666464484
transform 1 0 28060 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1666464484
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1666464484
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_332
timestamp 1666464484
transform 1 0 31648 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_344
timestamp 1666464484
transform 1 0 32752 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1666464484
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_89
timestamp 1666464484
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1666464484
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_126
timestamp 1666464484
transform 1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_136
timestamp 1666464484
transform 1 0 13616 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_148
timestamp 1666464484
transform 1 0 14720 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1666464484
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_177
timestamp 1666464484
transform 1 0 17388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_202
timestamp 1666464484
transform 1 0 19688 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_210
timestamp 1666464484
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1666464484
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_246
timestamp 1666464484
transform 1 0 23736 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_257
timestamp 1666464484
transform 1 0 24748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1666464484
transform 1 0 25668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1666464484
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_290
timestamp 1666464484
transform 1 0 27784 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1666464484
transform 1 0 28520 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_319
timestamp 1666464484
transform 1 0 30452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1666464484
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_345
timestamp 1666464484
transform 1 0 32844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_357
timestamp 1666464484
transform 1 0 33948 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_363
timestamp 1666464484
transform 1 0 34500 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_93
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_105
timestamp 1666464484
transform 1 0 10764 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1666464484
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_120
timestamp 1666464484
transform 1 0 12144 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_128
timestamp 1666464484
transform 1 0 12880 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1666464484
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1666464484
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1666464484
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_205
timestamp 1666464484
transform 1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1666464484
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_234
timestamp 1666464484
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1666464484
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_270
timestamp 1666464484
transform 1 0 25944 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_283
timestamp 1666464484
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_293
timestamp 1666464484
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1666464484
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_313
timestamp 1666464484
transform 1 0 29900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_334
timestamp 1666464484
transform 1 0 31832 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_344
timestamp 1666464484
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1666464484
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_92
timestamp 1666464484
transform 1 0 9568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1666464484
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_121
timestamp 1666464484
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_133
timestamp 1666464484
transform 1 0 13340 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_140
timestamp 1666464484
transform 1 0 13984 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1666464484
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_185
timestamp 1666464484
transform 1 0 18124 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_206
timestamp 1666464484
transform 1 0 20056 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1666464484
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_236
timestamp 1666464484
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_248
timestamp 1666464484
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_256
timestamp 1666464484
transform 1 0 24656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1666464484
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_288
timestamp 1666464484
transform 1 0 27600 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_300
timestamp 1666464484
transform 1 0 28704 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_308
timestamp 1666464484
transform 1 0 29440 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1666464484
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_99
timestamp 1666464484
transform 1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_111
timestamp 1666464484
transform 1 0 11316 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_123
timestamp 1666464484
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1666464484
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_152
timestamp 1666464484
transform 1 0 15088 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_160
timestamp 1666464484
transform 1 0 15824 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1666464484
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1666464484
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_282
timestamp 1666464484
transform 1 0 27048 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_292
timestamp 1666464484
transform 1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1666464484
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_328
timestamp 1666464484
transform 1 0 31280 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_340
timestamp 1666464484
transform 1 0 32384 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_352
timestamp 1666464484
transform 1 0 33488 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_78
timestamp 1666464484
transform 1 0 8280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_89
timestamp 1666464484
transform 1 0 9292 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_96
timestamp 1666464484
transform 1 0 9936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1666464484
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_134
timestamp 1666464484
transform 1 0 13432 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_143
timestamp 1666464484
transform 1 0 14260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1666464484
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_162
timestamp 1666464484
transform 1 0 16008 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_200
timestamp 1666464484
transform 1 0 19504 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1666464484
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1666464484
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1666464484
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1666464484
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_246
timestamp 1666464484
transform 1 0 23736 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1666464484
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_288
timestamp 1666464484
transform 1 0 27600 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_300
timestamp 1666464484
transform 1 0 28704 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_312
timestamp 1666464484
transform 1 0 29808 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_319
timestamp 1666464484
transform 1 0 30452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1666464484
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_93
timestamp 1666464484
transform 1 0 9660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_105
timestamp 1666464484
transform 1 0 10764 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_124
timestamp 1666464484
transform 1 0 12512 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1666464484
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_157
timestamp 1666464484
transform 1 0 15548 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_170
timestamp 1666464484
transform 1 0 16744 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_182
timestamp 1666464484
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1666464484
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1666464484
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_219
timestamp 1666464484
transform 1 0 21252 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_227
timestamp 1666464484
transform 1 0 21988 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1666464484
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_271
timestamp 1666464484
transform 1 0 26036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_293
timestamp 1666464484
transform 1 0 28060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_299
timestamp 1666464484
transform 1 0 28612 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_303
timestamp 1666464484
transform 1 0 28980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_92
timestamp 1666464484
transform 1 0 9568 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_104
timestamp 1666464484
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_136
timestamp 1666464484
transform 1 0 13616 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_144
timestamp 1666464484
transform 1 0 14352 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_151
timestamp 1666464484
transform 1 0 14996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_160
timestamp 1666464484
transform 1 0 15824 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_177
timestamp 1666464484
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1666464484
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_214
timestamp 1666464484
transform 1 0 20792 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1666464484
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_236
timestamp 1666464484
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_248
timestamp 1666464484
transform 1 0 23920 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_260
timestamp 1666464484
transform 1 0 25024 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_267
timestamp 1666464484
transform 1 0 25668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1666464484
transform 1 0 27416 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_296
timestamp 1666464484
transform 1 0 28336 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_105
timestamp 1666464484
transform 1 0 10764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_117
timestamp 1666464484
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_125
timestamp 1666464484
transform 1 0 12604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_132
timestamp 1666464484
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1666464484
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_212
timestamp 1666464484
transform 1 0 20608 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_223
timestamp 1666464484
transform 1 0 21620 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_235
timestamp 1666464484
transform 1 0 22724 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1666464484
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_262
timestamp 1666464484
transform 1 0 25208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_274
timestamp 1666464484
transform 1 0 26312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_282
timestamp 1666464484
transform 1 0 27048 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_292
timestamp 1666464484
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1666464484
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_316
timestamp 1666464484
transform 1 0 30176 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_328
timestamp 1666464484
transform 1 0 31280 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_340
timestamp 1666464484
transform 1 0 32384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_352
timestamp 1666464484
transform 1 0 33488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_133
timestamp 1666464484
transform 1 0 13340 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_156
timestamp 1666464484
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_187
timestamp 1666464484
transform 1 0 18308 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_210
timestamp 1666464484
transform 1 0 20424 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_255
timestamp 1666464484
transform 1 0 24564 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_294
timestamp 1666464484
transform 1 0 28152 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_306
timestamp 1666464484
transform 1 0 29256 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_315
timestamp 1666464484
transform 1 0 30084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1666464484
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_92
timestamp 1666464484
transform 1 0 9568 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1666464484
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_106
timestamp 1666464484
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_118
timestamp 1666464484
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_130
timestamp 1666464484
transform 1 0 13064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1666464484
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1666464484
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_167
timestamp 1666464484
transform 1 0 16468 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_174
timestamp 1666464484
transform 1 0 17112 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_186
timestamp 1666464484
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1666464484
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_217
timestamp 1666464484
transform 1 0 21068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_229
timestamp 1666464484
transform 1 0 22172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_241
timestamp 1666464484
transform 1 0 23276 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1666464484
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_276
timestamp 1666464484
transform 1 0 26496 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_284
timestamp 1666464484
transform 1 0 27232 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1666464484
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666464484
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1666464484
transform 1 0 9568 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1666464484
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1666464484
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_156
timestamp 1666464484
transform 1 0 15456 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_162
timestamp 1666464484
transform 1 0 16008 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1666464484
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1666464484
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_182
timestamp 1666464484
transform 1 0 17848 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_194
timestamp 1666464484
transform 1 0 18952 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1666464484
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_246
timestamp 1666464484
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_250
timestamp 1666464484
transform 1 0 24104 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1666464484
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1666464484
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666464484
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_292
timestamp 1666464484
transform 1 0 27968 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1666464484
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_98
timestamp 1666464484
transform 1 0 10120 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_106
timestamp 1666464484
transform 1 0 10856 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_117
timestamp 1666464484
transform 1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1666464484
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_146
timestamp 1666464484
transform 1 0 14536 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_154
timestamp 1666464484
transform 1 0 15272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_162
timestamp 1666464484
transform 1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_180
timestamp 1666464484
transform 1 0 17664 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1666464484
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1666464484
transform 1 0 20608 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_220
timestamp 1666464484
transform 1 0 21344 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_226
timestamp 1666464484
transform 1 0 21896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_239
timestamp 1666464484
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1666464484
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_264
timestamp 1666464484
transform 1 0 25392 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_292
timestamp 1666464484
transform 1 0 27968 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1666464484
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_89
timestamp 1666464484
transform 1 0 9292 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_97
timestamp 1666464484
transform 1 0 10028 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_124
timestamp 1666464484
transform 1 0 12512 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1666464484
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_187
timestamp 1666464484
transform 1 0 18308 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_199
timestamp 1666464484
transform 1 0 19412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_211
timestamp 1666464484
transform 1 0 20516 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1666464484
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_230
timestamp 1666464484
transform 1 0 22264 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_241
timestamp 1666464484
transform 1 0 23276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_253
timestamp 1666464484
transform 1 0 24380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_257
timestamp 1666464484
transform 1 0 24748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1666464484
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1666464484
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_313
timestamp 1666464484
transform 1 0 29900 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_320
timestamp 1666464484
transform 1 0 30544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1666464484
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_345
timestamp 1666464484
transform 1 0 32844 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_351
timestamp 1666464484
transform 1 0 33396 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_363
timestamp 1666464484
transform 1 0 34500 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_100
timestamp 1666464484
transform 1 0 10304 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_112
timestamp 1666464484
transform 1 0 11408 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_124
timestamp 1666464484
transform 1 0 12512 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1666464484
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_159
timestamp 1666464484
transform 1 0 15732 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_172
timestamp 1666464484
transform 1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_184
timestamp 1666464484
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_216
timestamp 1666464484
transform 1 0 20976 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_228
timestamp 1666464484
transform 1 0 22080 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666464484
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_29
timestamp 1666464484
transform 1 0 3772 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_37
timestamp 1666464484
transform 1 0 4508 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1666464484
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_76
timestamp 1666464484
transform 1 0 8096 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_85
timestamp 1666464484
transform 1 0 8924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_97
timestamp 1666464484
transform 1 0 10028 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_103
timestamp 1666464484
transform 1 0 10580 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1666464484
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1666464484
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_147
timestamp 1666464484
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1666464484
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_175
timestamp 1666464484
transform 1 0 17204 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_187
timestamp 1666464484
transform 1 0 18308 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_195
timestamp 1666464484
transform 1 0 19044 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_197
timestamp 1666464484
transform 1 0 19228 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_204
timestamp 1666464484
transform 1 0 19872 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_216
timestamp 1666464484
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_231
timestamp 1666464484
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_236
timestamp 1666464484
transform 1 0 22816 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_248
timestamp 1666464484
transform 1 0 23920 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_253
timestamp 1666464484
transform 1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_261
timestamp 1666464484
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_268
timestamp 1666464484
transform 1 0 25760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_300
timestamp 1666464484
transform 1 0 28704 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_309
timestamp 1666464484
transform 1 0 29532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_321
timestamp 1666464484
transform 1 0 30636 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_327
timestamp 1666464484
transform 1 0 31188 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1666464484
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_349
timestamp 1666464484
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_357
timestamp 1666464484
transform 1 0 33948 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_362
timestamp 1666464484
transform 1 0 34408 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 34868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 34868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 34868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 34868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 34868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 34868 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 34868 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 34868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 34868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 34868 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 34868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 34868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 34868 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 34868 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 34868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 34868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 34868 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 34868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 34868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 34868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 34868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 34868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 34868 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 34868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 34868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 34868 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 34868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 34868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 34868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 34868 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 34868 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1666464484
transform -1 0 4232 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4416 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1666464484
transform 1 0 14444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1666464484
transform 1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0471_
timestamp 1666464484
transform 1 0 12604 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1666464484
transform 1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _0473_
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _0474_
timestamp 1666464484
transform 1 0 9568 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0475_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13616 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1666464484
transform -1 0 25576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1666464484
transform -1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1666464484
transform 1 0 28704 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0480_
timestamp 1666464484
transform -1 0 33396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0481_
timestamp 1666464484
transform -1 0 30544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0482__1
timestamp 1666464484
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1666464484
transform -1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1666464484
transform 1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1666464484
transform -1 0 2300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26128 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0488_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5336 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9568 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10304 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__mux2_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0493_
timestamp 1666464484
transform -1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0494_
timestamp 1666464484
transform 1 0 22080 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0495_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11868 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20700 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0499_
timestamp 1666464484
transform -1 0 12604 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10672 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_4  _0501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _0502_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15824 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0503_
timestamp 1666464484
transform 1 0 14168 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0504_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15364 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1666464484
transform -1 0 13616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0506_
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0507_
timestamp 1666464484
transform 1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0508_
timestamp 1666464484
transform 1 0 7360 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0509_
timestamp 1666464484
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0510_
timestamp 1666464484
transform -1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0511_
timestamp 1666464484
transform 1 0 19780 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0512_
timestamp 1666464484
transform 1 0 7268 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0513_
timestamp 1666464484
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1666464484
transform 1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6624 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0516_
timestamp 1666464484
transform -1 0 7360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0517_
timestamp 1666464484
transform 1 0 18032 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0518_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8648 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1666464484
transform 1 0 16928 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0520_
timestamp 1666464484
transform 1 0 12144 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0521_
timestamp 1666464484
transform 1 0 15548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0522_
timestamp 1666464484
transform 1 0 12328 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1666464484
transform -1 0 14812 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _0524_
timestamp 1666464484
transform 1 0 6624 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0525_
timestamp 1666464484
transform 1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0526_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3036 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0527_
timestamp 1666464484
transform 1 0 26404 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_2  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11040 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0529_
timestamp 1666464484
transform 1 0 11684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0530_
timestamp 1666464484
transform 1 0 12880 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16928 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0532_
timestamp 1666464484
transform 1 0 2576 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1666464484
transform 1 0 8740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0535_
timestamp 1666464484
transform -1 0 4232 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0536_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2944 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0537_
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0538_
timestamp 1666464484
transform -1 0 3128 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0539_
timestamp 1666464484
transform 1 0 2852 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_2  _0540_
timestamp 1666464484
transform -1 0 3404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0541_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1666464484
transform -1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0543_
timestamp 1666464484
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0546_
timestamp 1666464484
transform -1 0 15916 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0547_
timestamp 1666464484
transform -1 0 13248 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0548_
timestamp 1666464484
transform -1 0 14260 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0549_
timestamp 1666464484
transform -1 0 25484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27508 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0551_
timestamp 1666464484
transform 1 0 25944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0552_
timestamp 1666464484
transform 1 0 27140 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0553_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27140 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0554_
timestamp 1666464484
transform -1 0 28612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0555_
timestamp 1666464484
transform -1 0 27600 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0556_
timestamp 1666464484
transform -1 0 24748 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0557_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26680 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0559_
timestamp 1666464484
transform 1 0 27140 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_2  _0560_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25116 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _0561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26312 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__a32o_4  _0562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26496 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28704 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0564_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0565_
timestamp 1666464484
transform 1 0 29716 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _0566_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27048 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_2  _0567_
timestamp 1666464484
transform 1 0 24656 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1666464484
transform 1 0 24472 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0569_
timestamp 1666464484
transform -1 0 25668 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0570_
timestamp 1666464484
transform -1 0 27968 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_8  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26128 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27968 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0573_
timestamp 1666464484
transform -1 0 27416 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0574_
timestamp 1666464484
transform 1 0 29624 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0575_
timestamp 1666464484
transform -1 0 28336 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28520 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_2  _0577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_4  _0578_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24932 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o31a_2  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27232 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28980 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__o311a_4  _0581_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24656 0 -1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _0582_
timestamp 1666464484
transform -1 0 22816 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0583_
timestamp 1666464484
transform -1 0 23276 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0584_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27324 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _0585_
timestamp 1666464484
transform -1 0 26036 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0586_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25944 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29164 0 -1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1666464484
transform -1 0 22540 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0589_
timestamp 1666464484
transform -1 0 19504 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0590_
timestamp 1666464484
transform 1 0 20240 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1666464484
transform -1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0592_
timestamp 1666464484
transform 1 0 19780 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0593_
timestamp 1666464484
transform -1 0 23736 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_4  _0594_
timestamp 1666464484
transform -1 0 24104 0 1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_2  _0595_
timestamp 1666464484
transform -1 0 21620 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _0596_
timestamp 1666464484
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1666464484
transform 1 0 20608 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0598_
timestamp 1666464484
transform -1 0 21252 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1666464484
transform -1 0 21344 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23920 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0601_
timestamp 1666464484
transform 1 0 22724 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_4  _0602_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 22172 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__or3b_1  _0603_
timestamp 1666464484
transform 1 0 24196 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0604_
timestamp 1666464484
transform 1 0 24564 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0606_
timestamp 1666464484
transform -1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_4  _0607_
timestamp 1666464484
transform 1 0 20056 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 20608 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1666464484
transform -1 0 17848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0610_
timestamp 1666464484
transform -1 0 15824 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0611_
timestamp 1666464484
transform -1 0 14996 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0612_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15180 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0614_
timestamp 1666464484
transform -1 0 19688 0 -1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_1  _0615_
timestamp 1666464484
transform -1 0 13800 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _0616_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20056 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _0617_
timestamp 1666464484
transform -1 0 20424 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0618_
timestamp 1666464484
transform -1 0 16376 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16468 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _0620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 1666464484
transform -1 0 22264 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0622_
timestamp 1666464484
transform 1 0 20700 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _0623_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17664 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__a21boi_2  _0625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16008 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0626_
timestamp 1666464484
transform -1 0 15548 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _0627_
timestamp 1666464484
transform -1 0 13432 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0628_
timestamp 1666464484
transform 1 0 12972 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1666464484
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0630_
timestamp 1666464484
transform -1 0 13800 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1666464484
transform -1 0 10304 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 1666464484
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13984 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_4  _0634_
timestamp 1666464484
transform -1 0 15456 0 -1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0635_
timestamp 1666464484
transform -1 0 10212 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _0636_
timestamp 1666464484
transform 1 0 11684 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _0637_
timestamp 1666464484
transform -1 0 9568 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0638_
timestamp 1666464484
transform 1 0 15548 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0639_
timestamp 1666464484
transform 1 0 16836 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1666464484
transform -1 0 17112 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0641_
timestamp 1666464484
transform -1 0 18308 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0642_
timestamp 1666464484
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0643_
timestamp 1666464484
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_4  _0644_
timestamp 1666464484
transform 1 0 9936 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__o211ai_4  _0645_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12512 0 1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _0646_
timestamp 1666464484
transform 1 0 9476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10764 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9568 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0649_
timestamp 1666464484
transform 1 0 9108 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0650_
timestamp 1666464484
transform -1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0651_
timestamp 1666464484
transform 1 0 7728 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0652_
timestamp 1666464484
transform 1 0 12880 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11868 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _0654_
timestamp 1666464484
transform -1 0 13708 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0655_
timestamp 1666464484
transform -1 0 17296 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0656_
timestamp 1666464484
transform -1 0 15916 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1666464484
transform -1 0 14444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0658_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16376 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0659_
timestamp 1666464484
transform -1 0 15640 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0660_
timestamp 1666464484
transform -1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1666464484
transform -1 0 16192 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0662_
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0663_
timestamp 1666464484
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0664_
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1666464484
transform -1 0 8648 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0666_
timestamp 1666464484
transform 1 0 8924 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 1666464484
transform 1 0 9292 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0668_
timestamp 1666464484
transform -1 0 9292 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0669_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1666464484
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0671_
timestamp 1666464484
transform -1 0 8556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0672_
timestamp 1666464484
transform -1 0 9568 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0673_
timestamp 1666464484
transform 1 0 16192 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0674_
timestamp 1666464484
transform -1 0 16376 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0675_
timestamp 1666464484
transform -1 0 10764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1666464484
transform -1 0 10028 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15364 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0678_
timestamp 1666464484
transform -1 0 16652 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0679_
timestamp 1666464484
transform -1 0 16376 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_4  _0680_
timestamp 1666464484
transform 1 0 17664 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0681_
timestamp 1666464484
transform -1 0 32568 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0682_
timestamp 1666464484
transform 1 0 31832 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1666464484
transform -1 0 32660 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0684_
timestamp 1666464484
transform 1 0 32292 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1666464484
transform -1 0 29624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31096 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0688_
timestamp 1666464484
transform 1 0 32292 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _0689_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31924 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0690_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1666464484
transform -1 0 33212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0692_
timestamp 1666464484
transform -1 0 33120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1666464484
transform -1 0 31832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0694_
timestamp 1666464484
transform -1 0 32660 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0695_
timestamp 1666464484
transform -1 0 31648 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0696_
timestamp 1666464484
transform -1 0 31740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0697_
timestamp 1666464484
transform 1 0 31464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0698_
timestamp 1666464484
transform -1 0 31556 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0699_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32568 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0700_
timestamp 1666464484
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1666464484
transform -1 0 33396 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1666464484
transform -1 0 33672 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0703_
timestamp 1666464484
transform -1 0 33212 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0704_
timestamp 1666464484
transform 1 0 33120 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _0705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0706_
timestamp 1666464484
transform -1 0 32200 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1666464484
transform 1 0 33580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0708_
timestamp 1666464484
transform 1 0 33488 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0709_
timestamp 1666464484
transform -1 0 30176 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28520 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ba_1  _0711_
timestamp 1666464484
transform 1 0 28336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1666464484
transform -1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32384 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_4  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28336 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_1  _0715_
timestamp 1666464484
transform -1 0 28152 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0717_
timestamp 1666464484
transform 1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0718_
timestamp 1666464484
transform -1 0 31188 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0719_
timestamp 1666464484
transform 1 0 28428 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1666464484
transform -1 0 27968 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0721_
timestamp 1666464484
transform -1 0 29348 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1666464484
transform -1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27508 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1666464484
transform 1 0 29716 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0725_
timestamp 1666464484
transform 1 0 30820 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0726_
timestamp 1666464484
transform -1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1666464484
transform -1 0 27508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _0728_
timestamp 1666464484
transform 1 0 14536 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0729_
timestamp 1666464484
transform 1 0 17756 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _0730_
timestamp 1666464484
transform 1 0 15916 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _0731_
timestamp 1666464484
transform 1 0 17572 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0732_
timestamp 1666464484
transform 1 0 15732 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0733_
timestamp 1666464484
transform 1 0 17664 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30360 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0735_
timestamp 1666464484
transform 1 0 17480 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0736_
timestamp 1666464484
transform 1 0 16836 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26312 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0738_
timestamp 1666464484
transform 1 0 17480 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0739_
timestamp 1666464484
transform -1 0 17112 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0740_
timestamp 1666464484
transform 1 0 17756 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0741_
timestamp 1666464484
transform 1 0 18768 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0742_
timestamp 1666464484
transform -1 0 22632 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0743_
timestamp 1666464484
transform 1 0 20608 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0744_
timestamp 1666464484
transform 1 0 17388 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0745_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0746_
timestamp 1666464484
transform 1 0 20516 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0747_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1666464484
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0749_
timestamp 1666464484
transform -1 0 25484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0750_
timestamp 1666464484
transform 1 0 24656 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0751_
timestamp 1666464484
transform 1 0 25300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0752_
timestamp 1666464484
transform 1 0 25852 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0754_
timestamp 1666464484
transform -1 0 14812 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_4  _0755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12788 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _0756_
timestamp 1666464484
transform 1 0 3220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0757_
timestamp 1666464484
transform -1 0 3496 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1666464484
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 1666464484
transform -1 0 12880 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0760_
timestamp 1666464484
transform 1 0 12052 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0761_
timestamp 1666464484
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1666464484
transform 1 0 12052 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0763_
timestamp 1666464484
transform -1 0 30360 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0764_
timestamp 1666464484
transform -1 0 28428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0765_
timestamp 1666464484
transform -1 0 28888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0767_
timestamp 1666464484
transform 1 0 27508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0768_
timestamp 1666464484
transform 1 0 18308 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0769_
timestamp 1666464484
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0770_
timestamp 1666464484
transform -1 0 25300 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0771_
timestamp 1666464484
transform 1 0 25024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1666464484
transform -1 0 28060 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0773_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0774_
timestamp 1666464484
transform 1 0 14260 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0775_
timestamp 1666464484
transform 1 0 12236 0 -1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1666464484
transform -1 0 3496 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0777_
timestamp 1666464484
transform 1 0 2668 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0778_
timestamp 1666464484
transform -1 0 4416 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0779_
timestamp 1666464484
transform -1 0 4416 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0780_
timestamp 1666464484
transform -1 0 15640 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0781_
timestamp 1666464484
transform -1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1666464484
transform -1 0 17572 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0783_
timestamp 1666464484
transform -1 0 16560 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 1666464484
transform -1 0 27784 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0785_
timestamp 1666464484
transform -1 0 28980 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1666464484
transform 1 0 20424 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1666464484
transform -1 0 23000 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0788_
timestamp 1666464484
transform 1 0 27232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0789_
timestamp 1666464484
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0790_
timestamp 1666464484
transform 1 0 27968 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0791_
timestamp 1666464484
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0792_
timestamp 1666464484
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0793_
timestamp 1666464484
transform -1 0 23460 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1666464484
transform 1 0 15088 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0795_
timestamp 1666464484
transform -1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0796_
timestamp 1666464484
transform 1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _0797_
timestamp 1666464484
transform 1 0 12420 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1666464484
transform -1 0 8648 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0799_
timestamp 1666464484
transform -1 0 8648 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_2  _0800_
timestamp 1666464484
transform -1 0 9476 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0801_
timestamp 1666464484
transform -1 0 6992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18676 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0803_
timestamp 1666464484
transform 1 0 17756 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0804_
timestamp 1666464484
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0805_
timestamp 1666464484
transform 1 0 28244 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0806_
timestamp 1666464484
transform -1 0 27876 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__a32o_1  _0807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0808_
timestamp 1666464484
transform -1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1666464484
transform 1 0 19412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0810_
timestamp 1666464484
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0811_
timestamp 1666464484
transform 1 0 23000 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0812_
timestamp 1666464484
transform -1 0 21160 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0813_
timestamp 1666464484
transform 1 0 19780 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _0814_
timestamp 1666464484
transform -1 0 20976 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1666464484
transform 1 0 11684 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _0816_
timestamp 1666464484
transform 1 0 12420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0817_
timestamp 1666464484
transform -1 0 11960 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1666464484
transform -1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1666464484
transform 1 0 10212 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0820_
timestamp 1666464484
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0821_
timestamp 1666464484
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0822_
timestamp 1666464484
transform 1 0 9108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0823_
timestamp 1666464484
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0824_
timestamp 1666464484
transform -1 0 8096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0825_
timestamp 1666464484
transform 1 0 5520 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1666464484
transform 1 0 6348 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0827_
timestamp 1666464484
transform -1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1666464484
transform -1 0 7912 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _0829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6808 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _0830_
timestamp 1666464484
transform 1 0 9844 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0831_
timestamp 1666464484
transform 1 0 4416 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _0832_
timestamp 1666464484
transform -1 0 5796 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0833_
timestamp 1666464484
transform -1 0 4692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1666464484
transform 1 0 2852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _0835_
timestamp 1666464484
transform -1 0 7636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _0836_
timestamp 1666464484
transform 1 0 6992 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 1666464484
transform 1 0 3128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1666464484
transform -1 0 7728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0839_
timestamp 1666464484
transform -1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0840_
timestamp 1666464484
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0841_
timestamp 1666464484
transform -1 0 10856 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0842_
timestamp 1666464484
transform 1 0 7636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0843_
timestamp 1666464484
transform 1 0 7176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1666464484
transform -1 0 8648 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1666464484
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0846_
timestamp 1666464484
transform -1 0 8556 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0847_
timestamp 1666464484
transform 1 0 6900 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0848_
timestamp 1666464484
transform 1 0 4140 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0849_
timestamp 1666464484
transform 1 0 3128 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0850_
timestamp 1666464484
transform 1 0 5060 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1666464484
transform -1 0 2392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0852_
timestamp 1666464484
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0853_
timestamp 1666464484
transform 1 0 5060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0856_
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0857_
timestamp 1666464484
transform -1 0 5520 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0858_
timestamp 1666464484
transform -1 0 3496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1666464484
transform 1 0 3956 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 1666464484
transform 1 0 3956 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _0862_
timestamp 1666464484
transform 1 0 3956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0863_
timestamp 1666464484
transform 1 0 4048 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1666464484
transform 1 0 6992 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0865_
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _0866_
timestamp 1666464484
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0867_
timestamp 1666464484
transform 1 0 8648 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _0868_
timestamp 1666464484
transform 1 0 9108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 1666464484
transform -1 0 3496 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0870_
timestamp 1666464484
transform -1 0 3496 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0871_
timestamp 1666464484
transform 1 0 20424 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0872_
timestamp 1666464484
transform 1 0 30820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0873_
timestamp 1666464484
transform 1 0 19412 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0874_
timestamp 1666464484
transform 1 0 23092 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0875_
timestamp 1666464484
transform 1 0 28704 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1666464484
transform 1 0 21988 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0877_
timestamp 1666464484
transform 1 0 19412 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0878_
timestamp 1666464484
transform 1 0 28612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0879_
timestamp 1666464484
transform 1 0 20608 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0880_
timestamp 1666464484
transform 1 0 22724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0881_
timestamp 1666464484
transform 1 0 25668 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0882_
timestamp 1666464484
transform 1 0 15548 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0883_
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0884_
timestamp 1666464484
transform 1 0 20424 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0885_
timestamp 1666464484
transform 1 0 14352 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0886_
timestamp 1666464484
transform -1 0 18952 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1666464484
transform -1 0 15916 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0888_
timestamp 1666464484
transform 1 0 25576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0889_
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0890_
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0891_
timestamp 1666464484
transform 1 0 11960 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1666464484
transform 1 0 28336 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 1666464484
transform -1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0895_
timestamp 1666464484
transform 1 0 29716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1666464484
transform 1 0 23552 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 1666464484
transform 1 0 17388 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1666464484
transform 1 0 17296 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1666464484
transform 1 0 16836 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1666464484
transform -1 0 29256 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0902_
timestamp 1666464484
transform 1 0 30452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1666464484
transform -1 0 29256 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1666464484
transform 1 0 29716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 1666464484
transform 1 0 22448 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1666464484
transform 1 0 21988 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1666464484
transform 1 0 17296 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1666464484
transform 1 0 20424 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1666464484
transform -1 0 31648 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0910_
timestamp 1666464484
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1666464484
transform -1 0 31832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1666464484
transform -1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0913_
timestamp 1666464484
transform -1 0 14904 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0914_
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0915_
timestamp 1666464484
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1666464484
transform 1 0 15732 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1666464484
transform -1 0 18952 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1666464484
transform 1 0 20424 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0919_
timestamp 1666464484
transform -1 0 19596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0920_
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1666464484
transform -1 0 26036 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1666464484
transform -1 0 25116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0923_
timestamp 1666464484
transform -1 0 26680 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0924_
timestamp 1666464484
transform -1 0 28336 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1666464484
transform -1 0 19964 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0926_
timestamp 1666464484
transform 1 0 20976 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1666464484
transform 1 0 23000 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0928_
timestamp 1666464484
transform 1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0929_
timestamp 1666464484
transform 1 0 26036 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1666464484
transform -1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0931_
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0932_
timestamp 1666464484
transform -1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1666464484
transform -1 0 30176 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1666464484
transform 1 0 32292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0935_
timestamp 1666464484
transform -1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1666464484
transform -1 0 31832 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1666464484
transform 1 0 23552 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1666464484
transform 1 0 23552 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0941_
timestamp 1666464484
transform 1 0 17664 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0942_
timestamp 1666464484
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0943_
timestamp 1666464484
transform -1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1666464484
transform 1 0 19412 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1666464484
transform 1 0 29900 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0946_
timestamp 1666464484
transform 1 0 32200 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1666464484
transform 1 0 32292 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0948_
timestamp 1666464484
transform 1 0 30544 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0949_
timestamp 1666464484
transform -1 0 21528 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0950_
timestamp 1666464484
transform 1 0 23276 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0951_
timestamp 1666464484
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0952_
timestamp 1666464484
transform -1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1666464484
transform -1 0 25116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0954_
timestamp 1666464484
transform 1 0 23552 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0956_
timestamp 1666464484
transform 1 0 3956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0957_
timestamp 1666464484
transform -1 0 3220 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1666464484
transform -1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0959_
timestamp 1666464484
transform -1 0 12144 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0960_
timestamp 1666464484
transform 1 0 9292 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0961_
timestamp 1666464484
transform 1 0 12144 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0962_
timestamp 1666464484
transform -1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0963_
timestamp 1666464484
transform 1 0 2944 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0964_
timestamp 1666464484
transform 1 0 7820 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0965_
timestamp 1666464484
transform -1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0966_
timestamp 1666464484
transform 1 0 9752 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0967_
timestamp 1666464484
transform 1 0 6992 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0968_
timestamp 1666464484
transform 1 0 9476 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0969_
timestamp 1666464484
transform -1 0 14536 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0970_
timestamp 1666464484
transform 1 0 12696 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0971_
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1666464484
transform -1 0 4416 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0973_
timestamp 1666464484
transform -1 0 5704 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0974__2
timestamp 1666464484
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975__3
timestamp 1666464484
transform -1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976__4
timestamp 1666464484
transform -1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977__5
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978__6
timestamp 1666464484
transform -1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979__7
timestamp 1666464484
transform -1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980__8
timestamp 1666464484
transform -1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1666464484
transform 1 0 24564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1666464484
transform 1 0 27416 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1666464484
transform 1 0 23828 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1666464484
transform -1 0 28796 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1666464484
transform 1 0 24564 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1666464484
transform 1 0 15548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1666464484
transform 1 0 16836 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1666464484
transform -1 0 16376 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1666464484
transform 1 0 14996 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1666464484
transform -1 0 29900 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1666464484
transform -1 0 29256 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1666464484
transform 1 0 30084 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1666464484
transform 1 0 28612 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1666464484
transform 1 0 21252 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1666464484
transform 1 0 19596 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1666464484
transform 1 0 19412 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1666464484
transform 1 0 19872 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1666464484
transform -1 0 32936 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1666464484
transform 1 0 32292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1666464484
transform 1 0 32292 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1666464484
transform -1 0 33764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1666464484
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1666464484
transform 1 0 15272 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1666464484
transform 1 0 14904 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1666464484
transform 1 0 15272 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_4  _1007_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1564 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1009_
timestamp 1666464484
transform 1 0 1656 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1010_
timestamp 1666464484
transform -1 0 12052 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1011_
timestamp 1666464484
transform -1 0 12144 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1012_
timestamp 1666464484
transform -1 0 13616 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1013_
timestamp 1666464484
transform -1 0 13156 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1014_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1666464484
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1666464484
transform 1 0 11684 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1666464484
transform 1 0 10764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1666464484
transform 1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1666464484
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1666464484
transform 1 0 11684 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1666464484
transform 1 0 11684 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1666464484
transform 1 0 5428 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1666464484
transform 1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1666464484
transform 1 0 11224 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1666464484
transform 1 0 10304 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1666464484
transform 1 0 5520 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1027_
timestamp 1666464484
transform 1 0 7084 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1028_
timestamp 1666464484
transform 1 0 9108 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1029_
timestamp 1666464484
transform 1 0 8924 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1030_
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1031_
timestamp 1666464484
transform 1 0 9108 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1032_
timestamp 1666464484
transform 1 0 11776 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1033_
timestamp 1666464484
transform 1 0 11776 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1034_
timestamp 1666464484
transform -1 0 9752 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  _1035_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2300 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1036_
timestamp 1666464484
transform 1 0 6808 0 -1 23936
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1037_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7084 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _1038_
timestamp 1666464484
transform 1 0 2668 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _1039_
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_2  _1040_
timestamp 1666464484
transform 1 0 4140 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1666464484
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1666464484
transform -1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1666464484
transform 1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1666464484
transform 1 0 16652 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1666464484
transform 1 0 17664 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1666464484
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1666464484
transform -1 0 21528 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1666464484
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1666464484
transform 1 0 19412 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1666464484
transform 1 0 19412 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1666464484
transform 1 0 18952 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1666464484
transform -1 0 26036 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1666464484
transform 1 0 24288 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1666464484
transform 1 0 25852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1666464484
transform 1 0 27140 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1666464484
transform 1 0 19688 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1666464484
transform 1 0 20056 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1666464484
transform 1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1666464484
transform 1 0 19688 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1666464484
transform 1 0 26404 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1666464484
transform 1 0 24564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1666464484
transform -1 0 25484 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1065_
timestamp 1666464484
transform -1 0 31464 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1066_
timestamp 1666464484
transform 1 0 31832 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1666464484
transform 1 0 32292 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1068_
timestamp 1666464484
transform 1 0 32292 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1069_
timestamp 1666464484
transform 1 0 23184 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1666464484
transform 1 0 23092 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1071_
timestamp 1666464484
transform 1 0 23184 0 -1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1072_
timestamp 1666464484
transform 1 0 23092 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1666464484
transform 1 0 17296 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1666464484
transform -1 0 18124 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1666464484
transform -1 0 18308 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1666464484
transform 1 0 17848 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1666464484
transform 1 0 29716 0 -1 27200
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1666464484
transform 1 0 29808 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1666464484
transform 1 0 30084 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1080_
timestamp 1666464484
transform 1 0 30084 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1081_
timestamp 1666464484
transform 1 0 21988 0 -1 25024
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1666464484
transform -1 0 21252 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1666464484
transform 1 0 21988 0 -1 26112
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1666464484
transform -1 0 25116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1666464484
transform -1 0 25024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 20240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 25116 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform 1 0 32292 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 23184 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform -1 0 19688 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 29992 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform 1 0 21620 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 24564 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 26036 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 21620 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 19228 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0460_
timestamp 1666464484
transform 1 0 20608 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1666464484
transform 1 0 15548 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform -1 0 33764 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 18216 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform -1 0 33028 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 20792 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform -1 0 17480 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 28612 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform -1 0 22632 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 23368 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform -1 0 25208 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform -1 0 14812 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform -1 0 30452 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 18216 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 18216 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0460_
timestamp 1666464484
transform -1 0 20056 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result
timestamp 1666464484
transform -1 0 33028 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result
timestamp 1666464484
transform 1 0 18216 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result
timestamp 1666464484
transform -1 0 25208 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result
timestamp 1666464484
transform -1 0 33028 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result
timestamp 1666464484
transform 1 0 20792 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result
timestamp 1666464484
transform 1 0 18216 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result
timestamp 1666464484
transform 1 0 28612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result
timestamp 1666464484
transform -1 0 22632 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result
timestamp 1666464484
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result
timestamp 1666464484
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result
timestamp 1666464484
transform 1 0 18216 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result
timestamp 1666464484
transform -1 0 30452 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result
timestamp 1666464484
transform 1 0 18216 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result
timestamp 1666464484
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result
timestamp 1666464484
transform 1 0 18216 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0460_
timestamp 1666464484
transform 1 0 20792 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1666464484
transform -1 0 9660 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1666464484
transform -1 0 12236 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1666464484
transform 1 0 20792 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20700 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout29
timestamp 1666464484
transform -1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout30
timestamp 1666464484
transform 1 0 21988 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27508 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout32
timestamp 1666464484
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout33
timestamp 1666464484
transform -1 0 22816 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout34
timestamp 1666464484
transform 1 0 17112 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  fanout35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 1666464484
transform -1 0 16376 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 1666464484
transform 1 0 14996 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1666464484
transform 1 0 19688 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout40
timestamp 1666464484
transform 1 0 16192 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1666464484
transform 1 0 18400 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp 1666464484
transform 1 0 18768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout43
timestamp 1666464484
transform -1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout44
timestamp 1666464484
transform 1 0 13984 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1666464484
transform -1 0 22540 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 1666464484
transform -1 0 12788 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 1666464484
transform -1 0 29808 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout49
timestamp 1666464484
transform 1 0 26128 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1666464484
transform -1 0 29992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout51
timestamp 1666464484
transform 1 0 26404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 1666464484
transform 1 0 13248 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  fanout53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout54
timestamp 1666464484
transform -1 0 4784 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout55
timestamp 1666464484
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout56
timestamp 1666464484
transform 1 0 12512 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1666464484
transform 1 0 7728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1666464484
transform 1 0 10672 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1666464484
transform -1 0 14628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform -1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1666464484
transform -1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform -1 0 22816 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1666464484
transform -1 0 25760 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1666464484
transform -1 0 28704 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1666464484
transform -1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1666464484
transform -1 0 34408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1666464484
transform 1 0 4784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output12
timestamp 1666464484
transform -1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp 1666464484
transform 1 0 15456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp 1666464484
transform 1 0 16836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp 1666464484
transform 1 0 18032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp 1666464484
transform 1 0 19412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output19
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp 1666464484
transform -1 0 25116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp 1666464484
transform -1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp 1666464484
transform -1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp 1666464484
transform -1 0 27692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp 1666464484
transform 1 0 28336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp 1666464484
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp 1666464484
transform -1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_58
timestamp 1666464484
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_59
timestamp 1666464484
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_60
timestamp 1666464484
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_61
timestamp 1666464484
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_62
timestamp 1666464484
transform -1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_63
timestamp 1666464484
transform -1 0 29992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_64
timestamp 1666464484
transform -1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_65
timestamp 1666464484
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_66
timestamp 1666464484
transform -1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_67
timestamp 1666464484
transform -1 0 34408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tholin_avalonsemi_5401_68
timestamp 1666464484
transform -1 0 34408 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 1766 35200 1822 36000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 7654 35200 7710 36000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 10598 35200 10654 36000 0 FreeSans 224 90 0 0 io_in[1]
port 2 nsew signal input
flabel metal2 s 13542 35200 13598 36000 0 FreeSans 224 90 0 0 io_in[2]
port 3 nsew signal input
flabel metal2 s 16486 35200 16542 36000 0 FreeSans 224 90 0 0 io_in[3]
port 4 nsew signal input
flabel metal2 s 19430 35200 19486 36000 0 FreeSans 224 90 0 0 io_in[4]
port 5 nsew signal input
flabel metal2 s 22374 35200 22430 36000 0 FreeSans 224 90 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 25318 35200 25374 36000 0 FreeSans 224 90 0 0 io_in[6]
port 7 nsew signal input
flabel metal2 s 28262 35200 28318 36000 0 FreeSans 224 90 0 0 io_in[7]
port 8 nsew signal input
flabel metal2 s 31206 35200 31262 36000 0 FreeSans 224 90 0 0 io_in[8]
port 9 nsew signal input
flabel metal2 s 34150 35200 34206 36000 0 FreeSans 224 90 0 0 io_in[9]
port 10 nsew signal input
flabel metal3 s 35200 17824 36000 17944 0 FreeSans 480 0 0 0 io_oeb
port 11 nsew signal tristate
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 io_out[0]
port 12 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 io_out[10]
port 13 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 io_out[11]
port 14 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[12]
port 15 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 io_out[13]
port 16 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 io_out[14]
port 17 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[15]
port 18 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 io_out[16]
port 19 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 io_out[17]
port 20 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[18]
port 21 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 io_out[19]
port 22 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 io_out[1]
port 23 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 io_out[20]
port 24 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_out[21]
port 25 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 io_out[22]
port 26 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 io_out[23]
port 27 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_out[24]
port 28 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 io_out[25]
port 29 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 io_out[26]
port 30 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal2 s 4710 35200 4766 36000 0 FreeSans 224 90 0 0 rst
port 39 nsew signal input
flabel metal4 s 5164 2128 5484 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 13605 2128 13925 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 22046 2128 22366 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 30487 2128 30807 33776 0 FreeSans 1920 90 0 0 vccd1
port 40 nsew power bidirectional
flabel metal4 s 9384 2128 9704 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 17825 2128 18145 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 26266 2128 26586 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
flabel metal4 s 34707 2128 35027 33776 0 FreeSans 1920 90 0 0 vssd1
port 41 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
