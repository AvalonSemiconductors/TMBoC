magic
tech sky130B
magscale 1 2
timestamp 1680006818
<< obsli1 >>
rect 1104 2159 83812 77809
<< obsm1 >>
rect 934 2128 83812 77840
<< metal2 >>
rect 4342 0 4398 800
rect 12806 0 12862 800
rect 21270 0 21326 800
rect 29734 0 29790 800
rect 38198 0 38254 800
rect 46662 0 46718 800
rect 55126 0 55182 800
rect 63590 0 63646 800
rect 72054 0 72110 800
rect 80518 0 80574 800
<< obsm2 >>
rect 938 856 83056 78577
rect 938 800 4286 856
rect 4454 800 12750 856
rect 12918 800 21214 856
rect 21382 800 29678 856
rect 29846 800 38142 856
rect 38310 800 46606 856
rect 46774 800 55070 856
rect 55238 800 63534 856
rect 63702 800 71998 856
rect 72166 800 80462 856
rect 80630 800 83056 856
<< metal3 >>
rect 0 78480 800 78600
rect 0 75624 800 75744
rect 0 72768 800 72888
rect 0 69912 800 70032
rect 0 67056 800 67176
rect 0 64200 800 64320
rect 0 61344 800 61464
rect 0 58488 800 58608
rect 0 55632 800 55752
rect 0 52776 800 52896
rect 0 49920 800 50040
rect 0 47064 800 47184
rect 0 44208 800 44328
rect 0 41352 800 41472
rect 0 38496 800 38616
rect 0 35640 800 35760
rect 0 32784 800 32904
rect 0 29928 800 30048
rect 0 27072 800 27192
rect 0 24216 800 24336
rect 0 21360 800 21480
rect 0 18504 800 18624
rect 0 15648 800 15768
rect 0 12792 800 12912
rect 0 9936 800 10056
rect 0 7080 800 7200
rect 0 4224 800 4344
rect 0 1368 800 1488
<< obsm3 >>
rect 880 78400 81326 78573
rect 800 75824 81326 78400
rect 880 75544 81326 75824
rect 800 72968 81326 75544
rect 880 72688 81326 72968
rect 800 70112 81326 72688
rect 880 69832 81326 70112
rect 800 67256 81326 69832
rect 880 66976 81326 67256
rect 800 64400 81326 66976
rect 880 64120 81326 64400
rect 800 61544 81326 64120
rect 880 61264 81326 61544
rect 800 58688 81326 61264
rect 880 58408 81326 58688
rect 800 55832 81326 58408
rect 880 55552 81326 55832
rect 800 52976 81326 55552
rect 880 52696 81326 52976
rect 800 50120 81326 52696
rect 880 49840 81326 50120
rect 800 47264 81326 49840
rect 880 46984 81326 47264
rect 800 44408 81326 46984
rect 880 44128 81326 44408
rect 800 41552 81326 44128
rect 880 41272 81326 41552
rect 800 38696 81326 41272
rect 880 38416 81326 38696
rect 800 35840 81326 38416
rect 880 35560 81326 35840
rect 800 32984 81326 35560
rect 880 32704 81326 32984
rect 800 30128 81326 32704
rect 880 29848 81326 30128
rect 800 27272 81326 29848
rect 880 26992 81326 27272
rect 800 24416 81326 26992
rect 880 24136 81326 24416
rect 800 21560 81326 24136
rect 880 21280 81326 21560
rect 800 18704 81326 21280
rect 880 18424 81326 18704
rect 800 15848 81326 18424
rect 880 15568 81326 15848
rect 800 12992 81326 15568
rect 880 12712 81326 12992
rect 800 10136 81326 12712
rect 880 9856 81326 10136
rect 800 7280 81326 9856
rect 880 7000 81326 7280
rect 800 4424 81326 7000
rect 880 4144 81326 4424
rect 800 1568 81326 4144
rect 880 1395 81326 1568
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
rect 81008 2128 81328 77840
<< obsm4 >>
rect 2267 11051 4128 63749
rect 4608 11051 19488 63749
rect 19968 11051 34848 63749
rect 35328 11051 50208 63749
rect 50688 11051 63605 63749
<< labels >>
rlabel metal2 s 72054 0 72110 800 6 clk
port 1 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 io_in[7]
port 9 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 io_oeb
port 10 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_out[10]
port 12 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 io_out[11]
port 13 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 io_out[12]
port 14 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_out[13]
port 15 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 io_out[14]
port 16 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_out[15]
port 17 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 io_out[16]
port 18 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 io_out[17]
port 19 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 io_out[18]
port 20 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_out[19]
port 21 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_out[1]
port 22 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 io_out[20]
port 23 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 io_out[21]
port 24 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 io_out[22]
port 25 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 io_out[23]
port 26 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_out[24]
port 27 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 io_out[25]
port 28 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 io_out[26]
port 29 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 io_out[2]
port 30 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 io_out[3]
port 31 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 io_out[4]
port 32 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_out[5]
port 33 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 io_out[6]
port 34 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_out[7]
port 35 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 io_out[8]
port 36 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 io_out[9]
port 37 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 rst
port 38 nsew signal input
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 40 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 77840 6 vssd1
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 85000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15615394
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS2650/runs/23_03_28_14_27/results/signoff/wrapped_as2650.magic.gds
string GDS_START 1381514
<< end >>

