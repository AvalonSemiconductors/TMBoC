magic
tech sky130B
magscale 1 2
timestamp 1680517358
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 429838 700748 429844 700800
rect 429896 700788 429902 700800
rect 449158 700788 449164 700800
rect 429896 700760 449164 700788
rect 429896 700748 429902 700760
rect 449158 700748 449164 700760
rect 449216 700748 449222 700800
rect 364978 700680 364984 700732
rect 365036 700720 365042 700732
rect 445018 700720 445024 700732
rect 365036 700692 445024 700720
rect 365036 700680 365042 700692
rect 445018 700680 445024 700692
rect 445076 700680 445082 700732
rect 348786 700612 348792 700664
rect 348844 700652 348850 700664
rect 446398 700652 446404 700664
rect 348844 700624 446404 700652
rect 348844 700612 348850 700624
rect 446398 700612 446404 700624
rect 446456 700612 446462 700664
rect 235166 700544 235172 700596
rect 235224 700584 235230 700596
rect 450538 700584 450544 700596
rect 235224 700556 450544 700584
rect 235224 700544 235230 700556
rect 450538 700544 450544 700556
rect 450596 700544 450602 700596
rect 218974 700476 218980 700528
rect 219032 700516 219038 700528
rect 449250 700516 449256 700528
rect 219032 700488 449256 700516
rect 219032 700476 219038 700488
rect 449250 700476 449256 700488
rect 449308 700476 449314 700528
rect 170306 700408 170312 700460
rect 170364 700448 170370 700460
rect 444282 700448 444288 700460
rect 170364 700420 444288 700448
rect 170364 700408 170370 700420
rect 444282 700408 444288 700420
rect 444340 700408 444346 700460
rect 105446 700340 105452 700392
rect 105504 700380 105510 700392
rect 445110 700380 445116 700392
rect 105504 700352 445116 700380
rect 105504 700340 105510 700352
rect 445110 700340 445116 700352
rect 445168 700340 445174 700392
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 445202 700312 445208 700324
rect 73028 700284 445208 700312
rect 73028 700272 73034 700284
rect 445202 700272 445208 700284
rect 445260 700272 445266 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 573358 696940 573364 696992
rect 573416 696980 573422 696992
rect 580166 696980 580172 696992
rect 573416 696952 580172 696980
rect 573416 696940 573422 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 299474 687896 299480 687948
rect 299532 687936 299538 687948
rect 449342 687936 449348 687948
rect 299532 687908 449348 687936
rect 299532 687896 299538 687908
rect 449342 687896 449348 687908
rect 449400 687896 449406 687948
rect 266354 686468 266360 686520
rect 266412 686508 266418 686520
rect 446490 686508 446496 686520
rect 266412 686480 446496 686508
rect 266412 686468 266418 686480
rect 446490 686468 446496 686480
rect 446548 686468 446554 686520
rect 88334 685244 88340 685296
rect 88392 685284 88398 685296
rect 418798 685284 418804 685296
rect 88392 685256 418804 685284
rect 88392 685244 88398 685256
rect 418798 685244 418804 685256
rect 418856 685244 418862 685296
rect 23474 685176 23480 685228
rect 23532 685216 23538 685228
rect 446582 685216 446588 685228
rect 23532 685188 446588 685216
rect 23532 685176 23538 685188
rect 446582 685176 446588 685188
rect 446640 685176 446646 685228
rect 6914 685108 6920 685160
rect 6972 685148 6978 685160
rect 446766 685148 446772 685160
rect 6972 685120 446772 685148
rect 6972 685108 6978 685120
rect 446766 685108 446772 685120
rect 446824 685108 446830 685160
rect 3970 684700 3976 684752
rect 4028 684740 4034 684752
rect 420362 684740 420368 684752
rect 4028 684712 420368 684740
rect 4028 684700 4034 684712
rect 420362 684700 420368 684712
rect 420420 684700 420426 684752
rect 3142 684632 3148 684684
rect 3200 684672 3206 684684
rect 420178 684672 420184 684684
rect 3200 684644 420184 684672
rect 3200 684632 3206 684644
rect 420178 684632 420184 684644
rect 420236 684632 420242 684684
rect 3326 684564 3332 684616
rect 3384 684604 3390 684616
rect 420546 684604 420552 684616
rect 3384 684576 420552 684604
rect 3384 684564 3390 684576
rect 420546 684564 420552 684576
rect 420604 684564 420610 684616
rect 3878 684496 3884 684548
rect 3936 684536 3942 684548
rect 446950 684536 446956 684548
rect 3936 684508 446956 684536
rect 3936 684496 3942 684508
rect 446950 684496 446956 684508
rect 447008 684496 447014 684548
rect 331214 683748 331220 683800
rect 331272 683788 331278 683800
rect 418890 683788 418896 683800
rect 331272 683760 418896 683788
rect 331272 683748 331278 683760
rect 418890 683748 418896 683760
rect 418948 683748 418954 683800
rect 20898 683544 20904 683596
rect 20956 683584 20962 683596
rect 359458 683584 359464 683596
rect 20956 683556 359464 683584
rect 20956 683544 20962 683556
rect 359458 683544 359464 683556
rect 359516 683544 359522 683596
rect 19978 683476 19984 683528
rect 20036 683516 20042 683528
rect 417418 683516 417424 683528
rect 20036 683488 417424 683516
rect 20036 683476 20042 683488
rect 417418 683476 417424 683488
rect 417476 683476 417482 683528
rect 4062 683408 4068 683460
rect 4120 683448 4126 683460
rect 420730 683448 420736 683460
rect 4120 683420 420736 683448
rect 4120 683408 4126 683420
rect 420730 683408 420736 683420
rect 420788 683408 420794 683460
rect 3786 683340 3792 683392
rect 3844 683380 3850 683392
rect 420638 683380 420644 683392
rect 3844 683352 420644 683380
rect 3844 683340 3850 683352
rect 420638 683340 420644 683352
rect 420696 683340 420702 683392
rect 3694 683272 3700 683324
rect 3752 683312 3758 683324
rect 445294 683312 445300 683324
rect 3752 683284 445300 683312
rect 3752 683272 3758 683284
rect 445294 683272 445300 683284
rect 445352 683272 445358 683324
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 445478 683244 445484 683256
rect 3476 683216 445484 683244
rect 3476 683204 3482 683216
rect 445478 683204 445484 683216
rect 445536 683204 445542 683256
rect 3510 683136 3516 683188
rect 3568 683176 3574 683188
rect 446674 683176 446680 683188
rect 3568 683148 446680 683176
rect 3568 683136 3574 683148
rect 446674 683136 446680 683148
rect 446732 683136 446738 683188
rect 576118 683136 576124 683188
rect 576176 683176 576182 683188
rect 580166 683176 580172 683188
rect 576176 683148 580172 683176
rect 576176 683136 576182 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 2866 682728 2872 682780
rect 2924 682768 2930 682780
rect 420822 682768 420828 682780
rect 2924 682740 420828 682768
rect 2924 682728 2930 682740
rect 420822 682728 420828 682740
rect 420880 682728 420886 682780
rect 2958 682660 2964 682712
rect 3016 682700 3022 682712
rect 447042 682700 447048 682712
rect 3016 682672 447048 682700
rect 3016 682660 3022 682672
rect 447042 682660 447048 682672
rect 447100 682660 447106 682712
rect 18138 680348 18144 680400
rect 18196 680388 18202 680400
rect 20898 680388 20904 680400
rect 18196 680360 20904 680388
rect 18196 680348 18202 680360
rect 20898 680348 20904 680360
rect 20956 680348 20962 680400
rect 361758 678988 361764 679040
rect 361816 679028 361822 679040
rect 382918 679028 382924 679040
rect 361816 679000 382924 679028
rect 361816 678988 361822 679000
rect 382918 678988 382924 679000
rect 382976 678988 382982 679040
rect 3510 678512 3516 678564
rect 3568 678512 3574 678564
rect 3528 678360 3556 678512
rect 3510 678308 3516 678360
rect 3568 678308 3574 678360
rect 16574 675248 16580 675300
rect 16632 675288 16638 675300
rect 18138 675288 18144 675300
rect 16632 675260 18144 675288
rect 16632 675248 16638 675260
rect 18138 675248 18144 675260
rect 18196 675248 18202 675300
rect 567838 670692 567844 670744
rect 567896 670732 567902 670744
rect 580166 670732 580172 670744
rect 567896 670704 580172 670732
rect 567896 670692 567902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 13078 667904 13084 667956
rect 13136 667944 13142 667956
rect 16482 667944 16488 667956
rect 13136 667916 16488 667944
rect 13136 667904 13142 667916
rect 16482 667904 16488 667916
rect 16540 667904 16546 667956
rect 361758 667904 361764 667956
rect 361816 667944 361822 667956
rect 378778 667944 378784 667956
rect 361816 667916 378784 667944
rect 361816 667904 361822 667916
rect 378778 667904 378784 667916
rect 378836 667904 378842 667956
rect 8938 662396 8944 662448
rect 8996 662436 9002 662448
rect 13078 662436 13084 662448
rect 8996 662408 13084 662436
rect 8996 662396 9002 662408
rect 13078 662396 13084 662408
rect 13136 662396 13142 662448
rect 361758 656888 361764 656940
rect 361816 656928 361822 656940
rect 400858 656928 400864 656940
rect 361816 656900 400864 656928
rect 361816 656888 361822 656900
rect 400858 656888 400864 656900
rect 400916 656888 400922 656940
rect 8938 652780 8944 652792
rect 6886 652752 8944 652780
rect 4798 652672 4804 652724
rect 4856 652712 4862 652724
rect 6886 652712 6914 652752
rect 8938 652740 8944 652752
rect 8996 652740 9002 652792
rect 4856 652684 6914 652712
rect 4856 652672 4862 652684
rect 361758 645872 361764 645924
rect 361816 645912 361822 645924
rect 376018 645912 376024 645924
rect 361816 645884 376024 645912
rect 361816 645872 361822 645884
rect 376018 645872 376024 645884
rect 376076 645872 376082 645924
rect 361574 634788 361580 634840
rect 361632 634828 361638 634840
rect 403618 634828 403624 634840
rect 361632 634800 403624 634828
rect 361632 634788 361638 634800
rect 403618 634788 403624 634800
rect 403676 634788 403682 634840
rect 3694 631320 3700 631372
rect 3752 631360 3758 631372
rect 19978 631360 19984 631372
rect 3752 631332 19984 631360
rect 3752 631320 3758 631332
rect 19978 631320 19984 631332
rect 20036 631320 20042 631372
rect 574738 630640 574744 630692
rect 574796 630680 574802 630692
rect 580166 630680 580172 630692
rect 574796 630652 580172 630680
rect 574796 630640 574802 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 361574 623772 361580 623824
rect 361632 623812 361638 623824
rect 374638 623812 374644 623824
rect 361632 623784 374644 623812
rect 361632 623772 361638 623784
rect 374638 623772 374644 623784
rect 374696 623772 374702 623824
rect 361574 612756 361580 612808
rect 361632 612796 361638 612808
rect 406378 612796 406384 612808
rect 361632 612768 406384 612796
rect 361632 612756 361638 612768
rect 406378 612756 406384 612768
rect 406436 612756 406442 612808
rect 359458 609968 359464 610020
rect 359516 610008 359522 610020
rect 359516 609980 361620 610008
rect 359516 609968 359522 609980
rect 361592 609940 361620 609980
rect 365714 609940 365720 609952
rect 361592 609912 365720 609940
rect 365714 609900 365720 609912
rect 365772 609900 365778 609952
rect 365714 607112 365720 607164
rect 365772 607152 365778 607164
rect 367830 607152 367836 607164
rect 365772 607124 367836 607152
rect 365772 607112 365778 607124
rect 367830 607112 367836 607124
rect 367888 607112 367894 607164
rect 458726 602760 458732 602812
rect 458784 602800 458790 602812
rect 459094 602800 459100 602812
rect 458784 602772 459100 602800
rect 458784 602760 458790 602772
rect 459094 602760 459100 602772
rect 459152 602760 459158 602812
rect 361574 601740 361580 601792
rect 361632 601780 361638 601792
rect 371878 601780 371884 601792
rect 361632 601752 371884 601780
rect 361632 601740 361638 601752
rect 371878 601740 371884 601752
rect 371936 601740 371942 601792
rect 367830 601672 367836 601724
rect 367888 601712 367894 601724
rect 369118 601712 369124 601724
rect 367888 601684 369124 601712
rect 367888 601672 367894 601684
rect 369118 601672 369124 601684
rect 369176 601672 369182 601724
rect 457806 600244 457812 600296
rect 457864 600284 457870 600296
rect 461670 600284 461676 600296
rect 457864 600256 461676 600284
rect 457864 600244 457870 600256
rect 461670 600244 461676 600256
rect 461728 600244 461734 600296
rect 457530 600176 457536 600228
rect 457588 600216 457594 600228
rect 461578 600216 461584 600228
rect 457588 600188 461584 600216
rect 457588 600176 457594 600188
rect 461578 600176 461584 600188
rect 461636 600176 461642 600228
rect 459186 599972 459192 600024
rect 459244 600012 459250 600024
rect 462498 600012 462504 600024
rect 459244 599984 462504 600012
rect 459244 599972 459250 599984
rect 462498 599972 462504 599984
rect 462556 599972 462562 600024
rect 458634 599700 458640 599752
rect 458692 599740 458698 599752
rect 465074 599740 465080 599752
rect 458692 599712 465080 599740
rect 458692 599700 458698 599712
rect 465074 599700 465080 599712
rect 465132 599700 465138 599752
rect 457254 599632 457260 599684
rect 457312 599672 457318 599684
rect 465166 599672 465172 599684
rect 457312 599644 465172 599672
rect 457312 599632 457318 599644
rect 465166 599632 465172 599644
rect 465224 599632 465230 599684
rect 457898 599564 457904 599616
rect 457956 599604 457962 599616
rect 468478 599604 468484 599616
rect 457956 599576 468484 599604
rect 457956 599564 457962 599576
rect 468478 599564 468484 599576
rect 468536 599564 468542 599616
rect 515398 599564 515404 599616
rect 515456 599604 515462 599616
rect 580350 599604 580356 599616
rect 515456 599576 580356 599604
rect 515456 599564 515462 599576
rect 580350 599564 580356 599576
rect 580408 599564 580414 599616
rect 459830 598408 459836 598460
rect 459888 598448 459894 598460
rect 463694 598448 463700 598460
rect 459888 598420 463700 598448
rect 459888 598408 459894 598420
rect 463694 598408 463700 598420
rect 463752 598408 463758 598460
rect 458818 598340 458824 598392
rect 458876 598380 458882 598392
rect 467926 598380 467932 598392
rect 458876 598352 467932 598380
rect 458876 598340 458882 598352
rect 467926 598340 467932 598352
rect 467984 598340 467990 598392
rect 484486 598340 484492 598392
rect 484544 598380 484550 598392
rect 494146 598380 494152 598392
rect 484544 598352 494152 598380
rect 484544 598340 484550 598352
rect 494146 598340 494152 598352
rect 494204 598340 494210 598392
rect 457622 598272 457628 598324
rect 457680 598312 457686 598324
rect 468570 598312 468576 598324
rect 457680 598284 468576 598312
rect 457680 598272 457686 598284
rect 468570 598272 468576 598284
rect 468628 598272 468634 598324
rect 477494 598272 477500 598324
rect 477552 598312 477558 598324
rect 494054 598312 494060 598324
rect 477552 598284 494060 598312
rect 477552 598272 477558 598284
rect 494054 598272 494060 598284
rect 494112 598272 494118 598324
rect 447962 598204 447968 598256
rect 448020 598244 448026 598256
rect 505462 598244 505468 598256
rect 448020 598216 505468 598244
rect 448020 598204 448026 598216
rect 505462 598204 505468 598216
rect 505520 598204 505526 598256
rect 491478 597796 491484 597848
rect 491536 597836 491542 597848
rect 494238 597836 494244 597848
rect 491536 597808 494244 597836
rect 491536 597796 491542 597808
rect 494238 597796 494244 597808
rect 494296 597796 494302 597848
rect 459738 596844 459744 596896
rect 459796 596884 459802 596896
rect 463786 596884 463792 596896
rect 459796 596856 463792 596884
rect 459796 596844 459802 596856
rect 463786 596844 463792 596856
rect 463844 596844 463850 596896
rect 457714 596572 457720 596624
rect 457772 596612 457778 596624
rect 461762 596612 461768 596624
rect 457772 596584 461768 596612
rect 457772 596572 457778 596584
rect 461762 596572 461768 596584
rect 461820 596572 461826 596624
rect 457438 595484 457444 595536
rect 457496 595524 457502 595536
rect 464338 595524 464344 595536
rect 457496 595496 464344 595524
rect 457496 595484 457502 595496
rect 464338 595484 464344 595496
rect 464396 595484 464402 595536
rect 449802 595416 449808 595468
rect 449860 595456 449866 595468
rect 469214 595456 469220 595468
rect 449860 595428 469220 595456
rect 449860 595416 449866 595428
rect 469214 595416 469220 595428
rect 469272 595416 469278 595468
rect 369118 595348 369124 595400
rect 369176 595388 369182 595400
rect 370682 595388 370688 595400
rect 369176 595360 370688 595388
rect 369176 595348 369182 595360
rect 370682 595348 370688 595360
rect 370740 595348 370746 595400
rect 459646 594056 459652 594108
rect 459704 594096 459710 594108
rect 466454 594096 466460 594108
rect 459704 594068 466460 594096
rect 459704 594056 459710 594068
rect 466454 594056 466460 594068
rect 466512 594056 466518 594108
rect 370682 593308 370688 593360
rect 370740 593348 370746 593360
rect 372614 593348 372620 593360
rect 370740 593320 372620 593348
rect 370740 593308 370746 593320
rect 372614 593308 372620 593320
rect 372672 593308 372678 593360
rect 361758 590656 361764 590708
rect 361816 590696 361822 590708
rect 370682 590696 370688 590708
rect 361816 590668 370688 590696
rect 361816 590656 361822 590668
rect 370682 590656 370688 590668
rect 370740 590656 370746 590708
rect 511258 590656 511264 590708
rect 511316 590696 511322 590708
rect 580166 590696 580172 590708
rect 511316 590668 580172 590696
rect 511316 590656 511322 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 372614 590588 372620 590640
rect 372672 590628 372678 590640
rect 376110 590628 376116 590640
rect 372672 590600 376116 590628
rect 372672 590588 372678 590600
rect 376110 590588 376116 590600
rect 376168 590588 376174 590640
rect 376110 582360 376116 582412
rect 376168 582400 376174 582412
rect 378870 582400 378876 582412
rect 376168 582372 378876 582400
rect 376168 582360 376174 582372
rect 378870 582360 378876 582372
rect 378928 582360 378934 582412
rect 361758 579640 361764 579692
rect 361816 579680 361822 579692
rect 367738 579680 367744 579692
rect 361816 579652 367744 579680
rect 361816 579640 361822 579652
rect 367738 579640 367744 579652
rect 367796 579640 367802 579692
rect 378870 574948 378876 575000
rect 378928 574988 378934 575000
rect 380802 574988 380808 575000
rect 378928 574960 380808 574988
rect 378928 574948 378934 574960
rect 380802 574948 380808 574960
rect 380860 574948 380866 575000
rect 380802 571344 380808 571396
rect 380860 571384 380866 571396
rect 380860 571356 380940 571384
rect 380860 571344 380866 571356
rect 380912 571316 380940 571356
rect 385678 571316 385684 571328
rect 380912 571288 385684 571316
rect 385678 571276 385684 571288
rect 385736 571276 385742 571328
rect 361574 568760 361580 568812
rect 361632 568800 361638 568812
rect 363598 568800 363604 568812
rect 361632 568772 363604 568800
rect 361632 568760 361638 568772
rect 363598 568760 363604 568772
rect 363656 568760 363662 568812
rect 515490 563048 515496 563100
rect 515548 563088 515554 563100
rect 579890 563088 579896 563100
rect 515548 563060 579896 563088
rect 515548 563048 515554 563060
rect 579890 563048 579896 563060
rect 579948 563048 579954 563100
rect 385678 560192 385684 560244
rect 385736 560232 385742 560244
rect 387150 560232 387156 560244
rect 385736 560204 387156 560232
rect 385736 560192 385742 560204
rect 387150 560192 387156 560204
rect 387208 560192 387214 560244
rect 361574 557744 361580 557796
rect 361632 557784 361638 557796
rect 363690 557784 363696 557796
rect 361632 557756 363696 557784
rect 361632 557744 361638 557756
rect 363690 557744 363696 557756
rect 363748 557744 363754 557796
rect 387150 556180 387156 556232
rect 387208 556220 387214 556232
rect 388438 556220 388444 556232
rect 387208 556192 388444 556220
rect 387208 556180 387214 556192
rect 388438 556180 388444 556192
rect 388496 556180 388502 556232
rect 361758 546456 361764 546508
rect 361816 546496 361822 546508
rect 407758 546496 407764 546508
rect 361816 546468 407764 546496
rect 361816 546456 361822 546468
rect 407758 546456 407764 546468
rect 407816 546456 407822 546508
rect 457346 542988 457352 543040
rect 457404 543028 457410 543040
rect 466546 543028 466552 543040
rect 457404 543000 466552 543028
rect 457404 542988 457410 543000
rect 466546 542988 466552 543000
rect 466604 542988 466610 543040
rect 514018 536800 514024 536852
rect 514076 536840 514082 536852
rect 580166 536840 580172 536852
rect 514076 536812 580172 536840
rect 514076 536800 514082 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 459554 536052 459560 536104
rect 459612 536092 459618 536104
rect 469398 536092 469404 536104
rect 459612 536064 469404 536092
rect 459612 536052 459618 536064
rect 469398 536052 469404 536064
rect 469456 536052 469462 536104
rect 361758 535440 361764 535492
rect 361816 535480 361822 535492
rect 410518 535480 410524 535492
rect 361816 535452 410524 535480
rect 361816 535440 361822 535452
rect 410518 535440 410524 535452
rect 410576 535440 410582 535492
rect 361758 524424 361764 524476
rect 361816 524464 361822 524476
rect 411898 524464 411904 524476
rect 361816 524436 411904 524464
rect 361816 524424 361822 524436
rect 411898 524424 411904 524436
rect 411956 524424 411962 524476
rect 457990 523676 457996 523728
rect 458048 523716 458054 523728
rect 467098 523716 467104 523728
rect 458048 523688 467104 523716
rect 458048 523676 458054 523688
rect 467098 523676 467104 523688
rect 467156 523676 467162 523728
rect 388438 522928 388444 522980
rect 388496 522968 388502 522980
rect 389818 522968 389824 522980
rect 388496 522940 389824 522968
rect 388496 522928 388502 522940
rect 389818 522928 389824 522940
rect 389876 522928 389882 522980
rect 458082 522316 458088 522368
rect 458140 522356 458146 522368
rect 468662 522356 468668 522368
rect 458140 522328 468668 522356
rect 458140 522316 458146 522328
rect 468662 522316 468668 522328
rect 468720 522316 468726 522368
rect 448054 522248 448060 522300
rect 448112 522288 448118 522300
rect 462406 522288 462412 522300
rect 448112 522260 462412 522288
rect 448112 522248 448118 522260
rect 462406 522248 462412 522260
rect 462464 522248 462470 522300
rect 459278 520888 459284 520940
rect 459336 520928 459342 520940
rect 470870 520928 470876 520940
rect 459336 520900 470876 520928
rect 459336 520888 459342 520900
rect 470870 520888 470876 520900
rect 470928 520888 470934 520940
rect 482922 520888 482928 520940
rect 482980 520928 482986 520940
rect 518894 520928 518900 520940
rect 482980 520900 518900 520928
rect 482980 520888 482986 520900
rect 518894 520888 518900 520900
rect 518952 520888 518958 520940
rect 449986 520344 449992 520396
rect 450044 520384 450050 520396
rect 488626 520384 488632 520396
rect 450044 520356 488632 520384
rect 450044 520344 450050 520356
rect 488626 520344 488632 520356
rect 488684 520344 488690 520396
rect 389818 520208 389824 520260
rect 389876 520248 389882 520260
rect 391198 520248 391204 520260
rect 389876 520220 391204 520248
rect 389876 520208 389882 520220
rect 391198 520208 391204 520220
rect 391256 520208 391262 520260
rect 450630 519528 450636 519580
rect 450688 519568 450694 519580
rect 511994 519568 512000 519580
rect 450688 519540 512000 519568
rect 450688 519528 450694 519540
rect 511994 519528 512000 519540
rect 512052 519528 512058 519580
rect 459370 518236 459376 518288
rect 459428 518276 459434 518288
rect 470686 518276 470692 518288
rect 459428 518248 470692 518276
rect 459428 518236 459434 518248
rect 470686 518236 470692 518248
rect 470744 518236 470750 518288
rect 448330 518168 448336 518220
rect 448388 518208 448394 518220
rect 498194 518208 498200 518220
rect 448388 518180 498200 518208
rect 448388 518168 448394 518180
rect 498194 518168 498200 518180
rect 498252 518168 498258 518220
rect 480162 517488 480168 517540
rect 480220 517528 480226 517540
rect 482646 517528 482652 517540
rect 480220 517500 482652 517528
rect 480220 517488 480226 517500
rect 482646 517488 482652 517500
rect 482704 517488 482710 517540
rect 448422 516128 448428 516180
rect 448480 516168 448486 516180
rect 491846 516168 491852 516180
rect 448480 516140 491852 516168
rect 448480 516128 448486 516140
rect 491846 516128 491852 516140
rect 491904 516128 491910 516180
rect 494146 515380 494152 515432
rect 494204 515420 494210 515432
rect 538214 515420 538220 515432
rect 494204 515392 538220 515420
rect 494204 515380 494210 515392
rect 538214 515380 538220 515392
rect 538272 515380 538278 515432
rect 3970 514768 3976 514820
rect 4028 514808 4034 514820
rect 4798 514808 4804 514820
rect 4028 514780 4804 514808
rect 4028 514768 4034 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 361758 513340 361764 513392
rect 361816 513380 361822 513392
rect 414658 513380 414664 513392
rect 361816 513352 414664 513380
rect 361816 513340 361822 513352
rect 414658 513340 414664 513352
rect 414716 513340 414722 513392
rect 494146 512592 494152 512644
rect 494204 512632 494210 512644
rect 494330 512632 494336 512644
rect 494204 512604 494336 512632
rect 494204 512592 494210 512604
rect 494330 512592 494336 512604
rect 494388 512632 494394 512644
rect 535454 512632 535460 512644
rect 494388 512604 535460 512632
rect 494388 512592 494394 512604
rect 535454 512592 535460 512604
rect 535512 512592 535518 512644
rect 494054 507832 494060 507884
rect 494112 507872 494118 507884
rect 532694 507872 532700 507884
rect 494112 507844 532700 507872
rect 494112 507832 494118 507844
rect 532694 507832 532700 507844
rect 532752 507832 532758 507884
rect 494238 505112 494244 505164
rect 494296 505152 494302 505164
rect 529934 505152 529940 505164
rect 494296 505124 529940 505152
rect 494296 505112 494302 505124
rect 529934 505112 529940 505124
rect 529992 505112 529998 505164
rect 361758 502324 361764 502376
rect 361816 502364 361822 502376
rect 416038 502364 416044 502376
rect 361816 502336 416044 502364
rect 361816 502324 361822 502336
rect 416038 502324 416044 502336
rect 416096 502324 416102 502376
rect 448054 501780 448060 501832
rect 448112 501820 448118 501832
rect 448330 501820 448336 501832
rect 448112 501792 448336 501820
rect 448112 501780 448118 501792
rect 448330 501780 448336 501792
rect 448388 501780 448394 501832
rect 391198 500556 391204 500608
rect 391256 500596 391262 500608
rect 393406 500596 393412 500608
rect 391256 500568 393412 500596
rect 391256 500556 391262 500568
rect 393406 500556 393412 500568
rect 393464 500556 393470 500608
rect 448514 500216 448520 500268
rect 448572 500256 448578 500268
rect 545114 500256 545120 500268
rect 448572 500228 545120 500256
rect 448572 500216 448578 500228
rect 545114 500216 545120 500228
rect 545172 500216 545178 500268
rect 447410 499536 447416 499588
rect 447468 499576 447474 499588
rect 449710 499576 449716 499588
rect 447468 499548 449716 499576
rect 447468 499536 447474 499548
rect 449710 499536 449716 499548
rect 449768 499536 449774 499588
rect 447962 499468 447968 499520
rect 448020 499508 448026 499520
rect 494054 499508 494060 499520
rect 448020 499480 494060 499508
rect 448020 499468 448026 499480
rect 494054 499468 494060 499480
rect 494112 499468 494118 499520
rect 448054 499400 448060 499452
rect 448112 499440 448118 499452
rect 494238 499440 494244 499452
rect 448112 499412 494244 499440
rect 448112 499400 448118 499412
rect 494238 499400 494244 499412
rect 494296 499400 494302 499452
rect 449710 498788 449716 498840
rect 449768 498828 449774 498840
rect 542446 498828 542452 498840
rect 449768 498800 542452 498828
rect 449768 498788 449774 498800
rect 542446 498788 542452 498800
rect 542504 498788 542510 498840
rect 457438 497564 457444 497616
rect 457496 497604 457502 497616
rect 482646 497604 482652 497616
rect 457496 497576 482652 497604
rect 457496 497564 457502 497576
rect 482646 497564 482652 497576
rect 482704 497564 482710 497616
rect 453298 497496 453304 497548
rect 453356 497536 453362 497548
rect 480254 497536 480260 497548
rect 453356 497508 480260 497536
rect 453356 497496 453362 497508
rect 480254 497496 480260 497508
rect 480312 497496 480318 497548
rect 451918 497428 451924 497480
rect 451976 497468 451982 497480
rect 491294 497468 491300 497480
rect 451976 497440 491300 497468
rect 451976 497428 451982 497440
rect 491294 497428 491300 497440
rect 491352 497428 491358 497480
rect 454126 497020 454132 497072
rect 454184 497060 454190 497072
rect 459554 497060 459560 497072
rect 454184 497032 459560 497060
rect 454184 497020 454190 497032
rect 459554 497020 459560 497032
rect 459612 497020 459618 497072
rect 454034 496952 454040 497004
rect 454092 496992 454098 497004
rect 458082 496992 458088 497004
rect 454092 496964 458088 496992
rect 454092 496952 454098 496964
rect 458082 496952 458088 496964
rect 458140 496952 458146 497004
rect 452838 496884 452844 496936
rect 452896 496924 452902 496936
rect 455138 496924 455144 496936
rect 452896 496896 455144 496924
rect 452896 496884 452902 496896
rect 455138 496884 455144 496896
rect 455196 496884 455202 496936
rect 455414 496884 455420 496936
rect 455472 496924 455478 496936
rect 461026 496924 461032 496936
rect 455472 496896 461032 496924
rect 455472 496884 455478 496896
rect 461026 496884 461032 496896
rect 461084 496884 461090 496936
rect 451366 496816 451372 496868
rect 451424 496856 451430 496868
rect 453666 496856 453672 496868
rect 451424 496828 453672 496856
rect 451424 496816 451430 496828
rect 453666 496816 453672 496828
rect 453724 496816 453730 496868
rect 454678 496816 454684 496868
rect 454736 496856 454742 496868
rect 456610 496856 456616 496868
rect 454736 496828 456616 496856
rect 454736 496816 454742 496828
rect 456610 496816 456616 496828
rect 456668 496816 456674 496868
rect 393406 496204 393412 496256
rect 393464 496244 393470 496256
rect 397546 496244 397552 496256
rect 393464 496216 397552 496244
rect 393464 496204 393470 496216
rect 397546 496204 397552 496216
rect 397604 496204 397610 496256
rect 449894 496068 449900 496120
rect 449952 496108 449958 496120
rect 547874 496108 547880 496120
rect 449952 496080 547880 496108
rect 449952 496068 449958 496080
rect 547874 496068 547880 496080
rect 547932 496068 547938 496120
rect 449894 494708 449900 494760
rect 449952 494748 449958 494760
rect 450630 494748 450636 494760
rect 449952 494720 450636 494748
rect 449952 494708 449958 494720
rect 450630 494708 450636 494720
rect 450688 494708 450694 494760
rect 361758 491308 361764 491360
rect 361816 491348 361822 491360
rect 417510 491348 417516 491360
rect 361816 491320 417516 491348
rect 361816 491308 361822 491320
rect 417510 491308 417516 491320
rect 417568 491308 417574 491360
rect 397546 489880 397552 489932
rect 397604 489920 397610 489932
rect 397604 489892 398880 489920
rect 397604 489880 397610 489892
rect 398852 489852 398880 489892
rect 400950 489852 400956 489864
rect 398852 489824 400956 489852
rect 400950 489812 400956 489824
rect 401008 489812 401014 489864
rect 518158 484372 518164 484424
rect 518216 484412 518222 484424
rect 580166 484412 580172 484424
rect 518216 484384 580172 484412
rect 518216 484372 518222 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 361758 480224 361764 480276
rect 361816 480264 361822 480276
rect 364978 480264 364984 480276
rect 361816 480236 364984 480264
rect 361816 480224 361822 480236
rect 364978 480224 364984 480236
rect 365036 480224 365042 480276
rect 400950 476756 400956 476808
rect 401008 476796 401014 476808
rect 402238 476796 402244 476808
rect 401008 476768 402244 476796
rect 401008 476756 401014 476768
rect 402238 476756 402244 476768
rect 402296 476756 402302 476808
rect 518250 470568 518256 470620
rect 518308 470608 518314 470620
rect 579982 470608 579988 470620
rect 518308 470580 579988 470608
rect 518308 470568 518314 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 402238 469820 402244 469872
rect 402296 469860 402302 469872
rect 406010 469860 406016 469872
rect 402296 469832 406016 469860
rect 402296 469820 402302 469832
rect 406010 469820 406016 469832
rect 406068 469820 406074 469872
rect 361758 469208 361764 469260
rect 361816 469248 361822 469260
rect 418982 469248 418988 469260
rect 361816 469220 418988 469248
rect 361816 469208 361822 469220
rect 418982 469208 418988 469220
rect 419040 469208 419046 469260
rect 406010 465060 406016 465112
rect 406068 465100 406074 465112
rect 406068 465072 407160 465100
rect 406068 465060 406074 465072
rect 407132 465032 407160 465072
rect 409138 465032 409144 465044
rect 407132 465004 409144 465032
rect 409138 464992 409144 465004
rect 409196 464992 409202 465044
rect 514110 464380 514116 464432
rect 514168 464420 514174 464432
rect 542354 464420 542360 464432
rect 514168 464392 542360 464420
rect 514168 464380 514174 464392
rect 542354 464380 542360 464392
rect 542412 464380 542418 464432
rect 450078 464312 450084 464364
rect 450136 464352 450142 464364
rect 525794 464352 525800 464364
rect 450136 464324 525800 464352
rect 450136 464312 450142 464324
rect 525794 464312 525800 464324
rect 525852 464312 525858 464364
rect 494698 462476 494704 462528
rect 494756 462516 494762 462528
rect 527634 462516 527640 462528
rect 494756 462488 527640 462516
rect 494756 462476 494762 462488
rect 527634 462476 527640 462488
rect 527692 462476 527698 462528
rect 436094 462408 436100 462460
rect 436152 462448 436158 462460
rect 554130 462448 554136 462460
rect 436152 462420 554136 462448
rect 436152 462408 436158 462420
rect 554130 462408 554136 462420
rect 554188 462408 554194 462460
rect 433242 462340 433248 462392
rect 433300 462380 433306 462392
rect 551186 462380 551192 462392
rect 433300 462352 551192 462380
rect 433300 462340 433306 462352
rect 551186 462340 551192 462352
rect 551244 462340 551250 462392
rect 480162 461592 480168 461644
rect 480220 461632 480226 461644
rect 521746 461632 521752 461644
rect 480220 461604 521752 461632
rect 480220 461592 480226 461604
rect 521746 461592 521752 461604
rect 521804 461592 521810 461644
rect 450170 460912 450176 460964
rect 450228 460952 450234 460964
rect 524414 460952 524420 460964
rect 450228 460924 524420 460952
rect 450228 460912 450234 460924
rect 524414 460912 524420 460924
rect 524472 460912 524478 460964
rect 361758 458192 361764 458244
rect 361816 458232 361822 458244
rect 381630 458232 381636 458244
rect 361816 458204 381636 458232
rect 361816 458192 361822 458204
rect 381630 458192 381636 458204
rect 381688 458192 381694 458244
rect 409138 458124 409144 458176
rect 409196 458164 409202 458176
rect 409874 458164 409880 458176
rect 409196 458136 409880 458164
rect 409196 458124 409202 458136
rect 409874 458124 409880 458136
rect 409932 458124 409938 458176
rect 449802 457444 449808 457496
rect 449860 457484 449866 457496
rect 488534 457484 488540 457496
rect 449860 457456 488540 457484
rect 449860 457444 449866 457456
rect 488534 457444 488540 457456
rect 488592 457444 488598 457496
rect 473722 456764 473728 456816
rect 473780 456804 473786 456816
rect 480162 456804 480168 456816
rect 473780 456776 480168 456804
rect 473780 456764 473786 456776
rect 480162 456764 480168 456776
rect 480220 456764 480226 456816
rect 488258 456016 488264 456068
rect 488316 456056 488322 456068
rect 494698 456056 494704 456068
rect 488316 456028 494704 456056
rect 488316 456016 488322 456028
rect 494698 456016 494704 456028
rect 494756 456016 494762 456068
rect 450630 455472 450636 455524
rect 450688 455512 450694 455524
rect 480990 455512 480996 455524
rect 450688 455484 480996 455512
rect 450688 455472 450694 455484
rect 480990 455472 480996 455484
rect 481048 455472 481054 455524
rect 409874 455404 409880 455456
rect 409932 455444 409938 455456
rect 409932 455416 412634 455444
rect 409932 455404 409938 455416
rect 412606 455376 412634 455416
rect 423582 455404 423588 455456
rect 423640 455444 423646 455456
rect 473722 455444 473728 455456
rect 423640 455416 473728 455444
rect 423640 455404 423646 455416
rect 473722 455404 473728 455416
rect 473780 455404 473786 455456
rect 414382 455376 414388 455388
rect 412606 455348 414388 455376
rect 414382 455336 414388 455348
rect 414440 455336 414446 455388
rect 450262 454792 450268 454844
rect 450320 454832 450326 454844
rect 481726 454832 481732 454844
rect 450320 454804 481732 454832
rect 450320 454792 450326 454804
rect 481726 454792 481732 454804
rect 481784 454792 481790 454844
rect 449710 454724 449716 454776
rect 449768 454764 449774 454776
rect 484394 454764 484400 454776
rect 449768 454736 484400 454764
rect 449768 454724 449774 454736
rect 484394 454724 484400 454736
rect 484452 454724 484458 454776
rect 449618 454656 449624 454708
rect 449676 454696 449682 454708
rect 487154 454696 487160 454708
rect 449676 454668 487160 454696
rect 449676 454656 449682 454668
rect 487154 454656 487160 454668
rect 487212 454656 487218 454708
rect 414382 453296 414388 453348
rect 414440 453336 414446 453348
rect 416682 453336 416688 453348
rect 414440 453308 416688 453336
rect 414440 453296 414446 453308
rect 416682 453296 416688 453308
rect 416740 453296 416746 453348
rect 416682 447924 416688 447976
rect 416740 447964 416746 447976
rect 419074 447964 419080 447976
rect 416740 447936 419080 447964
rect 416740 447924 416746 447936
rect 419074 447924 419080 447936
rect 419132 447924 419138 447976
rect 422478 447516 422484 447568
rect 422536 447556 422542 447568
rect 423582 447556 423588 447568
rect 422536 447528 423588 447556
rect 422536 447516 422542 447528
rect 423582 447516 423588 447528
rect 423640 447516 423646 447568
rect 432414 447516 432420 447568
rect 432472 447556 432478 447568
rect 433242 447556 433248 447568
rect 432472 447528 433248 447556
rect 432472 447516 432478 447528
rect 433242 447516 433248 447528
rect 433300 447516 433306 447568
rect 361574 447176 361580 447228
rect 361632 447216 361638 447228
rect 363782 447216 363788 447228
rect 361632 447188 363788 447216
rect 361632 447176 361638 447188
rect 363782 447176 363788 447188
rect 363840 447176 363846 447228
rect 433242 447176 433248 447228
rect 433300 447216 433306 447228
rect 444190 447216 444196 447228
rect 433300 447188 444196 447216
rect 433300 447176 433306 447188
rect 444190 447176 444196 447188
rect 444248 447176 444254 447228
rect 423582 447108 423588 447160
rect 423640 447148 423646 447160
rect 445570 447148 445576 447160
rect 423640 447120 445576 447148
rect 423640 447108 423646 447120
rect 445570 447108 445576 447120
rect 445628 447108 445634 447160
rect 436094 445680 436100 445732
rect 436152 445720 436158 445732
rect 437382 445720 437388 445732
rect 436152 445692 437388 445720
rect 436152 445680 436158 445692
rect 437382 445680 437388 445692
rect 437440 445680 437446 445732
rect 427722 444524 427728 444576
rect 427780 444564 427786 444576
rect 446214 444564 446220 444576
rect 427780 444536 446220 444564
rect 427780 444524 427786 444536
rect 446214 444524 446220 444536
rect 446272 444524 446278 444576
rect 437290 444456 437296 444508
rect 437348 444496 437354 444508
rect 444374 444496 444380 444508
rect 437348 444468 444380 444496
rect 437348 444456 437354 444468
rect 444374 444456 444380 444468
rect 444432 444456 444438 444508
rect 442626 444388 442632 444440
rect 442684 444428 442690 444440
rect 444098 444428 444104 444440
rect 442684 444400 444104 444428
rect 442684 444388 442690 444400
rect 444098 444388 444104 444400
rect 444156 444388 444162 444440
rect 444190 444320 444196 444372
rect 444248 444360 444254 444372
rect 447226 444360 447232 444372
rect 444248 444332 447232 444360
rect 444248 444320 444254 444332
rect 447226 444320 447232 444332
rect 447284 444320 447290 444372
rect 456886 429836 456892 429888
rect 456944 429876 456950 429888
rect 474274 429876 474280 429888
rect 456944 429848 474280 429876
rect 456944 429836 456950 429848
rect 474274 429836 474280 429848
rect 474332 429836 474338 429888
rect 480898 429156 480904 429208
rect 480956 429196 480962 429208
rect 482278 429196 482284 429208
rect 480956 429168 482284 429196
rect 480956 429156 480962 429168
rect 482278 429156 482284 429168
rect 482336 429156 482342 429208
rect 483658 429156 483664 429208
rect 483716 429196 483722 429208
rect 484946 429196 484952 429208
rect 483716 429168 484952 429196
rect 483716 429156 483722 429168
rect 484946 429156 484952 429168
rect 485004 429156 485010 429208
rect 486418 429156 486424 429208
rect 486476 429196 486482 429208
rect 487614 429196 487620 429208
rect 486476 429168 487620 429196
rect 486476 429156 486482 429168
rect 487614 429156 487620 429168
rect 487672 429156 487678 429208
rect 457530 428408 457536 428460
rect 457588 428448 457594 428460
rect 471606 428448 471612 428460
rect 457588 428420 471612 428448
rect 457588 428408 457594 428420
rect 471606 428408 471612 428420
rect 471664 428408 471670 428460
rect 502518 424328 502524 424380
rect 502576 424368 502582 424380
rect 557534 424368 557540 424380
rect 502576 424340 557540 424368
rect 502576 424328 502582 424340
rect 557534 424328 557540 424340
rect 557592 424328 557598 424380
rect 529198 423580 529204 423632
rect 529256 423620 529262 423632
rect 530210 423620 530216 423632
rect 529256 423592 530216 423620
rect 529256 423580 529262 423592
rect 530210 423580 530216 423592
rect 530268 423580 530274 423632
rect 530578 423580 530584 423632
rect 530636 423620 530642 423632
rect 532786 423620 532792 423632
rect 530636 423592 532792 423620
rect 530636 423580 530642 423592
rect 532786 423580 532792 423592
rect 532844 423580 532850 423632
rect 511442 423512 511448 423564
rect 511500 423552 511506 423564
rect 523770 423552 523776 423564
rect 511500 423524 523776 423552
rect 511500 423512 511506 423524
rect 523770 423512 523776 423524
rect 523828 423512 523834 423564
rect 522298 423444 522304 423496
rect 522356 423484 522362 423496
rect 549530 423484 549536 423496
rect 522356 423456 549536 423484
rect 522356 423444 522362 423456
rect 549530 423444 549536 423456
rect 549588 423444 549594 423496
rect 502978 423376 502984 423428
rect 503036 423416 503042 423428
rect 522482 423416 522488 423428
rect 503036 423388 522488 423416
rect 503036 423376 503042 423388
rect 522482 423376 522488 423388
rect 522540 423376 522546 423428
rect 523678 423376 523684 423428
rect 523736 423416 523742 423428
rect 552106 423416 552112 423428
rect 523736 423388 552112 423416
rect 523736 423376 523742 423388
rect 552106 423376 552112 423388
rect 552164 423376 552170 423428
rect 485774 423308 485780 423360
rect 485832 423348 485838 423360
rect 526346 423348 526352 423360
rect 485832 423320 526352 423348
rect 485832 423308 485838 423320
rect 526346 423308 526352 423320
rect 526404 423308 526410 423360
rect 526438 423308 526444 423360
rect 526496 423348 526502 423360
rect 554682 423348 554688 423360
rect 526496 423320 554688 423348
rect 526496 423308 526502 423320
rect 554682 423308 554688 423320
rect 554740 423308 554746 423360
rect 487154 423240 487160 423292
rect 487212 423280 487218 423292
rect 528922 423280 528928 423292
rect 487212 423252 528928 423280
rect 487212 423240 487218 423252
rect 528922 423240 528928 423252
rect 528980 423240 528986 423292
rect 488534 423172 488540 423224
rect 488592 423212 488598 423224
rect 531498 423212 531504 423224
rect 488592 423184 531504 423212
rect 488592 423172 488598 423184
rect 531498 423172 531504 423184
rect 531556 423172 531562 423224
rect 496814 423104 496820 423156
rect 496872 423144 496878 423156
rect 545666 423144 545672 423156
rect 496872 423116 545672 423144
rect 496872 423104 496878 423116
rect 545666 423104 545672 423116
rect 545724 423104 545730 423156
rect 498194 423036 498200 423088
rect 498252 423076 498258 423088
rect 548242 423076 548248 423088
rect 498252 423048 548248 423076
rect 498252 423036 498258 423048
rect 548242 423036 548248 423048
rect 548300 423036 548306 423088
rect 499574 422968 499580 423020
rect 499632 423008 499638 423020
rect 550818 423008 550824 423020
rect 499632 422980 550824 423008
rect 499632 422968 499638 422980
rect 550818 422968 550824 422980
rect 550876 422968 550882 423020
rect 501046 422900 501052 422952
rect 501104 422940 501110 422952
rect 553394 422940 553400 422952
rect 501104 422912 553400 422940
rect 501104 422900 501110 422912
rect 553394 422900 553400 422912
rect 553452 422900 553458 422952
rect 483014 421540 483020 421592
rect 483072 421580 483078 421592
rect 521194 421580 521200 421592
rect 483072 421552 521200 421580
rect 483072 421540 483078 421552
rect 521194 421540 521200 421552
rect 521252 421540 521258 421592
rect 419074 420588 419080 420640
rect 419132 420628 419138 420640
rect 423950 420628 423956 420640
rect 419132 420600 423956 420628
rect 419132 420588 419138 420600
rect 423950 420588 423956 420600
rect 424008 420588 424014 420640
rect 494054 420180 494060 420232
rect 494112 420220 494118 420232
rect 541802 420220 541808 420232
rect 494112 420192 541808 420220
rect 494112 420180 494118 420192
rect 541802 420180 541808 420192
rect 541860 420180 541866 420232
rect 362310 418752 362316 418804
rect 362368 418792 362374 418804
rect 440878 418792 440884 418804
rect 362368 418764 440884 418792
rect 362368 418752 362374 418764
rect 440878 418752 440884 418764
rect 440936 418752 440942 418804
rect 421466 417732 421472 417784
rect 421524 417772 421530 417784
rect 503714 417772 503720 417784
rect 421524 417744 503720 417772
rect 421524 417732 421530 417744
rect 503714 417732 503720 417744
rect 503772 417732 503778 417784
rect 425330 417664 425336 417716
rect 425388 417704 425394 417716
rect 507854 417704 507860 417716
rect 425388 417676 507860 417704
rect 425388 417664 425394 417676
rect 507854 417664 507860 417676
rect 507912 417664 507918 417716
rect 424042 417596 424048 417648
rect 424100 417636 424106 417648
rect 506474 417636 506480 417648
rect 424100 417608 506480 417636
rect 424100 417596 424106 417608
rect 506474 417596 506480 417608
rect 506532 417596 506538 417648
rect 424686 417528 424692 417580
rect 424744 417568 424750 417580
rect 506566 417568 506572 417580
rect 424744 417540 506572 417568
rect 424744 417528 424750 417540
rect 506566 417528 506572 417540
rect 506624 417528 506630 417580
rect 422110 417460 422116 417512
rect 422168 417500 422174 417512
rect 503990 417500 503996 417512
rect 422168 417472 503996 417500
rect 422168 417460 422174 417472
rect 503990 417460 503996 417472
rect 504048 417460 504054 417512
rect 425974 417392 425980 417444
rect 426032 417432 426038 417444
rect 507946 417432 507952 417444
rect 426032 417404 507952 417432
rect 426032 417392 426038 417404
rect 507946 417392 507952 417404
rect 508004 417392 508010 417444
rect 423950 416780 423956 416832
rect 424008 416820 424014 416832
rect 428458 416820 428464 416832
rect 424008 416792 428464 416820
rect 424008 416780 424014 416792
rect 428458 416780 428464 416792
rect 428516 416780 428522 416832
rect 362218 416032 362224 416084
rect 362276 416072 362282 416084
rect 436738 416072 436744 416084
rect 362276 416044 436744 416072
rect 362276 416032 362282 416044
rect 436738 416032 436744 416044
rect 436796 416032 436802 416084
rect 361574 413992 361580 414044
rect 361632 414032 361638 414044
rect 439498 414032 439504 414044
rect 361632 414004 439504 414032
rect 361632 413992 361638 414004
rect 439498 413992 439504 414004
rect 439556 413992 439562 414044
rect 428458 411272 428464 411324
rect 428516 411312 428522 411324
rect 431218 411312 431224 411324
rect 428516 411284 431224 411312
rect 428516 411272 428522 411284
rect 431218 411272 431224 411284
rect 431276 411272 431282 411324
rect 511350 404336 511356 404388
rect 511408 404376 511414 404388
rect 580166 404376 580172 404388
rect 511408 404348 580172 404376
rect 511408 404336 511414 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 361574 402976 361580 403028
rect 361632 403016 361638 403028
rect 442258 403016 442264 403028
rect 361632 402988 442264 403016
rect 361632 402976 361638 402988
rect 442258 402976 442264 402988
rect 442316 402976 442322 403028
rect 497458 400868 497464 400920
rect 497516 400908 497522 400920
rect 546494 400908 546500 400920
rect 497516 400880 546500 400908
rect 497516 400868 497522 400880
rect 546494 400868 546500 400880
rect 546552 400868 546558 400920
rect 431218 400120 431224 400172
rect 431276 400160 431282 400172
rect 432598 400160 432604 400172
rect 431276 400132 432604 400160
rect 431276 400120 431282 400132
rect 432598 400120 432604 400132
rect 432656 400120 432662 400172
rect 494146 399440 494152 399492
rect 494204 399480 494210 399492
rect 539594 399480 539600 399492
rect 494204 399452 539600 399480
rect 494204 399440 494210 399452
rect 539594 399440 539600 399452
rect 539652 399440 539658 399492
rect 459922 398080 459928 398132
rect 459980 398120 459986 398132
rect 483658 398120 483664 398132
rect 459980 398092 483664 398120
rect 459980 398080 459986 398092
rect 483658 398080 483664 398092
rect 483716 398080 483722 398132
rect 492674 398080 492680 398132
rect 492732 398120 492738 398132
rect 538214 398120 538220 398132
rect 492732 398092 538220 398120
rect 492732 398080 492738 398092
rect 538214 398080 538220 398092
rect 538272 398080 538278 398132
rect 458450 396720 458456 396772
rect 458508 396760 458514 396772
rect 478874 396760 478880 396772
rect 458508 396732 478880 396760
rect 458508 396720 458514 396732
rect 478874 396720 478880 396732
rect 478932 396720 478938 396772
rect 492766 396720 492772 396772
rect 492824 396760 492830 396772
rect 536834 396760 536840 396772
rect 492824 396732 536840 396760
rect 492824 396720 492830 396732
rect 536834 396720 536840 396732
rect 536892 396720 536898 396772
rect 458174 395292 458180 395344
rect 458232 395332 458238 395344
rect 476114 395332 476120 395344
rect 458232 395304 476120 395332
rect 458232 395292 458238 395304
rect 476114 395292 476120 395304
rect 476172 395292 476178 395344
rect 491570 395292 491576 395344
rect 491628 395332 491634 395344
rect 535454 395332 535460 395344
rect 491628 395304 535460 395332
rect 491628 395292 491634 395304
rect 535454 395292 535460 395304
rect 535512 395292 535518 395344
rect 465534 393932 465540 393984
rect 465592 393972 465598 393984
rect 490006 393972 490012 393984
rect 465592 393944 490012 393972
rect 465592 393932 465598 393944
rect 490006 393932 490012 393944
rect 490064 393932 490070 393984
rect 491294 393932 491300 393984
rect 491352 393972 491358 393984
rect 534166 393972 534172 393984
rect 491352 393944 534172 393972
rect 491352 393932 491358 393944
rect 534166 393932 534172 393944
rect 534224 393932 534230 393984
rect 496446 392640 496452 392692
rect 496504 392680 496510 392692
rect 543734 392680 543740 392692
rect 496504 392652 543740 392680
rect 496504 392640 496510 392652
rect 543734 392640 543740 392652
rect 543792 392640 543798 392692
rect 422386 392572 422392 392624
rect 422444 392612 422450 392624
rect 506014 392612 506020 392624
rect 422444 392584 506020 392612
rect 422444 392572 422450 392584
rect 506014 392572 506020 392584
rect 506072 392572 506078 392624
rect 361574 391960 361580 392012
rect 361632 392000 361638 392012
rect 440970 392000 440976 392012
rect 361632 391972 440976 392000
rect 361632 391960 361638 391972
rect 440970 391960 440976 391972
rect 441028 391960 441034 392012
rect 459646 391280 459652 391332
rect 459704 391320 459710 391332
rect 480898 391320 480904 391332
rect 459704 391292 480904 391320
rect 459704 391280 459710 391292
rect 480898 391280 480904 391292
rect 480956 391280 480962 391332
rect 495710 391280 495716 391332
rect 495768 391320 495774 391332
rect 542354 391320 542360 391332
rect 495768 391292 542360 391320
rect 495768 391280 495774 391292
rect 542354 391280 542360 391292
rect 542412 391280 542418 391332
rect 422294 391212 422300 391264
rect 422352 391252 422358 391264
rect 505278 391252 505284 391264
rect 422352 391224 505284 391252
rect 422352 391212 422358 391224
rect 505278 391212 505284 391224
rect 505336 391212 505342 391264
rect 461118 389784 461124 389836
rect 461176 389824 461182 389836
rect 486418 389824 486424 389836
rect 461176 389796 486424 389824
rect 461176 389784 461182 389796
rect 486418 389784 486424 389796
rect 486476 389784 486482 389836
rect 490558 389784 490564 389836
rect 490616 389824 490622 389836
rect 534074 389824 534080 389836
rect 490616 389796 534080 389824
rect 490616 389784 490622 389796
rect 534074 389784 534080 389796
rect 534132 389784 534138 389836
rect 449894 389240 449900 389292
rect 449952 389280 449958 389292
rect 450722 389280 450728 389292
rect 449952 389252 450728 389280
rect 449952 389240 449958 389252
rect 450722 389240 450728 389252
rect 450780 389240 450786 389292
rect 465074 389240 465080 389292
rect 465132 389280 465138 389292
rect 465902 389280 465908 389292
rect 465132 389252 465908 389280
rect 465132 389240 465138 389252
rect 465902 389240 465908 389252
rect 465960 389240 465966 389292
rect 492674 389240 492680 389292
rect 492732 389280 492738 389292
rect 493134 389280 493140 389292
rect 492732 389252 493140 389280
rect 492732 389240 492738 389252
rect 493134 389240 493140 389252
rect 493192 389240 493198 389292
rect 494054 389240 494060 389292
rect 494112 389280 494118 389292
rect 494606 389280 494612 389292
rect 494112 389252 494612 389280
rect 494112 389240 494118 389252
rect 494606 389240 494612 389252
rect 494664 389240 494670 389292
rect 453758 389104 453764 389156
rect 453816 389144 453822 389156
rect 454678 389144 454684 389156
rect 453816 389116 454684 389144
rect 453816 389104 453822 389116
rect 454678 389104 454684 389116
rect 454736 389104 454742 389156
rect 461670 389104 461676 389156
rect 461728 389144 461734 389156
rect 462590 389144 462596 389156
rect 461728 389116 462596 389144
rect 461728 389104 461734 389116
rect 462590 389104 462596 389116
rect 462648 389104 462654 389156
rect 464338 389104 464344 389156
rect 464396 389144 464402 389156
rect 469214 389144 469220 389156
rect 464396 389116 469220 389144
rect 464396 389104 464402 389116
rect 469214 389104 469220 389116
rect 469272 389104 469278 389156
rect 461854 389036 461860 389088
rect 461912 389076 461918 389088
rect 465534 389076 465540 389088
rect 461912 389048 465540 389076
rect 461912 389036 461918 389048
rect 465534 389036 465540 389048
rect 465592 389036 465598 389088
rect 483934 388968 483940 389020
rect 483992 389008 483998 389020
rect 502978 389008 502984 389020
rect 483992 388980 502984 389008
rect 483992 388968 483998 388980
rect 502978 388968 502984 388980
rect 503036 388968 503042 389020
rect 468478 388900 468484 388952
rect 468536 388940 468542 388952
rect 475102 388940 475108 388952
rect 468536 388912 475108 388940
rect 468536 388900 468542 388912
rect 475102 388900 475108 388912
rect 475160 388900 475166 388952
rect 499390 388900 499396 388952
rect 499448 388940 499454 388952
rect 522298 388940 522304 388952
rect 499448 388912 522304 388940
rect 499448 388900 499454 388912
rect 522298 388900 522304 388912
rect 522356 388900 522362 388952
rect 456702 388832 456708 388884
rect 456760 388872 456766 388884
rect 457530 388872 457536 388884
rect 456760 388844 457536 388872
rect 456760 388832 456766 388844
rect 457530 388832 457536 388844
rect 457588 388832 457594 388884
rect 468662 388832 468668 388884
rect 468720 388872 468726 388884
rect 480990 388872 480996 388884
rect 468720 388844 480996 388872
rect 468720 388832 468726 388844
rect 480990 388832 480996 388844
rect 481048 388832 481054 388884
rect 500862 388832 500868 388884
rect 500920 388872 500926 388884
rect 523678 388872 523684 388884
rect 500920 388844 523684 388872
rect 500920 388832 500926 388844
rect 523678 388832 523684 388844
rect 523736 388832 523742 388884
rect 468570 388764 468576 388816
rect 468628 388804 468634 388816
rect 478046 388804 478052 388816
rect 468628 388776 478052 388804
rect 468628 388764 468634 388776
rect 478046 388764 478052 388776
rect 478104 388764 478110 388816
rect 502334 388764 502340 388816
rect 502392 388804 502398 388816
rect 526438 388804 526444 388816
rect 502392 388776 526444 388804
rect 502392 388764 502398 388776
rect 526438 388764 526444 388776
rect 526496 388764 526502 388816
rect 467098 388696 467104 388748
rect 467156 388736 467162 388748
rect 480254 388736 480260 388748
rect 467156 388708 480260 388736
rect 467156 388696 467162 388708
rect 480254 388696 480260 388708
rect 480312 388696 480318 388748
rect 484670 388696 484676 388748
rect 484728 388736 484734 388748
rect 511442 388736 511448 388748
rect 484728 388708 511448 388736
rect 484728 388696 484734 388708
rect 511442 388696 511448 388708
rect 511500 388696 511506 388748
rect 467190 388628 467196 388680
rect 467248 388668 467254 388680
rect 481726 388668 481732 388680
rect 467248 388640 481732 388668
rect 467248 388628 467254 388640
rect 481726 388628 481732 388640
rect 481784 388628 481790 388680
rect 485406 388628 485412 388680
rect 485464 388668 485470 388680
rect 524414 388668 524420 388680
rect 485464 388640 524420 388668
rect 485464 388628 485470 388640
rect 524414 388628 524420 388640
rect 524472 388628 524478 388680
rect 461578 388560 461584 388612
rect 461636 388600 461642 388612
rect 476574 388600 476580 388612
rect 461636 388572 476580 388600
rect 461636 388560 461642 388572
rect 476574 388560 476580 388572
rect 476632 388560 476638 388612
rect 486878 388560 486884 388612
rect 486936 388600 486942 388612
rect 527174 388600 527180 388612
rect 486936 388572 527180 388600
rect 486936 388560 486942 388572
rect 527174 388560 527180 388572
rect 527232 388560 527238 388612
rect 461762 388492 461768 388544
rect 461820 388532 461826 388544
rect 478782 388532 478788 388544
rect 461820 388504 478788 388532
rect 461820 388492 461826 388504
rect 478782 388492 478788 388504
rect 478840 388492 478846 388544
rect 488350 388492 488356 388544
rect 488408 388532 488414 388544
rect 529198 388532 529204 388544
rect 488408 388504 529204 388532
rect 488408 388492 488414 388504
rect 529198 388492 529204 388504
rect 529256 388492 529262 388544
rect 462958 388424 462964 388476
rect 463016 388464 463022 388476
rect 482462 388464 482468 388476
rect 463016 388436 482468 388464
rect 463016 388424 463022 388436
rect 482462 388424 482468 388436
rect 482520 388424 482526 388476
rect 489822 388424 489828 388476
rect 489880 388464 489886 388476
rect 530578 388464 530584 388476
rect 489880 388436 530584 388464
rect 489880 388424 489886 388436
rect 530578 388424 530584 388436
rect 530636 388424 530642 388476
rect 447870 387132 447876 387184
rect 447928 387172 447934 387184
rect 457438 387172 457444 387184
rect 447928 387144 457444 387172
rect 447928 387132 447934 387144
rect 457438 387132 457444 387144
rect 457496 387132 457502 387184
rect 448974 387064 448980 387116
rect 449032 387104 449038 387116
rect 491110 387104 491116 387116
rect 449032 387076 491116 387104
rect 449032 387064 449038 387076
rect 491110 387064 491116 387076
rect 491168 387064 491174 387116
rect 445570 386520 445576 386572
rect 445628 386560 445634 386572
rect 553946 386560 553952 386572
rect 445628 386532 553952 386560
rect 445628 386520 445634 386532
rect 553946 386520 553952 386532
rect 554004 386520 554010 386572
rect 381538 386452 381544 386504
rect 381596 386492 381602 386504
rect 512178 386492 512184 386504
rect 381596 386464 512184 386492
rect 381596 386452 381602 386464
rect 512178 386452 512184 386464
rect 512236 386452 512242 386504
rect 370498 386384 370504 386436
rect 370556 386424 370562 386436
rect 511994 386424 512000 386436
rect 370556 386396 512000 386424
rect 370556 386384 370562 386396
rect 511994 386384 512000 386396
rect 512052 386384 512058 386436
rect 448422 385976 448428 386028
rect 448480 386016 448486 386028
rect 451918 386016 451924 386028
rect 448480 385988 451924 386016
rect 448480 385976 448486 385988
rect 451918 385976 451924 385988
rect 451976 385976 451982 386028
rect 447778 385364 447784 385416
rect 447836 385404 447842 385416
rect 453298 385404 453304 385416
rect 447836 385376 453304 385404
rect 447836 385364 447842 385376
rect 453298 385364 453304 385376
rect 453356 385364 453362 385416
rect 450354 385092 450360 385144
rect 450412 385132 450418 385144
rect 563422 385132 563428 385144
rect 450412 385104 563428 385132
rect 450412 385092 450418 385104
rect 563422 385092 563428 385104
rect 563480 385092 563486 385144
rect 370590 385024 370596 385076
rect 370648 385064 370654 385076
rect 512086 385064 512092 385076
rect 370648 385036 512092 385064
rect 370648 385024 370654 385036
rect 512086 385024 512092 385036
rect 512144 385024 512150 385076
rect 512730 383732 512736 383784
rect 512788 383772 512794 383784
rect 534718 383772 534724 383784
rect 512788 383744 534724 383772
rect 512788 383732 512794 383744
rect 534718 383732 534724 383744
rect 534776 383732 534782 383784
rect 513282 383664 513288 383716
rect 513340 383704 513346 383716
rect 547138 383704 547144 383716
rect 513340 383676 547144 383704
rect 513340 383664 513346 383676
rect 547138 383664 547144 383676
rect 547196 383664 547202 383716
rect 378778 383596 378784 383648
rect 378836 383636 378842 383648
rect 447318 383636 447324 383648
rect 378836 383608 447324 383636
rect 378836 383596 378842 383608
rect 447318 383596 447324 383608
rect 447376 383596 447382 383648
rect 382918 383528 382924 383580
rect 382976 383568 382982 383580
rect 447134 383568 447140 383580
rect 382976 383540 447140 383568
rect 382976 383528 382982 383540
rect 447134 383528 447140 383540
rect 447192 383528 447198 383580
rect 512454 382984 512460 383036
rect 512512 383024 512518 383036
rect 518342 383024 518348 383036
rect 512512 382996 518348 383024
rect 512512 382984 512518 382996
rect 518342 382984 518348 382996
rect 518400 382984 518406 383036
rect 513006 382440 513012 382492
rect 513064 382480 513070 382492
rect 519630 382480 519636 382492
rect 513064 382452 519636 382480
rect 513064 382440 513070 382452
rect 519630 382440 519636 382452
rect 519688 382440 519694 382492
rect 512270 382304 512276 382356
rect 512328 382344 512334 382356
rect 515582 382344 515588 382356
rect 512328 382316 515588 382344
rect 512328 382304 512334 382316
rect 515582 382304 515588 382316
rect 515640 382304 515646 382356
rect 376018 382168 376024 382220
rect 376076 382208 376082 382220
rect 447318 382208 447324 382220
rect 376076 382180 447324 382208
rect 376076 382168 376082 382180
rect 447318 382168 447324 382180
rect 447376 382168 447382 382220
rect 400858 382100 400864 382152
rect 400916 382140 400922 382152
rect 447134 382140 447140 382152
rect 400916 382112 447140 382140
rect 400916 382100 400922 382112
rect 447134 382100 447140 382112
rect 447192 382100 447198 382152
rect 361574 380876 361580 380928
rect 361632 380916 361638 380928
rect 442350 380916 442356 380928
rect 361632 380888 442356 380916
rect 361632 380876 361638 380888
rect 442350 380876 442356 380888
rect 442408 380876 442414 380928
rect 513282 380876 513288 380928
rect 513340 380916 513346 380928
rect 548518 380916 548524 380928
rect 513340 380888 548524 380916
rect 513340 380876 513346 380888
rect 548518 380876 548524 380888
rect 548576 380876 548582 380928
rect 374638 380808 374644 380860
rect 374696 380848 374702 380860
rect 447502 380848 447508 380860
rect 374696 380820 447508 380848
rect 374696 380808 374702 380820
rect 447502 380808 447508 380820
rect 447560 380808 447566 380860
rect 403618 380740 403624 380792
rect 403676 380780 403682 380792
rect 447134 380780 447140 380792
rect 403676 380752 447140 380780
rect 403676 380740 403682 380752
rect 447134 380740 447140 380752
rect 447192 380740 447198 380792
rect 406378 380672 406384 380724
rect 406436 380712 406442 380724
rect 447318 380712 447324 380724
rect 406436 380684 447324 380712
rect 406436 380672 406442 380684
rect 447318 380672 447324 380684
rect 447376 380672 447382 380724
rect 511994 380400 512000 380452
rect 512052 380440 512058 380452
rect 512362 380440 512368 380452
rect 512052 380412 512368 380440
rect 512052 380400 512058 380412
rect 512362 380400 512368 380412
rect 512420 380400 512426 380452
rect 511994 380264 512000 380316
rect 512052 380304 512058 380316
rect 514202 380304 514208 380316
rect 512052 380276 514208 380304
rect 512052 380264 512058 380276
rect 514202 380264 514208 380276
rect 514260 380264 514266 380316
rect 513282 379516 513288 379568
rect 513340 379556 513346 379568
rect 544378 379556 544384 379568
rect 513340 379528 544384 379556
rect 513340 379516 513346 379528
rect 544378 379516 544384 379528
rect 544436 379516 544442 379568
rect 370682 379448 370688 379500
rect 370740 379488 370746 379500
rect 447502 379488 447508 379500
rect 370740 379460 447508 379488
rect 370740 379448 370746 379460
rect 447502 379448 447508 379460
rect 447560 379448 447566 379500
rect 371878 379380 371884 379432
rect 371936 379420 371942 379432
rect 447134 379420 447140 379432
rect 371936 379392 447140 379420
rect 371936 379380 371942 379392
rect 447134 379380 447140 379392
rect 447192 379380 447198 379432
rect 512178 378292 512184 378344
rect 512236 378332 512242 378344
rect 522298 378332 522304 378344
rect 512236 378304 522304 378332
rect 512236 378292 512242 378304
rect 522298 378292 522304 378304
rect 522356 378292 522362 378344
rect 513282 378224 513288 378276
rect 513340 378264 513346 378276
rect 548610 378264 548616 378276
rect 513340 378236 548616 378264
rect 513340 378224 513346 378236
rect 548610 378224 548616 378236
rect 548668 378224 548674 378276
rect 516778 378156 516784 378208
rect 516836 378196 516842 378208
rect 580166 378196 580172 378208
rect 516836 378168 580172 378196
rect 516836 378156 516842 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 363598 378088 363604 378140
rect 363656 378128 363662 378140
rect 447318 378128 447324 378140
rect 363656 378100 447324 378128
rect 363656 378088 363662 378100
rect 447318 378088 447324 378100
rect 447376 378088 447382 378140
rect 367738 378020 367744 378072
rect 367796 378060 367802 378072
rect 447134 378060 447140 378072
rect 367796 378032 447140 378060
rect 367796 378020 367802 378032
rect 447134 378020 447140 378032
rect 447192 378020 447198 378072
rect 432598 377952 432604 378004
rect 432656 377992 432662 378004
rect 436830 377992 436836 378004
rect 432656 377964 436836 377992
rect 432656 377952 432662 377964
rect 436830 377952 436836 377964
rect 436888 377952 436894 378004
rect 512822 377408 512828 377460
rect 512880 377448 512886 377460
rect 549898 377448 549904 377460
rect 512880 377420 549904 377448
rect 512880 377408 512886 377420
rect 549898 377408 549904 377420
rect 549956 377408 549962 377460
rect 513190 376728 513196 376780
rect 513248 376768 513254 376780
rect 516962 376768 516968 376780
rect 513248 376740 516968 376768
rect 513248 376728 513254 376740
rect 516962 376728 516968 376740
rect 517020 376728 517026 376780
rect 363690 376660 363696 376712
rect 363748 376700 363754 376712
rect 447134 376700 447140 376712
rect 363748 376672 447140 376700
rect 363748 376660 363754 376672
rect 447134 376660 447140 376672
rect 447192 376660 447198 376712
rect 407758 376592 407764 376644
rect 407816 376632 407822 376644
rect 447318 376632 447324 376644
rect 407816 376604 447324 376632
rect 407816 376592 407822 376604
rect 447318 376592 447324 376604
rect 447376 376592 447382 376644
rect 512454 375980 512460 376032
rect 512512 376020 512518 376032
rect 547230 376020 547236 376032
rect 512512 375992 547236 376020
rect 512512 375980 512518 375992
rect 547230 375980 547236 375992
rect 547288 375980 547294 376032
rect 513282 375640 513288 375692
rect 513340 375680 513346 375692
rect 520274 375680 520280 375692
rect 513340 375652 520280 375680
rect 513340 375640 513346 375652
rect 520274 375640 520280 375652
rect 520332 375640 520338 375692
rect 410518 375300 410524 375352
rect 410576 375340 410582 375352
rect 447134 375340 447140 375352
rect 410576 375312 447140 375340
rect 410576 375300 410582 375312
rect 447134 375300 447140 375312
rect 447192 375300 447198 375352
rect 411898 375232 411904 375284
rect 411956 375272 411962 375284
rect 447318 375272 447324 375284
rect 411956 375244 447324 375272
rect 411956 375232 411962 375244
rect 447318 375232 447324 375244
rect 447376 375232 447382 375284
rect 512454 374144 512460 374196
rect 512512 374184 512518 374196
rect 515674 374184 515680 374196
rect 512512 374156 515680 374184
rect 512512 374144 512518 374156
rect 515674 374144 515680 374156
rect 515732 374144 515738 374196
rect 414658 373940 414664 373992
rect 414716 373980 414722 373992
rect 447134 373980 447140 373992
rect 414716 373952 447140 373980
rect 414716 373940 414722 373952
rect 447134 373940 447140 373952
rect 447192 373940 447198 373992
rect 416038 373872 416044 373924
rect 416096 373912 416102 373924
rect 447318 373912 447324 373924
rect 416096 373884 447324 373912
rect 416096 373872 416102 373884
rect 447318 373872 447324 373884
rect 447376 373872 447382 373924
rect 512638 373736 512644 373788
rect 512696 373776 512702 373788
rect 516226 373776 516232 373788
rect 512696 373748 516232 373776
rect 512696 373736 512702 373748
rect 516226 373736 516232 373748
rect 516284 373736 516290 373788
rect 513282 372716 513288 372768
rect 513340 372756 513346 372768
rect 521654 372756 521660 372768
rect 513340 372728 521660 372756
rect 513340 372716 513346 372728
rect 521654 372716 521660 372728
rect 521712 372716 521718 372768
rect 512086 372648 512092 372700
rect 512144 372688 512150 372700
rect 514846 372688 514852 372700
rect 512144 372660 514852 372688
rect 512144 372648 512150 372660
rect 514846 372648 514852 372660
rect 514904 372648 514910 372700
rect 364978 372512 364984 372564
rect 365036 372552 365042 372564
rect 447318 372552 447324 372564
rect 365036 372524 447324 372552
rect 365036 372512 365042 372524
rect 447318 372512 447324 372524
rect 447376 372512 447382 372564
rect 417510 372444 417516 372496
rect 417568 372484 417574 372496
rect 447134 372484 447140 372496
rect 417568 372456 447140 372484
rect 417568 372444 417574 372456
rect 447134 372444 447140 372456
rect 447192 372444 447198 372496
rect 512454 371764 512460 371816
rect 512512 371804 512518 371816
rect 516318 371804 516324 371816
rect 512512 371776 516324 371804
rect 512512 371764 512518 371776
rect 516318 371764 516324 371776
rect 516376 371764 516382 371816
rect 381630 371152 381636 371204
rect 381688 371192 381694 371204
rect 447318 371192 447324 371204
rect 381688 371164 447324 371192
rect 381688 371152 381694 371164
rect 447318 371152 447324 371164
rect 447376 371152 447382 371204
rect 418982 371084 418988 371136
rect 419040 371124 419046 371136
rect 447134 371124 447140 371136
rect 419040 371096 447140 371124
rect 419040 371084 419046 371096
rect 447134 371084 447140 371096
rect 447192 371084 447198 371136
rect 513282 370064 513288 370116
rect 513340 370104 513346 370116
rect 520366 370104 520372 370116
rect 513340 370076 520372 370104
rect 513340 370064 513346 370076
rect 520366 370064 520372 370076
rect 520424 370064 520430 370116
rect 512730 369928 512736 369980
rect 512788 369968 512794 369980
rect 516134 369968 516140 369980
rect 512788 369940 516140 369968
rect 512788 369928 512794 369940
rect 516134 369928 516140 369940
rect 516192 369928 516198 369980
rect 361574 369860 361580 369912
rect 361632 369900 361638 369912
rect 429194 369900 429200 369912
rect 361632 369872 429200 369900
rect 361632 369860 361638 369872
rect 429194 369860 429200 369872
rect 429252 369860 429258 369912
rect 363782 369792 363788 369844
rect 363840 369832 363846 369844
rect 447134 369832 447140 369844
rect 363840 369804 447140 369832
rect 363840 369792 363846 369804
rect 447134 369792 447140 369804
rect 447192 369792 447198 369844
rect 436738 369724 436744 369776
rect 436796 369764 436802 369776
rect 447318 369764 447324 369776
rect 436796 369736 447324 369764
rect 436796 369724 436802 369736
rect 447318 369724 447324 369736
rect 447376 369724 447382 369776
rect 513282 368500 513288 368552
rect 513340 368540 513346 368552
rect 520458 368540 520464 368552
rect 513340 368512 520464 368540
rect 513340 368500 513346 368512
rect 520458 368500 520464 368512
rect 520516 368500 520522 368552
rect 439498 368432 439504 368484
rect 439556 368472 439562 368484
rect 447318 368472 447324 368484
rect 439556 368444 447324 368472
rect 439556 368432 439562 368444
rect 447318 368432 447324 368444
rect 447376 368432 447382 368484
rect 440878 368364 440884 368416
rect 440936 368404 440942 368416
rect 447134 368404 447140 368416
rect 440936 368376 447140 368404
rect 440936 368364 440942 368376
rect 447134 368364 447140 368376
rect 447192 368364 447198 368416
rect 512638 367344 512644 367396
rect 512696 367384 512702 367396
rect 518986 367384 518992 367396
rect 512696 367356 518992 367384
rect 512696 367344 512702 367356
rect 518986 367344 518992 367356
rect 519044 367344 519050 367396
rect 511994 367208 512000 367260
rect 512052 367248 512058 367260
rect 514938 367248 514944 367260
rect 512052 367220 514944 367248
rect 512052 367208 512058 367220
rect 514938 367208 514944 367220
rect 514996 367208 515002 367260
rect 440970 367004 440976 367056
rect 441028 367044 441034 367056
rect 447134 367044 447140 367056
rect 441028 367016 447140 367044
rect 441028 367004 441034 367016
rect 447134 367004 447140 367016
rect 447192 367004 447198 367056
rect 442258 366936 442264 366988
rect 442316 366976 442322 366988
rect 447318 366976 447324 366988
rect 442316 366948 447324 366976
rect 442316 366936 442322 366948
rect 447318 366936 447324 366948
rect 447376 366936 447382 366988
rect 513282 365848 513288 365900
rect 513340 365888 513346 365900
rect 520550 365888 520556 365900
rect 513340 365860 520556 365888
rect 513340 365848 513346 365860
rect 520550 365848 520556 365860
rect 520608 365848 520614 365900
rect 513190 365712 513196 365764
rect 513248 365752 513254 365764
rect 518894 365752 518900 365764
rect 513248 365724 518900 365752
rect 513248 365712 513254 365724
rect 518894 365712 518900 365724
rect 518952 365712 518958 365764
rect 429194 365644 429200 365696
rect 429252 365684 429258 365696
rect 447134 365684 447140 365696
rect 429252 365656 447140 365684
rect 429252 365644 429258 365656
rect 447134 365644 447140 365656
rect 447192 365644 447198 365696
rect 442350 365576 442356 365628
rect 442408 365616 442414 365628
rect 447318 365616 447324 365628
rect 442408 365588 447324 365616
rect 442408 365576 442414 365588
rect 447318 365576 447324 365588
rect 447376 365576 447382 365628
rect 511994 364488 512000 364540
rect 512052 364528 512058 364540
rect 514294 364528 514300 364540
rect 512052 364500 514300 364528
rect 512052 364488 512058 364500
rect 514294 364488 514300 364500
rect 514352 364488 514358 364540
rect 513282 364352 513288 364404
rect 513340 364392 513346 364404
rect 523034 364392 523040 364404
rect 513340 364364 523040 364392
rect 513340 364352 513346 364364
rect 523034 364352 523040 364364
rect 523092 364352 523098 364404
rect 569218 364352 569224 364404
rect 569276 364392 569282 364404
rect 580166 364392 580172 364404
rect 569276 364364 580172 364392
rect 569276 364352 569282 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 512086 363536 512092 363588
rect 512144 363576 512150 363588
rect 513650 363576 513656 363588
rect 512144 363548 513656 363576
rect 512144 363536 512150 363548
rect 513650 363536 513656 363548
rect 513708 363536 513714 363588
rect 437014 362992 437020 363044
rect 437072 363032 437078 363044
rect 447134 363032 447140 363044
rect 437072 363004 447140 363032
rect 437072 362992 437078 363004
rect 447134 362992 447140 363004
rect 447192 362992 447198 363044
rect 432598 362924 432604 362976
rect 432656 362964 432662 362976
rect 447318 362964 447324 362976
rect 432656 362936 447324 362964
rect 432656 362924 432662 362936
rect 447318 362924 447324 362936
rect 447376 362924 447382 362976
rect 512362 362312 512368 362364
rect 512420 362352 512426 362364
rect 513742 362352 513748 362364
rect 512420 362324 513748 362352
rect 512420 362312 512426 362324
rect 513742 362312 513748 362324
rect 513800 362312 513806 362364
rect 513190 361768 513196 361820
rect 513248 361808 513254 361820
rect 519078 361808 519084 361820
rect 513248 361780 519084 361808
rect 513248 361768 513254 361780
rect 519078 361768 519084 361780
rect 519136 361768 519142 361820
rect 442258 361632 442264 361684
rect 442316 361672 442322 361684
rect 447318 361672 447324 361684
rect 442316 361644 447324 361672
rect 442316 361632 442322 361644
rect 447318 361632 447324 361644
rect 447376 361632 447382 361684
rect 439682 361564 439688 361616
rect 439740 361604 439746 361616
rect 447134 361604 447140 361616
rect 439740 361576 447140 361604
rect 439740 361564 439746 361576
rect 447134 361564 447140 361576
rect 447192 361564 447198 361616
rect 513282 361564 513288 361616
rect 513340 361604 513346 361616
rect 521746 361604 521752 361616
rect 513340 361576 521752 361604
rect 513340 361564 513346 361576
rect 521746 361564 521752 361576
rect 521804 361564 521810 361616
rect 522298 360816 522304 360868
rect 522356 360856 522362 360868
rect 550634 360856 550640 360868
rect 522356 360828 550640 360856
rect 522356 360816 522362 360828
rect 550634 360816 550640 360828
rect 550692 360816 550698 360868
rect 512822 360408 512828 360460
rect 512880 360448 512886 360460
rect 519170 360448 519176 360460
rect 512880 360420 519176 360448
rect 512880 360408 512886 360420
rect 519170 360408 519176 360420
rect 519228 360408 519234 360460
rect 513282 360340 513288 360392
rect 513340 360380 513346 360392
rect 523126 360380 523132 360392
rect 513340 360352 523132 360380
rect 513340 360340 513346 360352
rect 523126 360340 523132 360352
rect 523184 360340 523190 360392
rect 442350 360272 442356 360324
rect 442408 360312 442414 360324
rect 447318 360312 447324 360324
rect 442408 360284 447324 360312
rect 442408 360272 442414 360284
rect 447318 360272 447324 360284
rect 447376 360272 447382 360324
rect 512362 360272 512368 360324
rect 512420 360312 512426 360324
rect 515122 360312 515128 360324
rect 512420 360284 515128 360312
rect 512420 360272 512426 360284
rect 515122 360272 515128 360284
rect 515180 360272 515186 360324
rect 435450 360204 435456 360256
rect 435508 360244 435514 360256
rect 447134 360244 447140 360256
rect 435508 360216 447140 360244
rect 435508 360204 435514 360216
rect 447134 360204 447140 360216
rect 447192 360204 447198 360256
rect 548610 360136 548616 360188
rect 548668 360176 548674 360188
rect 552014 360176 552020 360188
rect 548668 360148 552020 360176
rect 548668 360136 548674 360148
rect 552014 360136 552020 360148
rect 552072 360136 552078 360188
rect 548518 359048 548524 359100
rect 548576 359088 548582 359100
rect 558178 359088 558184 359100
rect 548576 359060 558184 359088
rect 548576 359048 548582 359060
rect 558178 359048 558184 359060
rect 558236 359048 558242 359100
rect 544378 358980 544384 359032
rect 544436 359020 544442 359032
rect 553762 359020 553768 359032
rect 544436 358992 553768 359020
rect 544436 358980 544442 358992
rect 553762 358980 553768 358992
rect 553820 358980 553826 359032
rect 512362 358912 512368 358964
rect 512420 358952 512426 358964
rect 513834 358952 513840 358964
rect 512420 358924 513840 358952
rect 512420 358912 512426 358924
rect 513834 358912 513840 358924
rect 513892 358912 513898 358964
rect 547138 358912 547144 358964
rect 547196 358952 547202 358964
rect 565538 358952 565544 358964
rect 547196 358924 565544 358952
rect 547196 358912 547202 358924
rect 565538 358912 565544 358924
rect 565596 358912 565602 358964
rect 441062 358844 441068 358896
rect 441120 358884 441126 358896
rect 447318 358884 447324 358896
rect 441120 358856 447324 358884
rect 441120 358844 441126 358856
rect 447318 358844 447324 358856
rect 447376 358844 447382 358896
rect 512914 358844 512920 358896
rect 512972 358884 512978 358896
rect 519262 358884 519268 358896
rect 512972 358856 519268 358884
rect 512972 358844 512978 358856
rect 519262 358844 519268 358856
rect 519320 358844 519326 358896
rect 534718 358844 534724 358896
rect 534776 358884 534782 358896
rect 567010 358884 567016 358896
rect 534776 358856 567016 358884
rect 534776 358844 534782 358856
rect 567010 358844 567016 358856
rect 567068 358844 567074 358896
rect 436922 358776 436928 358828
rect 436980 358816 436986 358828
rect 447134 358816 447140 358828
rect 436980 358788 447140 358816
rect 436980 358776 436986 358788
rect 447134 358776 447140 358788
rect 447192 358776 447198 358828
rect 514202 358776 514208 358828
rect 514260 358816 514266 358828
rect 555234 358816 555240 358828
rect 514260 358788 555240 358816
rect 514260 358776 514266 358788
rect 555234 358776 555240 358788
rect 555292 358776 555298 358828
rect 549898 358708 549904 358760
rect 549956 358748 549962 358760
rect 556706 358748 556712 358760
rect 549956 358720 556712 358748
rect 549956 358708 549962 358720
rect 556706 358708 556712 358720
rect 556764 358708 556770 358760
rect 519630 358640 519636 358692
rect 519688 358680 519694 358692
rect 564066 358680 564072 358692
rect 519688 358652 564072 358680
rect 519688 358640 519694 358652
rect 564066 358640 564072 358652
rect 564124 358640 564130 358692
rect 518342 358572 518348 358624
rect 518400 358612 518406 358624
rect 562594 358612 562600 358624
rect 518400 358584 562600 358612
rect 518400 358572 518406 358584
rect 562594 358572 562600 358584
rect 562652 358572 562658 358624
rect 547230 358504 547236 358556
rect 547288 358544 547294 358556
rect 559650 358544 559656 358556
rect 547288 358516 559656 358544
rect 547288 358504 547294 358516
rect 559650 358504 559656 358516
rect 559708 358504 559714 358556
rect 515582 358436 515588 358488
rect 515640 358476 515646 358488
rect 561122 358476 561128 358488
rect 515640 358448 561128 358476
rect 515640 358436 515646 358448
rect 561122 358436 561128 358448
rect 561180 358436 561186 358488
rect 512914 356192 512920 356244
rect 512972 356232 512978 356244
rect 516502 356232 516508 356244
rect 512972 356204 516508 356232
rect 512972 356192 512978 356204
rect 516502 356192 516508 356204
rect 516560 356192 516566 356244
rect 513282 355104 513288 355156
rect 513340 355144 513346 355156
rect 517514 355144 517520 355156
rect 513340 355116 517520 355144
rect 513340 355104 513346 355116
rect 517514 355104 517520 355116
rect 517572 355104 517578 355156
rect 445570 354220 445576 354272
rect 445628 354260 445634 354272
rect 447318 354260 447324 354272
rect 445628 354232 447324 354260
rect 445628 354220 445634 354232
rect 447318 354220 447324 354232
rect 447376 354220 447382 354272
rect 512362 353608 512368 353660
rect 512420 353648 512426 353660
rect 515030 353648 515036 353660
rect 512420 353620 515036 353648
rect 512420 353608 512426 353620
rect 515030 353608 515036 353620
rect 515088 353608 515094 353660
rect 512822 353064 512828 353116
rect 512880 353104 512886 353116
rect 517606 353104 517612 353116
rect 512880 353076 517612 353104
rect 512880 353064 512886 353076
rect 517606 353064 517612 353076
rect 517664 353064 517670 353116
rect 512362 352384 512368 352436
rect 512420 352424 512426 352436
rect 515214 352424 515220 352436
rect 512420 352396 515220 352424
rect 512420 352384 512426 352396
rect 515214 352384 515220 352396
rect 515272 352384 515278 352436
rect 511442 352112 511448 352164
rect 511500 352152 511506 352164
rect 580166 352152 580172 352164
rect 511500 352124 580172 352152
rect 511500 352112 511506 352124
rect 580166 352112 580172 352124
rect 580224 352112 580230 352164
rect 513282 351976 513288 352028
rect 513340 352016 513346 352028
rect 519354 352016 519360 352028
rect 513340 351988 519360 352016
rect 513340 351976 513346 351988
rect 519354 351976 519360 351988
rect 519412 351976 519418 352028
rect 512362 350888 512368 350940
rect 512420 350928 512426 350940
rect 515306 350928 515312 350940
rect 512420 350900 515312 350928
rect 512420 350888 512426 350900
rect 515306 350888 515312 350900
rect 515364 350888 515370 350940
rect 513006 350616 513012 350668
rect 513064 350656 513070 350668
rect 517698 350656 517704 350668
rect 513064 350628 517704 350656
rect 513064 350616 513070 350628
rect 517698 350616 517704 350628
rect 517756 350616 517762 350668
rect 405734 350548 405740 350600
rect 405792 350588 405798 350600
rect 447134 350588 447140 350600
rect 405792 350560 447140 350588
rect 405792 350548 405798 350560
rect 447134 350548 447140 350560
rect 447192 350548 447198 350600
rect 513190 349528 513196 349580
rect 513248 349568 513254 349580
rect 520642 349568 520648 349580
rect 513248 349540 520648 349568
rect 513248 349528 513254 349540
rect 520642 349528 520648 349540
rect 520700 349528 520706 349580
rect 512362 349256 512368 349308
rect 512420 349296 512426 349308
rect 513926 349296 513932 349308
rect 512420 349268 513932 349296
rect 512420 349256 512426 349268
rect 513926 349256 513932 349268
rect 513984 349256 513990 349308
rect 513006 349188 513012 349240
rect 513064 349228 513070 349240
rect 516594 349228 516600 349240
rect 513064 349200 516600 349228
rect 513064 349188 513070 349200
rect 516594 349188 516600 349200
rect 516652 349188 516658 349240
rect 513006 348032 513012 348084
rect 513064 348072 513070 348084
rect 517790 348072 517796 348084
rect 513064 348044 517796 348072
rect 513064 348032 513070 348044
rect 517790 348032 517796 348044
rect 517848 348032 517854 348084
rect 361758 347760 361764 347812
rect 361816 347800 361822 347812
rect 402238 347800 402244 347812
rect 361816 347772 402244 347800
rect 361816 347760 361822 347772
rect 402238 347760 402244 347772
rect 402296 347760 402302 347812
rect 362218 347692 362224 347744
rect 362276 347732 362282 347744
rect 447134 347732 447140 347744
rect 362276 347704 447140 347732
rect 362276 347692 362282 347704
rect 447134 347692 447140 347704
rect 447192 347692 447198 347744
rect 513282 346672 513288 346724
rect 513340 346712 513346 346724
rect 519446 346712 519452 346724
rect 513340 346684 519452 346712
rect 513340 346672 513346 346684
rect 519446 346672 519452 346684
rect 519504 346672 519510 346724
rect 513098 346536 513104 346588
rect 513156 346576 513162 346588
rect 516870 346576 516876 346588
rect 513156 346548 516876 346576
rect 513156 346536 513162 346548
rect 516870 346536 516876 346548
rect 516928 346536 516934 346588
rect 446214 344904 446220 344956
rect 446272 344944 446278 344956
rect 448422 344944 448428 344956
rect 446272 344916 448428 344944
rect 446272 344904 446278 344916
rect 448422 344904 448428 344916
rect 448480 344904 448486 344956
rect 432690 344292 432696 344344
rect 432748 344332 432754 344344
rect 442258 344332 442264 344344
rect 432748 344304 442264 344332
rect 432748 344292 432754 344304
rect 442258 344292 442264 344304
rect 442316 344292 442322 344344
rect 447318 344224 447324 344276
rect 447376 344264 447382 344276
rect 447502 344264 447508 344276
rect 447376 344236 447508 344264
rect 447376 344224 447382 344236
rect 447502 344224 447508 344236
rect 447560 344224 447566 344276
rect 436830 343884 436836 343936
rect 436888 343924 436894 343936
rect 439130 343924 439136 343936
rect 436888 343896 439136 343924
rect 436888 343884 436894 343896
rect 439130 343884 439136 343896
rect 439188 343884 439194 343936
rect 512638 343680 512644 343732
rect 512696 343720 512702 343732
rect 520734 343720 520740 343732
rect 512696 343692 520740 343720
rect 512696 343680 512702 343692
rect 520734 343680 520740 343692
rect 520792 343680 520798 343732
rect 513006 343136 513012 343188
rect 513064 343176 513070 343188
rect 517882 343176 517888 343188
rect 513064 343148 517888 343176
rect 513064 343136 513070 343148
rect 517882 343136 517888 343148
rect 517940 343136 517946 343188
rect 402238 342864 402244 342916
rect 402296 342904 402302 342916
rect 447502 342904 447508 342916
rect 402296 342876 447508 342904
rect 402296 342864 402302 342876
rect 447502 342864 447508 342876
rect 447560 342864 447566 342916
rect 513282 342252 513288 342304
rect 513340 342292 513346 342304
rect 521838 342292 521844 342304
rect 513340 342264 521844 342292
rect 513340 342252 513346 342264
rect 521838 342252 521844 342264
rect 521896 342252 521902 342304
rect 447226 342184 447232 342236
rect 447284 342224 447290 342236
rect 447594 342224 447600 342236
rect 447284 342196 447600 342224
rect 447284 342184 447290 342196
rect 447594 342184 447600 342196
rect 447652 342184 447658 342236
rect 513006 341096 513012 341148
rect 513064 341136 513070 341148
rect 516686 341136 516692 341148
rect 513064 341108 516692 341136
rect 513064 341096 513070 341108
rect 516686 341096 516692 341108
rect 516744 341096 516750 341148
rect 418154 340960 418160 341012
rect 418212 341000 418218 341012
rect 447134 341000 447140 341012
rect 418212 340972 447140 341000
rect 418212 340960 418218 340972
rect 447134 340960 447140 340972
rect 447192 340960 447198 341012
rect 513282 340960 513288 341012
rect 513340 341000 513346 341012
rect 517974 341000 517980 341012
rect 513340 340972 517980 341000
rect 513340 340960 513346 340972
rect 517974 340960 517980 340972
rect 518032 340960 518038 341012
rect 361758 340892 361764 340944
rect 361816 340932 361822 340944
rect 447226 340932 447232 340944
rect 361816 340904 447232 340932
rect 361816 340892 361822 340904
rect 447226 340892 447232 340904
rect 447284 340892 447290 340944
rect 513282 339600 513288 339652
rect 513340 339640 513346 339652
rect 519630 339640 519636 339652
rect 513340 339612 519636 339640
rect 513340 339600 513346 339612
rect 519630 339600 519636 339612
rect 519688 339600 519694 339652
rect 443730 339532 443736 339584
rect 443788 339572 443794 339584
rect 447226 339572 447232 339584
rect 443788 339544 447232 339572
rect 443788 339532 443794 339544
rect 447226 339532 447232 339544
rect 447284 339532 447290 339584
rect 513098 339532 513104 339584
rect 513156 339572 513162 339584
rect 518066 339572 518072 339584
rect 513156 339544 518072 339572
rect 513156 339532 513162 339544
rect 518066 339532 518072 339544
rect 518124 339532 518130 339584
rect 399478 339464 399484 339516
rect 399536 339504 399542 339516
rect 447134 339504 447140 339516
rect 399536 339476 447140 339504
rect 399536 339464 399542 339476
rect 447134 339464 447140 339476
rect 447192 339464 447198 339516
rect 513190 339464 513196 339516
rect 513248 339504 513254 339516
rect 521930 339504 521936 339516
rect 513248 339476 521936 339504
rect 513248 339464 513254 339476
rect 521930 339464 521936 339476
rect 521988 339464 521994 339516
rect 512638 338240 512644 338292
rect 512696 338280 512702 338292
rect 520826 338280 520832 338292
rect 512696 338252 520832 338280
rect 512696 338240 512702 338252
rect 520826 338240 520832 338252
rect 520884 338240 520890 338292
rect 436830 338172 436836 338224
rect 436888 338212 436894 338224
rect 447134 338212 447140 338224
rect 436888 338184 447140 338212
rect 436888 338172 436894 338184
rect 447134 338172 447140 338184
rect 447192 338172 447198 338224
rect 385678 338104 385684 338156
rect 385736 338144 385742 338156
rect 447226 338144 447232 338156
rect 385736 338116 447232 338144
rect 385736 338104 385742 338116
rect 447226 338104 447232 338116
rect 447284 338104 447290 338156
rect 512822 338104 512828 338156
rect 512880 338144 512886 338156
rect 522022 338144 522028 338156
rect 512880 338116 522028 338144
rect 512880 338104 512886 338116
rect 522022 338104 522028 338116
rect 522080 338104 522086 338156
rect 439130 338036 439136 338088
rect 439188 338076 439194 338088
rect 441246 338076 441252 338088
rect 439188 338048 441252 338076
rect 439188 338036 439194 338048
rect 441246 338036 441252 338048
rect 441304 338036 441310 338088
rect 362218 337356 362224 337408
rect 362276 337396 362282 337408
rect 418154 337396 418160 337408
rect 362276 337368 418160 337396
rect 362276 337356 362282 337368
rect 418154 337356 418160 337368
rect 418212 337356 418218 337408
rect 513282 337016 513288 337068
rect 513340 337056 513346 337068
rect 518342 337056 518348 337068
rect 513340 337028 518348 337056
rect 513340 337016 513346 337028
rect 518342 337016 518348 337028
rect 518400 337016 518406 337068
rect 513282 336880 513288 336932
rect 513340 336920 513346 336932
rect 519722 336920 519728 336932
rect 513340 336892 519728 336920
rect 513340 336880 513346 336892
rect 519722 336880 519728 336892
rect 519780 336880 519786 336932
rect 420454 336812 420460 336864
rect 420512 336852 420518 336864
rect 429838 336852 429844 336864
rect 420512 336824 429844 336852
rect 420512 336812 420518 336824
rect 429838 336812 429844 336824
rect 429896 336812 429902 336864
rect 431218 336812 431224 336864
rect 431276 336852 431282 336864
rect 447226 336852 447232 336864
rect 431276 336824 447232 336852
rect 431276 336812 431282 336824
rect 447226 336812 447232 336824
rect 447284 336812 447290 336864
rect 416774 336744 416780 336796
rect 416832 336784 416838 336796
rect 439866 336784 439872 336796
rect 416832 336756 439872 336784
rect 416832 336744 416838 336756
rect 439866 336744 439872 336756
rect 439924 336744 439930 336796
rect 440970 336744 440976 336796
rect 441028 336784 441034 336796
rect 447134 336784 447140 336796
rect 441028 336756 447140 336784
rect 441028 336744 441034 336756
rect 447134 336744 447140 336756
rect 447192 336744 447198 336796
rect 418798 336200 418804 336252
rect 418856 336240 418862 336252
rect 438118 336240 438124 336252
rect 418856 336212 438124 336240
rect 418856 336200 418862 336212
rect 438118 336200 438124 336212
rect 438176 336200 438182 336252
rect 418890 336132 418896 336184
rect 418948 336172 418954 336184
rect 441338 336172 441344 336184
rect 418948 336144 441344 336172
rect 418948 336132 418954 336144
rect 441338 336132 441344 336144
rect 441396 336132 441402 336184
rect 412634 336064 412640 336116
rect 412692 336104 412698 336116
rect 449434 336104 449440 336116
rect 412692 336076 449440 336104
rect 412692 336064 412698 336076
rect 449434 336064 449440 336076
rect 449492 336064 449498 336116
rect 397454 335996 397460 336048
rect 397512 336036 397518 336048
rect 441154 336036 441160 336048
rect 397512 336008 441160 336036
rect 397512 335996 397518 336008
rect 441154 335996 441160 336008
rect 441212 335996 441218 336048
rect 413094 335384 413100 335436
rect 413152 335424 413158 335436
rect 435542 335424 435548 335436
rect 413152 335396 435548 335424
rect 413152 335384 413158 335396
rect 435542 335384 435548 335396
rect 435600 335384 435606 335436
rect 439774 335384 439780 335436
rect 439832 335424 439838 335436
rect 447134 335424 447140 335436
rect 439832 335396 447140 335424
rect 439832 335384 439838 335396
rect 447134 335384 447140 335396
rect 447192 335384 447198 335436
rect 409414 335316 409420 335368
rect 409472 335356 409478 335368
rect 431310 335356 431316 335368
rect 409472 335328 431316 335356
rect 409472 335316 409478 335328
rect 431310 335316 431316 335328
rect 431368 335316 431374 335368
rect 435358 335316 435364 335368
rect 435416 335356 435422 335368
rect 447226 335356 447232 335368
rect 435416 335328 447232 335356
rect 435416 335316 435422 335328
rect 447226 335316 447232 335328
rect 447284 335316 447290 335368
rect 420362 335044 420368 335096
rect 420420 335044 420426 335096
rect 420822 335044 420828 335096
rect 420880 335084 420886 335096
rect 443822 335084 443828 335096
rect 420880 335056 443828 335084
rect 420880 335044 420886 335056
rect 443822 335044 443828 335056
rect 443880 335044 443886 335096
rect 420380 335016 420408 335044
rect 443914 335016 443920 335028
rect 420380 334988 443920 335016
rect 443914 334976 443920 334988
rect 443972 334976 443978 335028
rect 420730 334908 420736 334960
rect 420788 334948 420794 334960
rect 446214 334948 446220 334960
rect 420788 334920 446220 334948
rect 420788 334908 420794 334920
rect 446214 334908 446220 334920
rect 446272 334908 446278 334960
rect 417418 334840 417424 334892
rect 417476 334880 417482 334892
rect 444006 334880 444012 334892
rect 417476 334852 444012 334880
rect 417476 334840 417482 334852
rect 444006 334840 444012 334852
rect 444064 334840 444070 334892
rect 420178 334772 420184 334824
rect 420236 334812 420242 334824
rect 449066 334812 449072 334824
rect 420236 334784 449072 334812
rect 420236 334772 420242 334784
rect 449066 334772 449072 334784
rect 449124 334772 449130 334824
rect 420546 334704 420552 334756
rect 420604 334744 420610 334756
rect 450446 334744 450452 334756
rect 420604 334716 450452 334744
rect 420604 334704 420610 334716
rect 450446 334704 450452 334716
rect 450504 334704 450510 334756
rect 420638 334636 420644 334688
rect 420696 334676 420702 334688
rect 450722 334676 450728 334688
rect 420696 334648 450728 334676
rect 420696 334636 420702 334648
rect 450722 334636 450728 334648
rect 450780 334636 450786 334688
rect 420270 334568 420276 334620
rect 420328 334608 420334 334620
rect 450630 334608 450636 334620
rect 420328 334580 450636 334608
rect 420328 334568 420334 334580
rect 450630 334568 450636 334580
rect 450688 334568 450694 334620
rect 428090 334364 428096 334416
rect 428148 334404 428154 334416
rect 428148 334376 431954 334404
rect 428148 334364 428154 334376
rect 431926 334132 431954 334376
rect 512730 334296 512736 334348
rect 512788 334336 512794 334348
rect 514754 334336 514760 334348
rect 512788 334308 514760 334336
rect 512788 334296 512794 334308
rect 514754 334296 514760 334308
rect 514812 334296 514818 334348
rect 447410 334132 447416 334144
rect 431926 334104 447416 334132
rect 447410 334092 447416 334104
rect 447468 334092 447474 334144
rect 442258 334024 442264 334076
rect 442316 334064 442322 334076
rect 447502 334064 447508 334076
rect 442316 334036 447508 334064
rect 442316 334024 442322 334036
rect 447502 334024 447508 334036
rect 447560 334024 447566 334076
rect 363598 333956 363604 334008
rect 363656 333996 363662 334008
rect 447226 333996 447232 334008
rect 363656 333968 447232 333996
rect 363656 333956 363662 333968
rect 447226 333956 447232 333968
rect 447284 333956 447290 334008
rect 439498 332800 439504 332852
rect 439556 332840 439562 332852
rect 447134 332840 447140 332852
rect 439556 332812 447140 332840
rect 439556 332800 439562 332812
rect 447134 332800 447140 332812
rect 447192 332800 447198 332852
rect 447410 332772 447416 332784
rect 443472 332744 447416 332772
rect 436738 332664 436744 332716
rect 436796 332704 436802 332716
rect 436796 332676 441614 332704
rect 436796 332664 436802 332676
rect 432966 332596 432972 332648
rect 433024 332636 433030 332648
rect 437014 332636 437020 332648
rect 433024 332608 437020 332636
rect 433024 332596 433030 332608
rect 437014 332596 437020 332608
rect 437072 332596 437078 332648
rect 441586 332636 441614 332676
rect 443472 332636 443500 332744
rect 447410 332732 447416 332744
rect 447468 332732 447474 332784
rect 441586 332608 443500 332636
rect 443638 332596 443644 332648
rect 443696 332636 443702 332648
rect 447226 332636 447232 332648
rect 443696 332608 447232 332636
rect 443696 332596 443702 332608
rect 447226 332596 447232 332608
rect 447284 332596 447290 332648
rect 512914 331440 512920 331492
rect 512972 331480 512978 331492
rect 516410 331480 516416 331492
rect 512972 331452 516416 331480
rect 512972 331440 512978 331452
rect 516410 331440 516416 331452
rect 516468 331440 516474 331492
rect 444098 331304 444104 331356
rect 444156 331344 444162 331356
rect 444282 331344 444288 331356
rect 444156 331316 444288 331344
rect 444156 331304 444162 331316
rect 444282 331304 444288 331316
rect 444340 331344 444346 331356
rect 447226 331344 447232 331356
rect 444340 331316 447232 331344
rect 444340 331304 444346 331316
rect 447226 331304 447232 331316
rect 447284 331304 447290 331356
rect 432782 331236 432788 331288
rect 432840 331276 432846 331288
rect 439682 331276 439688 331288
rect 432840 331248 439688 331276
rect 432840 331236 432846 331248
rect 439682 331236 439688 331248
rect 439740 331236 439746 331288
rect 440878 331236 440884 331288
rect 440936 331276 440942 331288
rect 447134 331276 447140 331288
rect 440936 331248 447140 331276
rect 440936 331236 440942 331248
rect 447134 331236 447140 331248
rect 447192 331236 447198 331288
rect 442902 330556 442908 330608
rect 442960 330596 442966 330608
rect 444374 330596 444380 330608
rect 442960 330568 444380 330596
rect 442960 330556 442966 330568
rect 444374 330556 444380 330568
rect 444432 330596 444438 330608
rect 447134 330596 447140 330608
rect 444432 330568 447140 330596
rect 444432 330556 444438 330568
rect 447134 330556 447140 330568
rect 447192 330556 447198 330608
rect 438762 330488 438768 330540
rect 438820 330528 438826 330540
rect 447594 330528 447600 330540
rect 438820 330500 447600 330528
rect 438820 330488 438826 330500
rect 447594 330488 447600 330500
rect 447652 330488 447658 330540
rect 432598 330012 432604 330064
rect 432656 330052 432662 330064
rect 435450 330052 435456 330064
rect 432656 330024 435456 330052
rect 432656 330012 432662 330024
rect 435450 330012 435456 330024
rect 435508 330012 435514 330064
rect 431862 329060 431868 329112
rect 431920 329100 431926 329112
rect 447410 329100 447416 329112
rect 431920 329072 447416 329100
rect 431920 329060 431926 329072
rect 447410 329060 447416 329072
rect 447468 329060 447474 329112
rect 436002 328448 436008 328500
rect 436060 328488 436066 328500
rect 447134 328488 447140 328500
rect 436060 328460 447140 328488
rect 436060 328448 436066 328460
rect 447134 328448 447140 328460
rect 447192 328448 447198 328500
rect 429194 328380 429200 328432
rect 429252 328420 429258 328432
rect 448238 328420 448244 328432
rect 429252 328392 448244 328420
rect 429252 328380 429258 328392
rect 448238 328380 448244 328392
rect 448296 328380 448302 328432
rect 429838 327020 429844 327072
rect 429896 327060 429902 327072
rect 447410 327060 447416 327072
rect 429896 327032 447416 327060
rect 429896 327020 429902 327032
rect 447410 327020 447416 327032
rect 447468 327060 447474 327072
rect 448146 327060 448152 327072
rect 447468 327032 448152 327060
rect 447468 327020 447474 327032
rect 448146 327020 448152 327032
rect 448204 327020 448210 327072
rect 439866 326952 439872 327004
rect 439924 326992 439930 327004
rect 447962 326992 447968 327004
rect 439924 326964 447968 326992
rect 439924 326952 439930 326964
rect 447962 326952 447968 326964
rect 448020 326952 448026 327004
rect 435542 325524 435548 325576
rect 435600 325564 435606 325576
rect 448054 325564 448060 325576
rect 435600 325536 448060 325564
rect 435600 325524 435606 325536
rect 448054 325524 448060 325536
rect 448112 325524 448118 325576
rect 431310 324912 431316 324964
rect 431368 324952 431374 324964
rect 448330 324952 448336 324964
rect 431368 324924 448336 324952
rect 431368 324912 431374 324924
rect 448330 324912 448336 324924
rect 448388 324952 448394 324964
rect 449526 324952 449532 324964
rect 448388 324924 449532 324952
rect 448388 324912 448394 324924
rect 449526 324912 449532 324924
rect 449584 324912 449590 324964
rect 432690 323552 432696 323604
rect 432748 323592 432754 323604
rect 442350 323592 442356 323604
rect 432748 323564 442356 323592
rect 432748 323552 432754 323564
rect 442350 323552 442356 323564
rect 442408 323552 442414 323604
rect 509694 323416 509700 323468
rect 509752 323456 509758 323468
rect 510246 323456 510252 323468
rect 509752 323428 510252 323456
rect 509752 323416 509758 323428
rect 510246 323416 510252 323428
rect 510304 323416 510310 323468
rect 507486 322668 507492 322720
rect 507544 322708 507550 322720
rect 510062 322708 510068 322720
rect 507544 322680 510068 322708
rect 507544 322668 507550 322680
rect 510062 322668 510068 322680
rect 510120 322668 510126 322720
rect 507578 322600 507584 322652
rect 507636 322640 507642 322652
rect 509602 322640 509608 322652
rect 507636 322612 509608 322640
rect 507636 322600 507642 322612
rect 509602 322600 509608 322612
rect 509660 322600 509666 322652
rect 507394 322532 507400 322584
rect 507452 322572 507458 322584
rect 510154 322572 510160 322584
rect 507452 322544 510160 322572
rect 507452 322532 507458 322544
rect 510154 322532 510160 322544
rect 510212 322532 510218 322584
rect 507302 322464 507308 322516
rect 507360 322504 507366 322516
rect 509970 322504 509976 322516
rect 507360 322476 509976 322504
rect 507360 322464 507366 322476
rect 509970 322464 509976 322476
rect 510028 322464 510034 322516
rect 463510 322436 463516 322448
rect 451246 322408 463516 322436
rect 450446 322328 450452 322380
rect 450504 322368 450510 322380
rect 451246 322368 451274 322408
rect 463510 322396 463516 322408
rect 463568 322396 463574 322448
rect 507118 322396 507124 322448
rect 507176 322436 507182 322448
rect 511166 322436 511172 322448
rect 507176 322408 511172 322436
rect 507176 322396 507182 322408
rect 511166 322396 511172 322408
rect 511224 322396 511230 322448
rect 464890 322368 464896 322380
rect 450504 322340 451274 322368
rect 456766 322340 464896 322368
rect 450504 322328 450510 322340
rect 441246 322260 441252 322312
rect 441304 322300 441310 322312
rect 456766 322300 456794 322340
rect 464890 322328 464896 322340
rect 464948 322328 464954 322380
rect 441304 322272 456794 322300
rect 441304 322260 441310 322272
rect 459646 322260 459652 322312
rect 459704 322300 459710 322312
rect 463510 322300 463516 322312
rect 459704 322272 463516 322300
rect 459704 322260 459710 322272
rect 463510 322260 463516 322272
rect 463568 322260 463574 322312
rect 443914 322192 443920 322244
rect 443972 322232 443978 322244
rect 463234 322232 463240 322244
rect 443972 322204 463240 322232
rect 443972 322192 443978 322204
rect 463234 322192 463240 322204
rect 463292 322192 463298 322244
rect 502150 322192 502156 322244
rect 502208 322232 502214 322244
rect 580442 322232 580448 322244
rect 502208 322204 580448 322232
rect 502208 322192 502214 322204
rect 580442 322192 580448 322204
rect 580500 322192 580506 322244
rect 449250 322124 449256 322176
rect 449308 322164 449314 322176
rect 471790 322164 471796 322176
rect 449308 322136 471796 322164
rect 449308 322124 449314 322136
rect 471790 322124 471796 322136
rect 471848 322124 471854 322176
rect 450722 322056 450728 322108
rect 450780 322096 450786 322108
rect 484210 322096 484216 322108
rect 450780 322068 484216 322096
rect 450780 322056 450786 322068
rect 484210 322056 484216 322068
rect 484268 322056 484274 322108
rect 445662 321988 445668 322040
rect 445720 322028 445726 322040
rect 481174 322028 481180 322040
rect 445720 322000 481180 322028
rect 445720 321988 445726 322000
rect 481174 321988 481180 322000
rect 481232 321988 481238 322040
rect 446214 321920 446220 321972
rect 446272 321960 446278 321972
rect 483934 321960 483940 321972
rect 446272 321932 483940 321960
rect 446272 321920 446278 321932
rect 483934 321920 483940 321932
rect 483992 321920 483998 321972
rect 449066 321852 449072 321904
rect 449124 321892 449130 321904
rect 474090 321892 474096 321904
rect 449124 321864 474096 321892
rect 449124 321852 449130 321864
rect 474090 321852 474096 321864
rect 474148 321852 474154 321904
rect 479610 321852 479616 321904
rect 479668 321892 479674 321904
rect 518158 321892 518164 321904
rect 479668 321864 518164 321892
rect 479668 321852 479674 321864
rect 518158 321852 518164 321864
rect 518216 321852 518222 321904
rect 444006 321784 444012 321836
rect 444064 321824 444070 321836
rect 463878 321824 463884 321836
rect 444064 321796 463884 321824
rect 444064 321784 444070 321796
rect 463878 321784 463884 321796
rect 463936 321784 463942 321836
rect 469122 321784 469128 321836
rect 469180 321824 469186 321836
rect 518250 321824 518256 321836
rect 469180 321796 518256 321824
rect 469180 321784 469186 321796
rect 518250 321784 518256 321796
rect 518308 321784 518314 321836
rect 459186 321716 459192 321768
rect 459244 321756 459250 321768
rect 515490 321756 515496 321768
rect 459244 321728 515496 321756
rect 459244 321716 459250 321728
rect 515490 321716 515496 321728
rect 515548 321716 515554 321768
rect 449158 321648 449164 321700
rect 449216 321688 449222 321700
rect 460566 321688 460572 321700
rect 449216 321660 460572 321688
rect 449216 321648 449222 321660
rect 460566 321648 460572 321660
rect 460624 321648 460630 321700
rect 567838 321688 567844 321700
rect 463068 321660 567844 321688
rect 459738 321580 459744 321632
rect 459796 321620 459802 321632
rect 463068 321620 463096 321660
rect 567838 321648 567844 321660
rect 567896 321648 567902 321700
rect 459796 321592 463096 321620
rect 459796 321580 459802 321592
rect 463510 321580 463516 321632
rect 463568 321620 463574 321632
rect 580258 321620 580264 321632
rect 463568 321592 580264 321620
rect 463568 321580 463574 321592
rect 580258 321580 580264 321592
rect 580316 321580 580322 321632
rect 458910 321512 458916 321564
rect 458968 321552 458974 321564
rect 580534 321552 580540 321564
rect 458968 321524 580540 321552
rect 458968 321512 458974 321524
rect 580534 321512 580540 321524
rect 580592 321512 580598 321564
rect 445018 321444 445024 321496
rect 445076 321484 445082 321496
rect 460842 321484 460848 321496
rect 445076 321456 460848 321484
rect 445076 321444 445082 321456
rect 460842 321444 460848 321456
rect 460900 321444 460906 321496
rect 470226 321444 470232 321496
rect 470284 321484 470290 321496
rect 576118 321484 576124 321496
rect 470284 321456 576124 321484
rect 470284 321444 470290 321456
rect 576118 321444 576124 321456
rect 576176 321444 576182 321496
rect 450538 321376 450544 321428
rect 450596 321416 450602 321428
rect 461394 321416 461400 321428
rect 450596 321388 461400 321416
rect 450596 321376 450602 321388
rect 461394 321376 461400 321388
rect 461452 321376 461458 321428
rect 469950 321376 469956 321428
rect 470008 321416 470014 321428
rect 574738 321416 574744 321428
rect 470008 321388 574744 321416
rect 470008 321376 470014 321388
rect 574738 321376 574744 321388
rect 574796 321376 574802 321428
rect 445478 321308 445484 321360
rect 445536 321348 445542 321360
rect 462498 321348 462504 321360
rect 445536 321320 462504 321348
rect 445536 321308 445542 321320
rect 462498 321308 462504 321320
rect 462556 321308 462562 321360
rect 468570 321308 468576 321360
rect 468628 321348 468634 321360
rect 569218 321348 569224 321360
rect 468628 321320 569224 321348
rect 468628 321308 468634 321320
rect 569218 321308 569224 321320
rect 569276 321308 569282 321360
rect 480714 321240 480720 321292
rect 480772 321280 480778 321292
rect 573358 321280 573364 321292
rect 480772 321252 573364 321280
rect 480772 321240 480778 321252
rect 573358 321240 573364 321252
rect 573416 321240 573422 321292
rect 458082 321172 458088 321224
rect 458140 321212 458146 321224
rect 511442 321212 511448 321224
rect 458140 321184 511448 321212
rect 458140 321172 458146 321184
rect 511442 321172 511448 321184
rect 511500 321172 511506 321224
rect 458358 321104 458364 321156
rect 458416 321144 458422 321156
rect 511350 321144 511356 321156
rect 458416 321116 511356 321144
rect 458416 321104 458422 321116
rect 511350 321104 511356 321116
rect 511408 321104 511414 321156
rect 446398 321036 446404 321088
rect 446456 321076 446462 321088
rect 471330 321076 471336 321088
rect 446456 321048 471336 321076
rect 446456 321036 446462 321048
rect 471330 321036 471336 321048
rect 471388 321036 471394 321088
rect 479058 321036 479064 321088
rect 479116 321076 479122 321088
rect 516778 321076 516784 321088
rect 479116 321048 516784 321076
rect 479116 321036 479122 321048
rect 516778 321036 516784 321048
rect 516836 321036 516842 321088
rect 450630 320968 450636 321020
rect 450688 321008 450694 321020
rect 484578 321008 484584 321020
rect 450688 320980 484584 321008
rect 450688 320968 450694 320980
rect 484578 320968 484584 320980
rect 484636 320968 484642 321020
rect 447042 320900 447048 320952
rect 447100 320940 447106 320952
rect 473538 320940 473544 320952
rect 447100 320912 473544 320940
rect 447100 320900 447106 320912
rect 473538 320900 473544 320912
rect 473596 320900 473602 320952
rect 496814 320900 496820 320952
rect 496872 320940 496878 320952
rect 580718 320940 580724 320952
rect 496872 320912 580724 320940
rect 496872 320900 496878 320912
rect 580718 320900 580724 320912
rect 580776 320900 580782 320952
rect 461854 320832 461860 320884
rect 461912 320872 461918 320884
rect 580626 320872 580632 320884
rect 461912 320844 580632 320872
rect 461912 320832 461918 320844
rect 580626 320832 580632 320844
rect 580684 320832 580690 320884
rect 441154 320764 441160 320816
rect 441212 320804 441218 320816
rect 481542 320804 481548 320816
rect 441212 320776 481548 320804
rect 441212 320764 441218 320776
rect 481542 320764 481548 320776
rect 481600 320764 481606 320816
rect 438118 320696 438124 320748
rect 438176 320736 438182 320748
rect 472434 320736 472440 320748
rect 438176 320708 472440 320736
rect 438176 320696 438182 320708
rect 472434 320696 472440 320708
rect 472492 320696 472498 320748
rect 446950 320628 446956 320680
rect 447008 320668 447014 320680
rect 473814 320668 473820 320680
rect 447008 320640 473820 320668
rect 447008 320628 447014 320640
rect 473814 320628 473820 320640
rect 473872 320628 473878 320680
rect 445110 320560 445116 320612
rect 445168 320600 445174 320612
rect 461946 320600 461952 320612
rect 445168 320572 461952 320600
rect 445168 320560 445174 320572
rect 461946 320560 461952 320572
rect 462004 320560 462010 320612
rect 441338 320492 441344 320544
rect 441396 320532 441402 320544
rect 481818 320532 481824 320544
rect 441396 320504 481824 320532
rect 441396 320492 441402 320504
rect 481818 320492 481824 320504
rect 481876 320492 481882 320544
rect 458634 320084 458640 320136
rect 458692 320124 458698 320136
rect 461854 320124 461860 320136
rect 458692 320096 461860 320124
rect 458692 320084 458698 320096
rect 461854 320084 461860 320096
rect 461912 320084 461918 320136
rect 464890 320084 464896 320136
rect 464948 320124 464954 320136
rect 474366 320124 474372 320136
rect 464948 320096 474372 320124
rect 464948 320084 464954 320096
rect 474366 320084 474372 320096
rect 474424 320084 474430 320136
rect 479334 320084 479340 320136
rect 479392 320124 479398 320136
rect 496814 320124 496820 320136
rect 479392 320096 496820 320124
rect 479392 320084 479398 320096
rect 496814 320084 496820 320096
rect 496872 320084 496878 320136
rect 449342 320016 449348 320068
rect 449400 320056 449406 320068
rect 461118 320056 461124 320068
rect 449400 320028 461124 320056
rect 449400 320016 449406 320028
rect 461118 320016 461124 320028
rect 461176 320016 461182 320068
rect 469674 320016 469680 320068
rect 469732 320056 469738 320068
rect 580350 320056 580356 320068
rect 469732 320028 580356 320056
rect 469732 320016 469738 320028
rect 580350 320016 580356 320028
rect 580408 320016 580414 320068
rect 444190 319948 444196 320000
rect 444248 319988 444254 320000
rect 460290 319988 460296 320000
rect 444248 319960 460296 319988
rect 444248 319948 444254 319960
rect 460290 319948 460296 319960
rect 460348 319948 460354 320000
rect 478782 319948 478788 320000
rect 478840 319988 478846 320000
rect 580166 319988 580172 320000
rect 478840 319960 580172 319988
rect 478840 319948 478846 319960
rect 580166 319948 580172 319960
rect 580224 319948 580230 320000
rect 470502 319880 470508 319932
rect 470560 319920 470566 319932
rect 514110 319920 514116 319932
rect 470560 319892 514116 319920
rect 470560 319880 470566 319892
rect 514110 319880 514116 319892
rect 514168 319880 514174 319932
rect 449434 319812 449440 319864
rect 449492 319852 449498 319864
rect 471054 319852 471060 319864
rect 449492 319824 471060 319852
rect 449492 319812 449498 319824
rect 471054 319812 471060 319824
rect 471112 319812 471118 319864
rect 480990 319812 480996 319864
rect 481048 319852 481054 319864
rect 519538 319852 519544 319864
rect 481048 319824 519544 319852
rect 481048 319812 481054 319824
rect 519538 319812 519544 319824
rect 519596 319812 519602 319864
rect 443822 319744 443828 319796
rect 443880 319784 443886 319796
rect 463050 319784 463056 319796
rect 443880 319756 463056 319784
rect 443880 319744 443886 319756
rect 463050 319744 463056 319756
rect 463108 319744 463114 319796
rect 480438 319744 480444 319796
rect 480496 319784 480502 319796
rect 515398 319784 515404 319796
rect 480496 319756 515404 319784
rect 480496 319744 480502 319756
rect 515398 319744 515404 319756
rect 515456 319744 515462 319796
rect 445294 319676 445300 319728
rect 445352 319716 445358 319728
rect 462774 319716 462780 319728
rect 445352 319688 462780 319716
rect 445352 319676 445358 319688
rect 462774 319676 462780 319688
rect 462832 319676 462838 319728
rect 479886 319676 479892 319728
rect 479944 319716 479950 319728
rect 514018 319716 514024 319728
rect 479944 319688 514024 319716
rect 479944 319676 479950 319688
rect 514018 319676 514024 319688
rect 514076 319676 514082 319728
rect 458910 319608 458916 319660
rect 458968 319648 458974 319660
rect 465534 319648 465540 319660
rect 458968 319620 465540 319648
rect 458968 319608 458974 319620
rect 465534 319608 465540 319620
rect 465592 319608 465598 319660
rect 469398 319608 469404 319660
rect 469456 319648 469462 319660
rect 502150 319648 502156 319660
rect 469456 319620 502156 319648
rect 469456 319608 469462 319620
rect 502150 319608 502156 319620
rect 502208 319608 502214 319660
rect 459094 319540 459100 319592
rect 459152 319580 459158 319592
rect 476022 319580 476028 319592
rect 459152 319552 476028 319580
rect 459152 319540 459158 319552
rect 476022 319540 476028 319552
rect 476080 319540 476086 319592
rect 480162 319540 480168 319592
rect 480220 319580 480226 319592
rect 511258 319580 511264 319592
rect 480220 319552 511264 319580
rect 480220 319540 480226 319552
rect 511258 319540 511264 319552
rect 511316 319540 511322 319592
rect 460382 319472 460388 319524
rect 460440 319512 460446 319524
rect 476298 319512 476304 319524
rect 460440 319484 476304 319512
rect 460440 319472 460446 319484
rect 476298 319472 476304 319484
rect 476356 319472 476362 319524
rect 498102 319472 498108 319524
rect 498160 319512 498166 319524
rect 530670 319512 530676 319524
rect 498160 319484 530676 319512
rect 498160 319472 498166 319484
rect 530670 319472 530676 319484
rect 530728 319472 530734 319524
rect 456150 319404 456156 319456
rect 456208 319444 456214 319456
rect 486510 319444 486516 319456
rect 456208 319416 486516 319444
rect 456208 319404 456214 319416
rect 486510 319404 486516 319416
rect 486568 319404 486574 319456
rect 502794 319404 502800 319456
rect 502852 319444 502858 319456
rect 538858 319444 538864 319456
rect 502852 319416 538864 319444
rect 502852 319404 502858 319416
rect 538858 319404 538864 319416
rect 538916 319404 538922 319456
rect 460290 319336 460296 319388
rect 460348 319376 460354 319388
rect 465810 319376 465816 319388
rect 460348 319348 465816 319376
rect 460348 319336 460354 319348
rect 465810 319336 465816 319348
rect 465868 319336 465874 319388
rect 498654 319336 498660 319388
rect 498712 319376 498718 319388
rect 530578 319376 530584 319388
rect 498712 319348 530584 319376
rect 498712 319336 498718 319348
rect 530578 319336 530584 319348
rect 530636 319336 530642 319388
rect 445386 319268 445392 319320
rect 445444 319308 445450 319320
rect 473262 319308 473268 319320
rect 445444 319280 473268 319308
rect 445444 319268 445450 319280
rect 473262 319268 473268 319280
rect 473320 319268 473326 319320
rect 487246 319268 487252 319320
rect 487304 319308 487310 319320
rect 487798 319308 487804 319320
rect 487304 319280 487804 319308
rect 487304 319268 487310 319280
rect 487798 319268 487804 319280
rect 487856 319268 487862 319320
rect 494422 319268 494428 319320
rect 494480 319308 494486 319320
rect 494698 319308 494704 319320
rect 494480 319280 494704 319308
rect 494480 319268 494486 319280
rect 494698 319268 494704 319280
rect 494756 319268 494762 319320
rect 455506 319200 455512 319252
rect 455564 319240 455570 319252
rect 456334 319240 456340 319252
rect 455564 319212 456340 319240
rect 455564 319200 455570 319212
rect 456334 319200 456340 319212
rect 456392 319200 456398 319252
rect 466546 319200 466552 319252
rect 466604 319240 466610 319252
rect 467374 319240 467380 319252
rect 466604 319212 467380 319240
rect 466604 319200 466610 319212
rect 467374 319200 467380 319212
rect 467432 319200 467438 319252
rect 468846 319200 468852 319252
rect 468904 319240 468910 319252
rect 580810 319240 580816 319252
rect 468904 319212 580816 319240
rect 468904 319200 468910 319212
rect 580810 319200 580816 319212
rect 580868 319200 580874 319252
rect 446674 319132 446680 319184
rect 446732 319172 446738 319184
rect 472986 319172 472992 319184
rect 446732 319144 472992 319172
rect 446732 319132 446738 319144
rect 472986 319132 472992 319144
rect 473044 319132 473050 319184
rect 474826 319132 474832 319184
rect 474884 319172 474890 319184
rect 475102 319172 475108 319184
rect 474884 319144 475108 319172
rect 474884 319132 474890 319144
rect 475102 319132 475108 319144
rect 475160 319132 475166 319184
rect 476206 319132 476212 319184
rect 476264 319172 476270 319184
rect 477310 319172 477316 319184
rect 476264 319144 477316 319172
rect 476264 319132 476270 319144
rect 477310 319132 477316 319144
rect 477368 319132 477374 319184
rect 477586 319132 477592 319184
rect 477644 319172 477650 319184
rect 478138 319172 478144 319184
rect 477644 319144 478144 319172
rect 477644 319132 477650 319144
rect 478138 319132 478144 319144
rect 478196 319132 478202 319184
rect 446858 319064 446864 319116
rect 446916 319104 446922 319116
rect 483474 319104 483480 319116
rect 446916 319076 483480 319104
rect 446916 319064 446922 319076
rect 483474 319064 483480 319076
rect 483532 319064 483538 319116
rect 485866 319064 485872 319116
rect 485924 319104 485930 319116
rect 486970 319104 486976 319116
rect 485924 319076 486976 319104
rect 485924 319064 485930 319076
rect 486970 319064 486976 319076
rect 487028 319064 487034 319116
rect 488902 319064 488908 319116
rect 488960 319104 488966 319116
rect 489730 319104 489736 319116
rect 488960 319076 489736 319104
rect 488960 319064 488966 319076
rect 489730 319064 489736 319076
rect 489788 319064 489794 319116
rect 493042 319064 493048 319116
rect 493100 319104 493106 319116
rect 493594 319104 493600 319116
rect 493100 319076 493600 319104
rect 493100 319064 493106 319076
rect 493594 319064 493600 319076
rect 493652 319064 493658 319116
rect 495802 319064 495808 319116
rect 495860 319104 495866 319116
rect 496354 319104 496360 319116
rect 495860 319076 496360 319104
rect 495860 319064 495866 319076
rect 496354 319064 496360 319076
rect 496412 319064 496418 319116
rect 496906 319064 496912 319116
rect 496964 319104 496970 319116
rect 497182 319104 497188 319116
rect 496964 319076 497188 319104
rect 496964 319064 496970 319076
rect 497182 319064 497188 319076
rect 497240 319064 497246 319116
rect 498562 319064 498568 319116
rect 498620 319104 498626 319116
rect 499390 319104 499396 319116
rect 498620 319076 499396 319104
rect 498620 319064 498626 319076
rect 499390 319064 499396 319076
rect 499448 319064 499454 319116
rect 499666 319064 499672 319116
rect 499724 319104 499730 319116
rect 500770 319104 500776 319116
rect 499724 319076 500776 319104
rect 499724 319064 499730 319076
rect 500770 319064 500776 319076
rect 500828 319064 500834 319116
rect 501046 319064 501052 319116
rect 501104 319104 501110 319116
rect 501322 319104 501328 319116
rect 501104 319076 501328 319104
rect 501104 319064 501110 319076
rect 501322 319064 501328 319076
rect 501380 319064 501386 319116
rect 502426 319064 502432 319116
rect 502484 319104 502490 319116
rect 503530 319104 503536 319116
rect 502484 319076 503536 319104
rect 502484 319064 502490 319076
rect 503530 319064 503536 319076
rect 503588 319064 503594 319116
rect 446490 318996 446496 319048
rect 446548 319036 446554 319048
rect 482094 319036 482100 319048
rect 446548 319008 482100 319036
rect 446548 318996 446554 319008
rect 482094 318996 482100 319008
rect 482152 318996 482158 319048
rect 492766 318996 492772 319048
rect 492824 319036 492830 319048
rect 493870 319036 493876 319048
rect 492824 319008 493876 319036
rect 492824 318996 492830 319008
rect 493870 318996 493876 319008
rect 493928 318996 493934 319048
rect 495526 318996 495532 319048
rect 495584 319036 495590 319048
rect 496630 319036 496636 319048
rect 495584 319008 496636 319036
rect 495584 318996 495590 319008
rect 496630 318996 496636 319008
rect 496688 318996 496694 319048
rect 498286 318996 498292 319048
rect 498344 319036 498350 319048
rect 499114 319036 499120 319048
rect 498344 319008 499120 319036
rect 498344 318996 498350 319008
rect 499114 318996 499120 319008
rect 499172 318996 499178 319048
rect 455598 318928 455604 318980
rect 455656 318968 455662 318980
rect 456058 318968 456064 318980
rect 455656 318940 456064 318968
rect 455656 318928 455662 318940
rect 456058 318928 456064 318940
rect 456116 318928 456122 318980
rect 456886 318928 456892 318980
rect 456944 318968 456950 318980
rect 457438 318968 457444 318980
rect 456944 318940 457444 318968
rect 456944 318928 456950 318940
rect 457438 318928 457444 318940
rect 457496 318928 457502 318980
rect 466822 318928 466828 318980
rect 466880 318968 466886 318980
rect 467098 318968 467104 318980
rect 466880 318940 467104 318968
rect 466880 318928 466886 318940
rect 467098 318928 467104 318940
rect 467156 318928 467162 318980
rect 476482 318928 476488 318980
rect 476540 318968 476546 318980
rect 476758 318968 476764 318980
rect 476540 318940 476764 318968
rect 476540 318928 476546 318940
rect 476758 318928 476764 318940
rect 476816 318928 476822 318980
rect 491938 318928 491944 318980
rect 491996 318968 492002 318980
rect 492490 318968 492496 318980
rect 491996 318940 492496 318968
rect 491996 318928 492002 318940
rect 492490 318928 492496 318940
rect 492548 318928 492554 318980
rect 497182 318928 497188 318980
rect 497240 318968 497246 318980
rect 497734 318968 497740 318980
rect 497240 318940 497740 318968
rect 497240 318928 497246 318940
rect 497734 318928 497740 318940
rect 497792 318928 497798 318980
rect 455414 318860 455420 318912
rect 455472 318900 455478 318912
rect 456610 318900 456616 318912
rect 455472 318872 456616 318900
rect 455472 318860 455478 318872
rect 456610 318860 456616 318872
rect 456668 318860 456674 318912
rect 442810 318724 442816 318776
rect 442868 318764 442874 318776
rect 470778 318764 470784 318776
rect 442868 318736 470784 318764
rect 442868 318724 442874 318736
rect 470778 318724 470784 318736
rect 470836 318724 470842 318776
rect 478506 318724 478512 318776
rect 478564 318764 478570 318776
rect 479518 318764 479524 318776
rect 478564 318736 479524 318764
rect 478564 318724 478570 318736
rect 479518 318724 479524 318736
rect 479576 318724 479582 318776
rect 457806 318316 457812 318368
rect 457864 318356 457870 318368
rect 461578 318356 461584 318368
rect 457864 318328 461584 318356
rect 457864 318316 457870 318328
rect 461578 318316 461584 318328
rect 461636 318316 461642 318368
rect 459186 318248 459192 318300
rect 459244 318288 459250 318300
rect 491478 318288 491484 318300
rect 459244 318260 491484 318288
rect 459244 318248 459250 318260
rect 491478 318248 491484 318260
rect 491536 318248 491542 318300
rect 501690 318248 501696 318300
rect 501748 318288 501754 318300
rect 540330 318288 540336 318300
rect 501748 318260 540336 318288
rect 501748 318248 501754 318260
rect 540330 318248 540336 318260
rect 540388 318248 540394 318300
rect 452102 318180 452108 318232
rect 452160 318220 452166 318232
rect 495618 318220 495624 318232
rect 452160 318192 495624 318220
rect 452160 318180 452166 318192
rect 495618 318180 495624 318192
rect 495676 318180 495682 318232
rect 496170 318180 496176 318232
rect 496228 318220 496234 318232
rect 540974 318220 540980 318232
rect 496228 318192 540980 318220
rect 496228 318180 496234 318192
rect 540974 318180 540980 318192
rect 541032 318180 541038 318232
rect 458818 318112 458824 318164
rect 458876 318152 458882 318164
rect 512270 318152 512276 318164
rect 458876 318124 512276 318152
rect 458876 318112 458882 318124
rect 512270 318112 512276 318124
rect 512328 318112 512334 318164
rect 448238 318044 448244 318096
rect 448296 318084 448302 318096
rect 455230 318084 455236 318096
rect 448296 318056 455236 318084
rect 448296 318044 448302 318056
rect 455230 318044 455236 318056
rect 455288 318044 455294 318096
rect 456058 318044 456064 318096
rect 456116 318084 456122 318096
rect 512454 318084 512460 318096
rect 456116 318056 512460 318084
rect 456116 318044 456122 318056
rect 512454 318044 512460 318056
rect 512512 318044 512518 318096
rect 456334 317364 456340 317416
rect 456392 317404 456398 317416
rect 475746 317404 475752 317416
rect 456392 317376 475752 317404
rect 456392 317364 456398 317376
rect 475746 317364 475752 317376
rect 475804 317364 475810 317416
rect 456518 317296 456524 317348
rect 456576 317336 456582 317348
rect 486234 317336 486240 317348
rect 456576 317308 486240 317336
rect 456576 317296 456582 317308
rect 486234 317296 486240 317308
rect 486292 317296 486298 317348
rect 453574 317228 453580 317280
rect 453632 317268 453638 317280
rect 485682 317268 485688 317280
rect 453632 317240 485688 317268
rect 453632 317228 453638 317240
rect 485682 317228 485688 317240
rect 485740 317228 485746 317280
rect 500310 317228 500316 317280
rect 500368 317268 500374 317280
rect 539686 317268 539692 317280
rect 500368 317240 539692 317268
rect 500368 317228 500374 317240
rect 539686 317228 539692 317240
rect 539744 317228 539750 317280
rect 454770 317160 454776 317212
rect 454828 317200 454834 317212
rect 491570 317200 491576 317212
rect 454828 317172 491576 317200
rect 454828 317160 454834 317172
rect 491570 317160 491576 317172
rect 491628 317160 491634 317212
rect 502518 317160 502524 317212
rect 502576 317200 502582 317212
rect 543090 317200 543096 317212
rect 502576 317172 543096 317200
rect 502576 317160 502582 317172
rect 543090 317160 543096 317172
rect 543148 317160 543154 317212
rect 453390 317092 453396 317144
rect 453448 317132 453454 317144
rect 485958 317132 485964 317144
rect 453448 317104 485964 317132
rect 453448 317092 453454 317104
rect 485958 317092 485964 317104
rect 486016 317092 486022 317144
rect 487338 317092 487344 317144
rect 487396 317132 487402 317144
rect 529934 317132 529940 317144
rect 487396 317104 529940 317132
rect 487396 317092 487402 317104
rect 529934 317092 529940 317104
rect 529992 317092 529998 317144
rect 455046 317024 455052 317076
rect 455104 317064 455110 317076
rect 509878 317064 509884 317076
rect 455104 317036 509884 317064
rect 455104 317024 455110 317036
rect 509878 317024 509884 317036
rect 509936 317024 509942 317076
rect 456242 316956 456248 317008
rect 456300 316996 456306 317008
rect 511074 316996 511080 317008
rect 456300 316968 511080 316996
rect 456300 316956 456306 316968
rect 511074 316956 511080 316968
rect 511132 316956 511138 317008
rect 454862 316888 454868 316940
rect 454920 316928 454926 316940
rect 510246 316928 510252 316940
rect 454920 316900 510252 316928
rect 454920 316888 454926 316900
rect 510246 316888 510252 316900
rect 510304 316888 510310 316940
rect 450722 316820 450728 316872
rect 450780 316860 450786 316872
rect 509694 316860 509700 316872
rect 450780 316832 509700 316860
rect 450780 316820 450786 316832
rect 509694 316820 509700 316832
rect 509752 316820 509758 316872
rect 450630 316752 450636 316804
rect 450688 316792 450694 316804
rect 512362 316792 512368 316804
rect 450688 316764 512368 316792
rect 450688 316752 450694 316764
rect 512362 316752 512368 316764
rect 512420 316752 512426 316804
rect 450538 316684 450544 316736
rect 450596 316724 450602 316736
rect 514754 316724 514760 316736
rect 450596 316696 514760 316724
rect 450596 316684 450602 316696
rect 514754 316684 514760 316696
rect 514812 316684 514818 316736
rect 456426 316616 456432 316668
rect 456484 316656 456490 316668
rect 475470 316656 475476 316668
rect 456484 316628 475476 316656
rect 456484 316616 456490 316628
rect 475470 316616 475476 316628
rect 475528 316616 475534 316668
rect 453482 316548 453488 316600
rect 453540 316588 453546 316600
rect 464982 316588 464988 316600
rect 453540 316560 464988 316588
rect 453540 316548 453546 316560
rect 464982 316548 464988 316560
rect 465040 316548 465046 316600
rect 459002 316480 459008 316532
rect 459060 316520 459066 316532
rect 465258 316520 465264 316532
rect 459060 316492 465264 316520
rect 459060 316480 459066 316492
rect 465258 316480 465264 316492
rect 465316 316480 465322 316532
rect 361758 315936 361764 315988
rect 361816 315976 361822 315988
rect 399478 315976 399484 315988
rect 361816 315948 399484 315976
rect 361816 315936 361822 315948
rect 399478 315936 399484 315948
rect 399536 315936 399542 315988
rect 452010 315324 452016 315376
rect 452068 315364 452074 315376
rect 494146 315364 494152 315376
rect 452068 315336 494152 315364
rect 452068 315324 452074 315336
rect 494146 315324 494152 315336
rect 494204 315324 494210 315376
rect 501138 315324 501144 315376
rect 501196 315364 501202 315376
rect 541066 315364 541072 315376
rect 501196 315336 541072 315364
rect 501196 315324 501202 315336
rect 541066 315324 541072 315336
rect 541124 315324 541130 315376
rect 455690 315256 455696 315308
rect 455748 315296 455754 315308
rect 562318 315296 562324 315308
rect 455748 315268 562324 315296
rect 455748 315256 455754 315268
rect 562318 315256 562324 315268
rect 562376 315256 562382 315308
rect 451090 314236 451096 314288
rect 451148 314276 451154 314288
rect 464706 314276 464712 314288
rect 451148 314248 464712 314276
rect 451148 314236 451154 314248
rect 464706 314236 464712 314248
rect 464764 314236 464770 314288
rect 450998 314168 451004 314220
rect 451056 314208 451062 314220
rect 475010 314208 475016 314220
rect 451056 314180 475016 314208
rect 451056 314168 451062 314180
rect 475010 314168 475016 314180
rect 475068 314168 475074 314220
rect 457438 314100 457444 314152
rect 457496 314140 457502 314152
rect 485314 314140 485320 314152
rect 457496 314112 485320 314140
rect 457496 314100 457502 314112
rect 485314 314100 485320 314112
rect 485372 314100 485378 314152
rect 502978 314100 502984 314152
rect 503036 314140 503042 314152
rect 538950 314140 538956 314152
rect 503036 314112 538956 314140
rect 503036 314100 503042 314112
rect 538950 314100 538956 314112
rect 539008 314100 539014 314152
rect 452194 314032 452200 314084
rect 452252 314072 452258 314084
rect 494974 314072 494980 314084
rect 452252 314044 494980 314072
rect 452252 314032 452258 314044
rect 494974 314032 494980 314044
rect 495032 314032 495038 314084
rect 501322 314032 501328 314084
rect 501380 314072 501386 314084
rect 542998 314072 543004 314084
rect 501380 314044 543004 314072
rect 501380 314032 501386 314044
rect 542998 314032 543004 314044
rect 543056 314032 543062 314084
rect 450814 313964 450820 314016
rect 450872 314004 450878 314016
rect 513374 314004 513380 314016
rect 450872 313976 513380 314004
rect 450872 313964 450878 313976
rect 513374 313964 513380 313976
rect 513432 313964 513438 314016
rect 450906 313896 450912 313948
rect 450964 313936 450970 313948
rect 474826 313936 474832 313948
rect 450964 313908 474832 313936
rect 450964 313896 450970 313908
rect 474826 313896 474832 313908
rect 474884 313896 474890 313948
rect 476758 313896 476764 313948
rect 476816 313936 476822 313948
rect 548518 313936 548524 313948
rect 476816 313908 548524 313936
rect 476816 313896 476822 313908
rect 548518 313896 548524 313908
rect 548576 313896 548582 313948
rect 482278 313284 482284 313336
rect 482336 313324 482342 313336
rect 484486 313324 484492 313336
rect 482336 313296 484492 313324
rect 482336 313284 482342 313296
rect 484486 313284 484492 313296
rect 484544 313284 484550 313336
rect 468202 313216 468208 313268
rect 468260 313256 468266 313268
rect 580166 313256 580172 313268
rect 468260 313228 580172 313256
rect 468260 313216 468266 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 466638 312536 466644 312588
rect 466696 312576 466702 312588
rect 544378 312576 544384 312588
rect 466696 312548 544384 312576
rect 466696 312536 466702 312548
rect 544378 312536 544384 312548
rect 544436 312536 544442 312588
rect 451918 311176 451924 311228
rect 451976 311216 451982 311228
rect 489454 311216 489460 311228
rect 451976 311188 489460 311216
rect 451976 311176 451982 311188
rect 489454 311176 489460 311188
rect 489512 311176 489518 311228
rect 502702 311176 502708 311228
rect 502760 311216 502766 311228
rect 542722 311216 542728 311228
rect 502760 311188 542728 311216
rect 502760 311176 502766 311188
rect 542722 311176 542728 311188
rect 542780 311176 542786 311228
rect 432598 311108 432604 311160
rect 432656 311148 432662 311160
rect 441062 311148 441068 311160
rect 432656 311120 441068 311148
rect 432656 311108 432662 311120
rect 441062 311108 441068 311120
rect 441120 311108 441126 311160
rect 477678 311108 477684 311160
rect 477736 311148 477742 311160
rect 547138 311148 547144 311160
rect 477736 311120 547144 311148
rect 477736 311108 477742 311120
rect 547138 311108 547144 311120
rect 547196 311108 547202 311160
rect 461670 310904 461676 310956
rect 461728 310944 461734 310956
rect 463786 310944 463792 310956
rect 461728 310916 463792 310944
rect 461728 310904 461734 310916
rect 463786 310904 463792 310916
rect 463844 310904 463850 310956
rect 495526 309816 495532 309868
rect 495584 309856 495590 309868
rect 539594 309856 539600 309868
rect 495584 309828 539600 309856
rect 495584 309816 495590 309828
rect 539594 309816 539600 309828
rect 539652 309816 539658 309868
rect 453666 309748 453672 309800
rect 453724 309788 453730 309800
rect 490834 309788 490840 309800
rect 453724 309760 490840 309788
rect 453724 309748 453730 309760
rect 490834 309748 490840 309760
rect 490892 309748 490898 309800
rect 496998 309748 497004 309800
rect 497056 309788 497062 309800
rect 542906 309788 542912 309800
rect 497056 309760 542912 309788
rect 497056 309748 497062 309760
rect 542906 309748 542912 309760
rect 542964 309748 542970 309800
rect 453758 308456 453764 308508
rect 453816 308496 453822 308508
rect 491110 308496 491116 308508
rect 453816 308468 491116 308496
rect 453816 308456 453822 308468
rect 491110 308456 491116 308468
rect 491168 308456 491174 308508
rect 487798 308388 487804 308440
rect 487856 308428 487862 308440
rect 529198 308428 529204 308440
rect 487856 308400 529204 308428
rect 487856 308388 487862 308400
rect 529198 308388 529204 308400
rect 529256 308388 529262 308440
rect 432414 307708 432420 307760
rect 432472 307748 432478 307760
rect 436922 307748 436928 307760
rect 432472 307720 436928 307748
rect 432472 307708 432478 307720
rect 436922 307708 436928 307720
rect 436980 307708 436986 307760
rect 471238 307708 471244 307760
rect 471296 307748 471302 307760
rect 473722 307748 473728 307760
rect 471296 307720 473728 307748
rect 471296 307708 471302 307720
rect 473722 307708 473728 307720
rect 473780 307708 473786 307760
rect 487522 307164 487528 307216
rect 487580 307204 487586 307216
rect 530026 307204 530032 307216
rect 487580 307176 530032 307204
rect 487580 307164 487586 307176
rect 530026 307164 530032 307176
rect 530084 307164 530090 307216
rect 449618 307096 449624 307148
rect 449676 307136 449682 307148
rect 536834 307136 536840 307148
rect 449676 307108 536840 307136
rect 449676 307096 449682 307108
rect 536834 307096 536840 307108
rect 536892 307096 536898 307148
rect 465718 307028 465724 307080
rect 465776 307068 465782 307080
rect 566458 307068 566464 307080
rect 465776 307040 566464 307068
rect 465776 307028 465782 307040
rect 566458 307028 566464 307040
rect 566516 307028 566522 307080
rect 409230 306280 409236 306332
rect 409288 306320 409294 306332
rect 454954 306320 454960 306332
rect 409288 306292 454960 306320
rect 409288 306280 409294 306292
rect 454954 306280 454960 306292
rect 455012 306280 455018 306332
rect 409138 306212 409144 306264
rect 409196 306252 409202 306264
rect 455046 306252 455052 306264
rect 409196 306224 455052 306252
rect 409196 306212 409202 306224
rect 455046 306212 455052 306224
rect 455104 306212 455110 306264
rect 406746 306144 406752 306196
rect 406804 306184 406810 306196
rect 454862 306184 454868 306196
rect 406804 306156 454868 306184
rect 406804 306144 406810 306156
rect 454862 306144 454868 306156
rect 454920 306144 454926 306196
rect 457530 306144 457536 306196
rect 457588 306184 457594 306196
rect 493042 306184 493048 306196
rect 457588 306156 493048 306184
rect 457588 306144 457594 306156
rect 493042 306144 493048 306156
rect 493100 306144 493106 306196
rect 400858 306076 400864 306128
rect 400916 306116 400922 306128
rect 465442 306116 465448 306128
rect 400916 306088 465448 306116
rect 400916 306076 400922 306088
rect 465442 306076 465448 306088
rect 465500 306076 465506 306128
rect 476482 306076 476488 306128
rect 476540 306116 476546 306128
rect 565078 306116 565084 306128
rect 476540 306088 565084 306116
rect 476540 306076 476546 306088
rect 565078 306076 565084 306088
rect 565136 306076 565142 306128
rect 406470 306008 406476 306060
rect 406528 306048 406534 306060
rect 510982 306048 510988 306060
rect 406528 306020 510988 306048
rect 406528 306008 406534 306020
rect 510982 306008 510988 306020
rect 511040 306008 511046 306060
rect 403986 305940 403992 305992
rect 404044 305980 404050 305992
rect 510890 305980 510896 305992
rect 404044 305952 510896 305980
rect 404044 305940 404050 305952
rect 510890 305940 510896 305952
rect 510948 305940 510954 305992
rect 403618 305872 403624 305924
rect 403676 305912 403682 305924
rect 510798 305912 510804 305924
rect 403676 305884 510804 305912
rect 403676 305872 403682 305884
rect 510798 305872 510804 305884
rect 510856 305872 510862 305924
rect 406562 305804 406568 305856
rect 406620 305844 406626 305856
rect 513926 305844 513932 305856
rect 406620 305816 513932 305844
rect 406620 305804 406626 305816
rect 513926 305804 513932 305816
rect 513984 305804 513990 305856
rect 406654 305736 406660 305788
rect 406712 305776 406718 305788
rect 515214 305776 515220 305788
rect 406712 305748 515220 305776
rect 406712 305736 406718 305748
rect 515214 305736 515220 305748
rect 515272 305736 515278 305788
rect 406378 305668 406384 305720
rect 406436 305708 406442 305720
rect 515306 305708 515312 305720
rect 406436 305680 515312 305708
rect 406436 305668 406442 305680
rect 515306 305668 515312 305680
rect 515364 305668 515370 305720
rect 359458 305600 359464 305652
rect 359516 305640 359522 305652
rect 512546 305640 512552 305652
rect 359516 305612 512552 305640
rect 359516 305600 359522 305612
rect 512546 305600 512552 305612
rect 512604 305600 512610 305652
rect 447778 305532 447784 305584
rect 447836 305572 447842 305584
rect 464062 305572 464068 305584
rect 447836 305544 464068 305572
rect 447836 305532 447842 305544
rect 464062 305532 464068 305544
rect 464120 305532 464126 305584
rect 3602 304988 3608 305040
rect 3660 305028 3666 305040
rect 4798 305028 4804 305040
rect 3660 305000 4804 305028
rect 3660 304988 3666 305000
rect 4798 304988 4804 305000
rect 4856 304988 4862 305040
rect 361758 304920 361764 304972
rect 361816 304960 361822 304972
rect 443730 304960 443736 304972
rect 361816 304932 443736 304960
rect 361816 304920 361822 304932
rect 443730 304920 443736 304932
rect 443788 304920 443794 304972
rect 446398 304444 446404 304496
rect 446456 304484 446462 304496
rect 461670 304484 461676 304496
rect 446456 304456 461676 304484
rect 446456 304444 446462 304456
rect 461670 304444 461676 304456
rect 461728 304444 461734 304496
rect 455598 304376 455604 304428
rect 455656 304416 455662 304428
rect 563698 304416 563704 304428
rect 455656 304388 563704 304416
rect 455656 304376 455662 304388
rect 563698 304376 563704 304388
rect 563756 304376 563762 304428
rect 362218 304308 362224 304360
rect 362276 304348 362282 304360
rect 512822 304348 512828 304360
rect 362276 304320 512828 304348
rect 362276 304308 362282 304320
rect 512822 304308 512828 304320
rect 512880 304308 512886 304360
rect 360838 304240 360844 304292
rect 360896 304280 360902 304292
rect 512178 304280 512184 304292
rect 360896 304252 512184 304280
rect 360896 304240 360902 304252
rect 512178 304240 512184 304252
rect 512236 304240 512242 304292
rect 401042 303560 401048 303612
rect 401100 303600 401106 303612
rect 510614 303600 510620 303612
rect 401100 303572 510620 303600
rect 401100 303560 401106 303572
rect 510614 303560 510620 303572
rect 510672 303560 510678 303612
rect 403802 303492 403808 303544
rect 403860 303532 403866 303544
rect 513834 303532 513840 303544
rect 403860 303504 513840 303532
rect 403860 303492 403866 303504
rect 513834 303492 513840 303504
rect 513892 303492 513898 303544
rect 398374 303424 398380 303476
rect 398432 303464 398438 303476
rect 509326 303464 509332 303476
rect 398432 303436 509332 303464
rect 398432 303424 398438 303436
rect 509326 303424 509332 303436
rect 509384 303424 509390 303476
rect 401226 303356 401232 303408
rect 401284 303396 401290 303408
rect 513650 303396 513656 303408
rect 401284 303368 513656 303396
rect 401284 303356 401290 303368
rect 513650 303356 513656 303368
rect 513708 303356 513714 303408
rect 400950 303288 400956 303340
rect 401008 303328 401014 303340
rect 513742 303328 513748 303340
rect 401008 303300 513748 303328
rect 401008 303288 401014 303300
rect 513742 303288 513748 303300
rect 513800 303288 513806 303340
rect 401318 303220 401324 303272
rect 401376 303260 401382 303272
rect 515122 303260 515128 303272
rect 401376 303232 515128 303260
rect 401376 303220 401382 303232
rect 515122 303220 515128 303232
rect 515180 303220 515186 303272
rect 401134 303152 401140 303204
rect 401192 303192 401198 303204
rect 514938 303192 514944 303204
rect 401192 303164 514944 303192
rect 401192 303152 401198 303164
rect 514938 303152 514944 303164
rect 514996 303152 515002 303204
rect 398282 303084 398288 303136
rect 398340 303124 398346 303136
rect 513466 303124 513472 303136
rect 398340 303096 513472 303124
rect 398340 303084 398346 303096
rect 513466 303084 513472 303096
rect 513524 303084 513530 303136
rect 398190 303016 398196 303068
rect 398248 303056 398254 303068
rect 516318 303056 516324 303068
rect 398248 303028 516324 303056
rect 398248 303016 398254 303028
rect 516318 303016 516324 303028
rect 516376 303016 516382 303068
rect 455506 302948 455512 303000
rect 455564 302988 455570 303000
rect 574738 302988 574744 303000
rect 455564 302960 574744 302988
rect 455564 302948 455570 302960
rect 574738 302948 574744 302960
rect 574796 302948 574802 303000
rect 360930 302880 360936 302932
rect 360988 302920 360994 302932
rect 512638 302920 512644 302932
rect 360988 302892 512644 302920
rect 360988 302880 360994 302892
rect 512638 302880 512644 302892
rect 512696 302880 512702 302932
rect 403710 302812 403716 302864
rect 403768 302852 403774 302864
rect 509418 302852 509424 302864
rect 403768 302824 509424 302852
rect 403768 302812 403774 302824
rect 509418 302812 509424 302824
rect 509476 302812 509482 302864
rect 396718 302744 396724 302796
rect 396776 302784 396782 302796
rect 485866 302784 485872 302796
rect 396776 302756 485872 302784
rect 396776 302744 396782 302756
rect 485866 302744 485872 302756
rect 485924 302744 485930 302796
rect 455414 301452 455420 301504
rect 455472 301492 455478 301504
rect 576118 301492 576124 301504
rect 455472 301464 576124 301492
rect 455472 301452 455478 301464
rect 576118 301452 576124 301464
rect 576176 301452 576182 301504
rect 456978 300704 456984 300756
rect 457036 300744 457042 300756
rect 537478 300744 537484 300756
rect 457036 300716 537484 300744
rect 457036 300704 457042 300716
rect 537478 300704 537484 300716
rect 537536 300704 537542 300756
rect 398098 300636 398104 300688
rect 398156 300676 398162 300688
rect 516226 300676 516232 300688
rect 398156 300648 516232 300676
rect 398156 300636 398162 300648
rect 516226 300636 516232 300648
rect 516284 300636 516290 300688
rect 395614 300568 395620 300620
rect 395672 300608 395678 300620
rect 517974 300608 517980 300620
rect 395672 300580 517980 300608
rect 395672 300568 395678 300580
rect 517974 300568 517980 300580
rect 518032 300568 518038 300620
rect 395798 300500 395804 300552
rect 395856 300540 395862 300552
rect 518342 300540 518348 300552
rect 395856 300512 518348 300540
rect 395856 300500 395862 300512
rect 518342 300500 518348 300512
rect 518400 300500 518406 300552
rect 395430 300432 395436 300484
rect 395488 300472 395494 300484
rect 518066 300472 518072 300484
rect 395488 300444 518072 300472
rect 395488 300432 395494 300444
rect 518066 300432 518072 300444
rect 518124 300432 518130 300484
rect 392762 300364 392768 300416
rect 392820 300404 392826 300416
rect 516594 300404 516600 300416
rect 392820 300376 516600 300404
rect 392820 300364 392826 300376
rect 516594 300364 516600 300376
rect 516652 300364 516658 300416
rect 392946 300296 392952 300348
rect 393004 300336 393010 300348
rect 516870 300336 516876 300348
rect 393004 300308 516876 300336
rect 393004 300296 393010 300308
rect 516870 300296 516876 300308
rect 516928 300296 516934 300348
rect 393038 300228 393044 300280
rect 393096 300268 393102 300280
rect 517790 300268 517796 300280
rect 393096 300240 517796 300268
rect 393096 300228 393102 300240
rect 517790 300228 517796 300240
rect 517848 300228 517854 300280
rect 392670 300160 392676 300212
rect 392728 300200 392734 300212
rect 517882 300200 517888 300212
rect 392728 300172 517888 300200
rect 392728 300160 392734 300172
rect 517882 300160 517888 300172
rect 517940 300160 517946 300212
rect 361022 300092 361028 300144
rect 361080 300132 361086 300144
rect 511994 300132 512000 300144
rect 361080 300104 512000 300132
rect 361080 300092 361086 300104
rect 511994 300092 512000 300104
rect 512052 300092 512058 300144
rect 461578 299412 461584 299464
rect 461636 299452 461642 299464
rect 580166 299452 580172 299464
rect 461636 299424 580172 299452
rect 461636 299412 461642 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 457162 298052 457168 298104
rect 457220 298092 457226 298104
rect 578878 298092 578884 298104
rect 457220 298064 578884 298092
rect 457220 298052 457226 298064
rect 578878 298052 578884 298064
rect 578936 298052 578942 298104
rect 392854 297984 392860 298036
rect 392912 298024 392918 298036
rect 517698 298024 517704 298036
rect 392912 297996 517704 298024
rect 392912 297984 392918 297996
rect 517698 297984 517704 297996
rect 517756 297984 517762 298036
rect 387242 297916 387248 297968
rect 387300 297956 387306 297968
rect 514294 297956 514300 297968
rect 387300 297928 514300 297956
rect 387300 297916 387306 297928
rect 514294 297916 514300 297928
rect 514352 297916 514358 297968
rect 389910 297848 389916 297900
rect 389968 297888 389974 297900
rect 516502 297888 516508 297900
rect 389968 297860 516508 297888
rect 389968 297848 389974 297860
rect 516502 297848 516508 297860
rect 516560 297848 516566 297900
rect 390186 297780 390192 297832
rect 390244 297820 390250 297832
rect 517606 297820 517612 297832
rect 390244 297792 517612 297820
rect 390244 297780 390250 297792
rect 517606 297780 517612 297792
rect 517664 297780 517670 297832
rect 390094 297712 390100 297764
rect 390152 297752 390158 297764
rect 519262 297752 519268 297764
rect 390152 297724 519268 297752
rect 390152 297712 390158 297724
rect 519262 297712 519268 297724
rect 519320 297712 519326 297764
rect 387518 297644 387524 297696
rect 387576 297684 387582 297696
rect 519170 297684 519176 297696
rect 387576 297656 519176 297684
rect 387576 297644 387582 297656
rect 519170 297644 519176 297656
rect 519228 297644 519234 297696
rect 387334 297576 387340 297628
rect 387392 297616 387398 297628
rect 519078 297616 519084 297628
rect 387392 297588 519084 297616
rect 387392 297576 387398 297588
rect 519078 297576 519084 297588
rect 519136 297576 519142 297628
rect 387150 297508 387156 297560
rect 387208 297548 387214 297560
rect 518986 297548 518992 297560
rect 387208 297520 518992 297548
rect 387208 297508 387214 297520
rect 518986 297508 518992 297520
rect 519044 297508 519050 297560
rect 387058 297440 387064 297492
rect 387116 297480 387122 297492
rect 520550 297480 520556 297492
rect 387116 297452 520556 297480
rect 387116 297440 387122 297452
rect 520550 297440 520556 297452
rect 520608 297440 520614 297492
rect 361114 297372 361120 297424
rect 361172 297412 361178 297424
rect 512086 297412 512092 297424
rect 361172 297384 512092 297412
rect 361172 297372 361178 297384
rect 512086 297372 512092 297384
rect 512144 297372 512150 297424
rect 390002 297304 390008 297356
rect 390060 297344 390066 297356
rect 511534 297344 511540 297356
rect 390060 297316 511540 297344
rect 390060 297304 390066 297316
rect 511534 297304 511540 297316
rect 511592 297304 511598 297356
rect 390278 297236 390284 297288
rect 390336 297276 390342 297288
rect 507578 297276 507584 297288
rect 390336 297248 507584 297276
rect 390336 297236 390342 297248
rect 507578 297236 507584 297248
rect 507636 297236 507642 297288
rect 456886 295944 456892 295996
rect 456944 295984 456950 295996
rect 571978 295984 571984 295996
rect 456944 295956 571984 295984
rect 456944 295944 456950 295956
rect 571978 295944 571984 295956
rect 572036 295944 572042 295996
rect 384298 295264 384304 295316
rect 384356 295304 384362 295316
rect 507394 295304 507400 295316
rect 384356 295276 507400 295304
rect 384356 295264 384362 295276
rect 507394 295264 507400 295276
rect 507452 295264 507458 295316
rect 381906 295196 381912 295248
rect 381964 295236 381970 295248
rect 507486 295236 507492 295248
rect 381964 295208 507492 295236
rect 381964 295196 381970 295208
rect 507486 295196 507492 295208
rect 507544 295196 507550 295248
rect 384574 295128 384580 295180
rect 384632 295168 384638 295180
rect 514846 295168 514852 295180
rect 384632 295140 514852 295168
rect 384632 295128 384638 295140
rect 514846 295128 514852 295140
rect 514904 295128 514910 295180
rect 384390 295060 384396 295112
rect 384448 295100 384454 295112
rect 515674 295100 515680 295112
rect 384448 295072 515680 295100
rect 384448 295060 384454 295072
rect 515674 295060 515680 295072
rect 515732 295060 515738 295112
rect 387426 294992 387432 295044
rect 387484 295032 387490 295044
rect 520458 295032 520464 295044
rect 387484 295004 520464 295032
rect 387484 294992 387490 295004
rect 520458 294992 520464 295004
rect 520516 294992 520522 295044
rect 384482 294924 384488 294976
rect 384540 294964 384546 294976
rect 520366 294964 520372 294976
rect 384540 294936 520372 294964
rect 384540 294924 384546 294936
rect 520366 294924 520372 294936
rect 520424 294924 520430 294976
rect 381998 294856 382004 294908
rect 382056 294896 382062 294908
rect 519722 294896 519728 294908
rect 382056 294868 519728 294896
rect 382056 294856 382062 294868
rect 519722 294856 519728 294868
rect 519780 294856 519786 294908
rect 378870 294788 378876 294840
rect 378928 294828 378934 294840
rect 516686 294828 516692 294840
rect 378928 294800 516692 294828
rect 378928 294788 378934 294800
rect 516686 294788 516692 294800
rect 516744 294788 516750 294840
rect 381722 294720 381728 294772
rect 381780 294760 381786 294772
rect 520274 294760 520280 294772
rect 381780 294732 520280 294760
rect 381780 294720 381786 294732
rect 520274 294720 520280 294732
rect 520332 294720 520338 294772
rect 378962 294652 378968 294704
rect 379020 294692 379026 294704
rect 519630 294692 519636 294704
rect 379020 294664 519636 294692
rect 379020 294652 379026 294664
rect 519630 294652 519636 294664
rect 519688 294652 519694 294704
rect 379054 294584 379060 294636
rect 379112 294624 379118 294636
rect 520826 294624 520832 294636
rect 379112 294596 520832 294624
rect 379112 294584 379118 294596
rect 520826 294584 520832 294596
rect 520884 294584 520890 294636
rect 476206 294516 476212 294568
rect 476264 294556 476270 294568
rect 573358 294556 573364 294568
rect 476264 294528 573364 294556
rect 476264 294516 476270 294528
rect 573358 294516 573364 294528
rect 573416 294516 573422 294568
rect 361758 293904 361764 293956
rect 361816 293944 361822 293956
rect 385678 293944 385684 293956
rect 361816 293916 385684 293944
rect 361816 293904 361822 293916
rect 385678 293904 385684 293916
rect 385736 293904 385742 293956
rect 467098 293224 467104 293276
rect 467156 293264 467162 293276
rect 559558 293264 559564 293276
rect 467156 293236 559564 293264
rect 467156 293224 467162 293236
rect 559558 293224 559564 293236
rect 559616 293224 559622 293276
rect 3602 292544 3608 292596
rect 3660 292584 3666 292596
rect 19978 292584 19984 292596
rect 3660 292556 19984 292584
rect 3660 292544 3666 292556
rect 19978 292544 19984 292556
rect 20036 292544 20042 292596
rect 373442 292476 373448 292528
rect 373500 292516 373506 292528
rect 513558 292516 513564 292528
rect 373500 292488 513564 292516
rect 373500 292476 373506 292488
rect 513558 292476 513564 292488
rect 513616 292476 513622 292528
rect 379146 292408 379152 292460
rect 379204 292448 379210 292460
rect 519446 292448 519452 292460
rect 379204 292420 519452 292448
rect 379204 292408 379210 292420
rect 519446 292408 519452 292420
rect 519504 292408 519510 292460
rect 376478 292340 376484 292392
rect 376536 292380 376542 292392
rect 517514 292380 517520 292392
rect 376536 292352 517520 292380
rect 376536 292340 376542 292352
rect 517514 292340 517520 292352
rect 517572 292340 517578 292392
rect 379238 292272 379244 292324
rect 379296 292312 379302 292324
rect 520734 292312 520740 292324
rect 379296 292284 520740 292312
rect 379296 292272 379302 292284
rect 520734 292272 520740 292284
rect 520792 292272 520798 292324
rect 376110 292204 376116 292256
rect 376168 292244 376174 292256
rect 519354 292244 519360 292256
rect 376168 292216 519360 292244
rect 376168 292204 376174 292216
rect 519354 292204 519360 292216
rect 519412 292204 519418 292256
rect 376294 292136 376300 292188
rect 376352 292176 376358 292188
rect 520642 292176 520648 292188
rect 376352 292148 520648 292176
rect 376352 292136 376358 292148
rect 520642 292136 520648 292148
rect 520700 292136 520706 292188
rect 370682 292068 370688 292120
rect 370740 292108 370746 292120
rect 516134 292108 516140 292120
rect 370740 292080 516140 292108
rect 370740 292068 370746 292080
rect 516134 292068 516140 292080
rect 516192 292068 516198 292120
rect 370774 292000 370780 292052
rect 370832 292040 370838 292052
rect 518894 292040 518900 292052
rect 370832 292012 518900 292040
rect 370832 292000 370838 292012
rect 518894 292000 518900 292012
rect 518952 292000 518958 292052
rect 373534 291932 373540 291984
rect 373592 291972 373598 291984
rect 521746 291972 521752 291984
rect 373592 291944 521752 291972
rect 373592 291932 373598 291944
rect 521746 291932 521752 291944
rect 521804 291932 521810 291984
rect 373350 291864 373356 291916
rect 373408 291904 373414 291916
rect 523034 291904 523040 291916
rect 373408 291876 523040 291904
rect 373408 291864 373414 291876
rect 523034 291864 523040 291876
rect 523092 291864 523098 291916
rect 373258 291796 373264 291848
rect 373316 291836 373322 291848
rect 523126 291836 523132 291848
rect 373316 291808 523132 291836
rect 373316 291796 373322 291808
rect 523126 291796 523132 291808
rect 523184 291796 523190 291848
rect 376202 291728 376208 291780
rect 376260 291768 376266 291780
rect 515030 291768 515036 291780
rect 376260 291740 515036 291768
rect 376260 291728 376266 291740
rect 515030 291728 515036 291740
rect 515088 291728 515094 291780
rect 466914 291660 466920 291712
rect 466972 291700 466978 291712
rect 569218 291700 569224 291712
rect 466972 291672 569224 291700
rect 466972 291660 466978 291672
rect 569218 291660 569224 291672
rect 569276 291660 569282 291712
rect 399478 291592 399484 291644
rect 399536 291632 399542 291644
rect 486142 291632 486148 291644
rect 399536 291604 486148 291632
rect 399536 291592 399542 291604
rect 486142 291592 486148 291604
rect 486200 291592 486206 291644
rect 477862 290436 477868 290488
rect 477920 290476 477926 290488
rect 551278 290476 551284 290488
rect 477920 290448 551284 290476
rect 477920 290436 477926 290448
rect 551278 290436 551284 290448
rect 551336 290436 551342 290488
rect 439682 289620 439688 289672
rect 439740 289660 439746 289672
rect 446398 289660 446404 289672
rect 439740 289632 446404 289660
rect 439740 289620 439746 289632
rect 446398 289620 446404 289632
rect 446456 289620 446462 289672
rect 477586 289620 477592 289672
rect 477644 289660 477650 289672
rect 570598 289660 570604 289672
rect 477644 289632 570604 289660
rect 477644 289620 477650 289632
rect 570598 289620 570604 289632
rect 570656 289620 570662 289672
rect 404998 289552 405004 289604
rect 405056 289592 405062 289604
rect 516410 289592 516416 289604
rect 405056 289564 516416 289592
rect 405056 289552 405062 289564
rect 516410 289552 516416 289564
rect 516468 289552 516474 289604
rect 368106 289484 368112 289536
rect 368164 289524 368170 289536
rect 507118 289524 507124 289536
rect 368164 289496 507124 289524
rect 368164 289484 368170 289496
rect 507118 289484 507124 289496
rect 507176 289484 507182 289536
rect 368198 289416 368204 289468
rect 368256 289456 368262 289468
rect 507302 289456 507308 289468
rect 368256 289428 507308 289456
rect 368256 289416 368262 289428
rect 507302 289416 507308 289428
rect 507360 289416 507366 289468
rect 367738 289348 367744 289400
rect 367796 289388 367802 289400
rect 507210 289388 507216 289400
rect 367796 289360 507216 289388
rect 367796 289348 367802 289360
rect 507210 289348 507216 289360
rect 507268 289348 507274 289400
rect 370958 289280 370964 289332
rect 371016 289320 371022 289332
rect 521654 289320 521660 289332
rect 371016 289292 521660 289320
rect 371016 289280 371022 289292
rect 521654 289280 521660 289292
rect 521712 289280 521718 289332
rect 368014 289212 368020 289264
rect 368072 289252 368078 289264
rect 521838 289252 521844 289264
rect 368072 289224 521844 289252
rect 368072 289212 368078 289224
rect 521838 289212 521844 289224
rect 521896 289212 521902 289264
rect 367922 289144 367928 289196
rect 367980 289184 367986 289196
rect 522022 289184 522028 289196
rect 367980 289156 522028 289184
rect 367980 289144 367986 289156
rect 522022 289144 522028 289156
rect 522080 289144 522086 289196
rect 367830 289076 367836 289128
rect 367888 289116 367894 289128
rect 521930 289116 521936 289128
rect 367888 289088 521936 289116
rect 367888 289076 367894 289088
rect 521930 289076 521936 289088
rect 521988 289076 521994 289128
rect 465718 288396 465724 288448
rect 465776 288436 465782 288448
rect 471238 288436 471244 288448
rect 465776 288408 471244 288436
rect 465776 288396 465782 288408
rect 471238 288396 471244 288408
rect 471296 288396 471302 288448
rect 476758 288396 476764 288448
rect 476816 288436 476822 288448
rect 482278 288436 482284 288448
rect 476816 288408 482284 288436
rect 476816 288396 476822 288408
rect 482278 288396 482284 288408
rect 482336 288396 482342 288448
rect 445018 288328 445024 288380
rect 445076 288368 445082 288380
rect 447778 288368 447784 288380
rect 445076 288340 447784 288368
rect 445076 288328 445082 288340
rect 447778 288328 447784 288340
rect 447836 288328 447842 288380
rect 487246 287648 487252 287700
rect 487304 287688 487310 287700
rect 531314 287688 531320 287700
rect 487304 287660 531320 287688
rect 487304 287648 487310 287660
rect 531314 287648 531320 287660
rect 531372 287648 531378 287700
rect 453850 284996 453856 285048
rect 453908 285036 453914 285048
rect 489178 285036 489184 285048
rect 453908 285008 489184 285036
rect 453908 284996 453914 285008
rect 489178 284996 489184 285008
rect 489236 284996 489242 285048
rect 376018 284928 376024 284980
rect 376076 284968 376082 284980
rect 476574 284968 476580 284980
rect 376076 284940 476580 284968
rect 376076 284928 376082 284940
rect 476574 284928 476580 284940
rect 476632 284928 476638 284980
rect 498378 284928 498384 284980
rect 498436 284968 498442 284980
rect 539870 284968 539876 284980
rect 498436 284940 539876 284968
rect 498436 284928 498442 284940
rect 539870 284928 539876 284940
rect 539928 284928 539934 284980
rect 452470 283568 452476 283620
rect 452528 283608 452534 283620
rect 494514 283608 494520 283620
rect 452528 283580 494520 283608
rect 452528 283568 452534 283580
rect 494514 283568 494520 283580
rect 494572 283568 494578 283620
rect 361758 282820 361764 282872
rect 361816 282860 361822 282872
rect 436830 282860 436836 282872
rect 361816 282832 436836 282860
rect 361816 282820 361822 282832
rect 436830 282820 436836 282832
rect 436888 282820 436894 282872
rect 455046 282208 455052 282260
rect 455104 282248 455110 282260
rect 493318 282248 493324 282260
rect 455104 282220 493324 282248
rect 455104 282208 455110 282220
rect 493318 282208 493324 282220
rect 493376 282208 493382 282260
rect 466822 282140 466828 282192
rect 466880 282180 466886 282192
rect 554038 282180 554044 282192
rect 466880 282152 554044 282180
rect 466880 282140 466886 282152
rect 554038 282140 554044 282152
rect 554096 282140 554102 282192
rect 457622 280780 457628 280832
rect 457680 280820 457686 280832
rect 492858 280820 492864 280832
rect 457680 280792 492864 280820
rect 457680 280780 457686 280792
rect 492858 280780 492864 280792
rect 492916 280780 492922 280832
rect 502426 280780 502432 280832
rect 502484 280820 502490 280832
rect 539042 280820 539048 280832
rect 502484 280792 539048 280820
rect 502484 280780 502490 280792
rect 539042 280780 539048 280792
rect 539100 280780 539106 280832
rect 459278 279488 459284 279540
rect 459336 279528 459342 279540
rect 492214 279528 492220 279540
rect 459336 279500 492220 279528
rect 459336 279488 459342 279500
rect 492214 279488 492220 279500
rect 492272 279488 492278 279540
rect 453942 279420 453948 279472
rect 454000 279460 454006 279472
rect 490558 279460 490564 279472
rect 454000 279432 490564 279460
rect 454000 279420 454006 279432
rect 490558 279420 490564 279432
rect 490616 279420 490622 279472
rect 500218 279420 500224 279472
rect 500276 279460 500282 279472
rect 540146 279460 540152 279472
rect 500276 279432 540152 279460
rect 500276 279420 500282 279432
rect 540146 279420 540152 279432
rect 540204 279420 540210 279472
rect 460474 277992 460480 278044
rect 460532 278032 460538 278044
rect 494698 278032 494704 278044
rect 460532 278004 494704 278032
rect 460532 277992 460538 278004
rect 494698 277992 494704 278004
rect 494756 277992 494762 278044
rect 499942 277992 499948 278044
rect 500000 278032 500006 278044
rect 541434 278032 541440 278044
rect 500000 278004 541440 278032
rect 500000 277992 500006 278004
rect 541434 277992 541440 278004
rect 541492 277992 541498 278044
rect 454862 276632 454868 276684
rect 454920 276672 454926 276684
rect 488994 276672 489000 276684
rect 454920 276644 489000 276672
rect 454920 276632 454926 276644
rect 488994 276632 489000 276644
rect 489052 276632 489058 276684
rect 499758 276632 499764 276684
rect 499816 276672 499822 276684
rect 539962 276672 539968 276684
rect 499816 276644 539968 276672
rect 499816 276632 499822 276644
rect 539962 276632 539968 276644
rect 540020 276632 540026 276684
rect 459462 275340 459468 275392
rect 459520 275380 459526 275392
rect 492766 275380 492772 275392
rect 459520 275352 492772 275380
rect 459520 275340 459526 275352
rect 492766 275340 492772 275352
rect 492824 275340 492830 275392
rect 452286 275272 452292 275324
rect 452344 275312 452350 275324
rect 490006 275312 490012 275324
rect 452344 275284 490012 275312
rect 452344 275272 452350 275284
rect 490006 275272 490012 275284
rect 490064 275272 490070 275324
rect 498838 275272 498844 275324
rect 498896 275312 498902 275324
rect 541250 275312 541256 275324
rect 498896 275284 541256 275312
rect 498896 275272 498902 275284
rect 541250 275272 541256 275284
rect 541308 275272 541314 275324
rect 460566 274048 460572 274100
rect 460624 274088 460630 274100
rect 465718 274088 465724 274100
rect 460624 274060 465724 274088
rect 460624 274048 460630 274060
rect 465718 274048 465724 274060
rect 465776 274048 465782 274100
rect 455138 273980 455144 274032
rect 455196 274020 455202 274032
rect 491938 274020 491944 274032
rect 455196 273992 491944 274020
rect 455196 273980 455202 273992
rect 491938 273980 491944 273992
rect 491996 273980 492002 274032
rect 498562 273980 498568 274032
rect 498620 274020 498626 274032
rect 541342 274020 541348 274032
rect 498620 273992 541348 274020
rect 498620 273980 498626 273992
rect 541342 273980 541348 273992
rect 541400 273980 541406 274032
rect 456610 273912 456616 273964
rect 456668 273952 456674 273964
rect 495894 273952 495900 273964
rect 456668 273924 495900 273952
rect 456668 273912 456674 273924
rect 495894 273912 495900 273924
rect 495952 273912 495958 273964
rect 497458 273912 497464 273964
rect 497516 273952 497522 273964
rect 541158 273952 541164 273964
rect 497516 273924 541164 273952
rect 497516 273912 497522 273924
rect 541158 273912 541164 273924
rect 541216 273912 541222 273964
rect 479518 273164 479524 273216
rect 479576 273204 479582 273216
rect 580166 273204 580172 273216
rect 479576 273176 580172 273204
rect 479576 273164 479582 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 457714 272552 457720 272604
rect 457772 272592 457778 272604
rect 491662 272592 491668 272604
rect 457772 272564 491668 272592
rect 457772 272552 457778 272564
rect 491662 272552 491668 272564
rect 491720 272552 491726 272604
rect 457806 272484 457812 272536
rect 457864 272524 457870 272536
rect 494422 272524 494428 272536
rect 457864 272496 494428 272524
rect 457864 272484 457870 272496
rect 494422 272484 494428 272496
rect 494480 272484 494486 272536
rect 501046 272484 501052 272536
rect 501104 272524 501110 272536
rect 540238 272524 540244 272536
rect 501104 272496 540244 272524
rect 501104 272484 501110 272496
rect 540238 272484 540244 272496
rect 540296 272484 540302 272536
rect 361758 271804 361764 271856
rect 361816 271844 361822 271856
rect 431218 271844 431224 271856
rect 361816 271816 431224 271844
rect 361816 271804 361822 271816
rect 431218 271804 431224 271816
rect 431276 271804 431282 271856
rect 459370 271260 459376 271312
rect 459428 271300 459434 271312
rect 493134 271300 493140 271312
rect 459428 271272 493140 271300
rect 459428 271260 459434 271272
rect 493134 271260 493140 271272
rect 493192 271260 493198 271312
rect 454954 271192 454960 271244
rect 455012 271232 455018 271244
rect 488626 271232 488632 271244
rect 455012 271204 488632 271232
rect 455012 271192 455018 271204
rect 488626 271192 488632 271204
rect 488684 271192 488690 271244
rect 498286 271192 498292 271244
rect 498344 271232 498350 271244
rect 540054 271232 540060 271244
rect 498344 271204 540060 271232
rect 498344 271192 498350 271204
rect 540054 271192 540060 271204
rect 540112 271192 540118 271244
rect 453206 271124 453212 271176
rect 453264 271164 453270 271176
rect 488902 271164 488908 271176
rect 453264 271136 488908 271164
rect 453264 271124 453270 271136
rect 488902 271124 488908 271136
rect 488960 271124 488966 271176
rect 499666 271124 499672 271176
rect 499724 271164 499730 271176
rect 541526 271164 541532 271176
rect 499724 271136 541532 271164
rect 499724 271124 499730 271136
rect 541526 271124 541532 271136
rect 541584 271124 541590 271176
rect 503806 269968 503812 270020
rect 503864 270008 503870 270020
rect 543734 270008 543740 270020
rect 503864 269980 543740 270008
rect 503864 269968 503870 269980
rect 543734 269968 543740 269980
rect 543792 269968 543798 270020
rect 456702 269900 456708 269952
rect 456760 269940 456766 269952
rect 488074 269940 488080 269952
rect 456760 269912 488080 269940
rect 456760 269900 456766 269912
rect 488074 269900 488080 269912
rect 488132 269900 488138 269952
rect 497182 269900 497188 269952
rect 497240 269940 497246 269952
rect 542814 269940 542820 269952
rect 497240 269912 542820 269940
rect 497240 269900 497246 269912
rect 542814 269900 542820 269912
rect 542872 269900 542878 269952
rect 467926 269832 467932 269884
rect 467984 269872 467990 269884
rect 580258 269872 580264 269884
rect 467984 269844 580264 269872
rect 467984 269832 467990 269844
rect 580258 269832 580264 269844
rect 580316 269832 580322 269884
rect 359550 269764 359556 269816
rect 359608 269804 359614 269816
rect 512730 269804 512736 269816
rect 359608 269776 512736 269804
rect 359608 269764 359614 269776
rect 512730 269764 512736 269776
rect 512788 269764 512794 269816
rect 481082 269288 481088 269340
rect 481140 269328 481146 269340
rect 484762 269328 484768 269340
rect 481140 269300 484768 269328
rect 481140 269288 481146 269300
rect 484762 269288 484768 269300
rect 484820 269288 484826 269340
rect 445662 268540 445668 268592
rect 445720 268580 445726 268592
rect 476758 268580 476764 268592
rect 445720 268552 476764 268580
rect 445720 268540 445726 268552
rect 476758 268540 476764 268552
rect 476816 268540 476822 268592
rect 447778 268472 447784 268524
rect 447836 268512 447842 268524
rect 481082 268512 481088 268524
rect 447836 268484 481088 268512
rect 447836 268472 447842 268484
rect 481082 268472 481088 268484
rect 481140 268472 481146 268524
rect 452378 268404 452384 268456
rect 452436 268444 452442 268456
rect 490282 268444 490288 268456
rect 452436 268416 490288 268444
rect 452436 268404 452442 268416
rect 490282 268404 490288 268416
rect 490340 268404 490346 268456
rect 496906 268404 496912 268456
rect 496964 268444 496970 268456
rect 542630 268444 542636 268456
rect 496964 268416 542636 268444
rect 496964 268404 496970 268416
rect 542630 268404 542636 268416
rect 542688 268404 542694 268456
rect 466546 268336 466552 268388
rect 466604 268376 466610 268388
rect 555418 268376 555424 268388
rect 466604 268348 555424 268376
rect 466604 268336 466610 268348
rect 555418 268336 555424 268348
rect 555476 268336 555482 268388
rect 435450 266976 435456 267028
rect 435508 267016 435514 267028
rect 460566 267016 460572 267028
rect 435508 266988 460572 267016
rect 435508 266976 435514 266988
rect 460566 266976 460572 266988
rect 460624 266976 460630 267028
rect 3510 266364 3516 266416
rect 3568 266404 3574 266416
rect 4890 266404 4896 266416
rect 3568 266376 4896 266404
rect 3568 266364 3574 266376
rect 4890 266364 4896 266376
rect 4948 266364 4954 266416
rect 447962 265616 447968 265668
rect 448020 265656 448026 265668
rect 457898 265656 457904 265668
rect 448020 265628 457904 265656
rect 448020 265616 448026 265628
rect 457898 265616 457904 265628
rect 457956 265616 457962 265668
rect 420914 264256 420920 264308
rect 420972 264296 420978 264308
rect 439682 264296 439688 264308
rect 420972 264268 439688 264296
rect 420972 264256 420978 264268
rect 439682 264256 439688 264268
rect 439740 264256 439746 264308
rect 422938 264188 422944 264240
rect 422996 264228 423002 264240
rect 445662 264228 445668 264240
rect 422996 264200 445668 264228
rect 422996 264188 423002 264200
rect 445662 264188 445668 264200
rect 445720 264188 445726 264240
rect 449710 263508 449716 263560
rect 449768 263548 449774 263560
rect 456794 263548 456800 263560
rect 449768 263520 456800 263548
rect 449768 263508 449774 263520
rect 456794 263508 456800 263520
rect 456852 263508 456858 263560
rect 431218 262828 431224 262880
rect 431276 262868 431282 262880
rect 445018 262868 445024 262880
rect 431276 262840 445024 262868
rect 431276 262828 431282 262840
rect 445018 262828 445024 262840
rect 445076 262828 445082 262880
rect 411898 261468 411904 261520
rect 411956 261508 411962 261520
rect 420914 261508 420920 261520
rect 411956 261480 420920 261508
rect 411956 261468 411962 261480
rect 420914 261468 420920 261480
rect 420972 261468 420978 261520
rect 361758 260788 361764 260840
rect 361816 260828 361822 260840
rect 440970 260828 440976 260840
rect 361816 260800 440976 260828
rect 361816 260788 361822 260800
rect 440970 260788 440976 260800
rect 441028 260788 441034 260840
rect 401410 255960 401416 256012
rect 401468 256000 401474 256012
rect 411898 256000 411904 256012
rect 401468 255972 411904 256000
rect 401468 255960 401474 255972
rect 411898 255960 411904 255972
rect 411956 255960 411962 256012
rect 428458 253920 428464 253972
rect 428516 253960 428522 253972
rect 431218 253960 431224 253972
rect 428516 253932 431224 253960
rect 428516 253920 428522 253932
rect 431218 253920 431224 253932
rect 431276 253920 431282 253972
rect 361758 249704 361764 249756
rect 361816 249744 361822 249756
rect 435358 249744 435364 249756
rect 361816 249716 435364 249744
rect 361816 249704 361822 249716
rect 435358 249704 435364 249716
rect 435416 249704 435422 249756
rect 449802 249704 449808 249756
rect 449860 249744 449866 249756
rect 449986 249744 449992 249756
rect 449860 249716 449992 249744
rect 449860 249704 449866 249716
rect 449986 249704 449992 249716
rect 450044 249704 450050 249756
rect 449986 248412 449992 248464
rect 450044 248452 450050 248464
rect 456794 248452 456800 248464
rect 450044 248424 456800 248452
rect 450044 248412 450050 248424
rect 456794 248412 456800 248424
rect 456852 248412 456858 248464
rect 571978 245556 571984 245608
rect 572036 245596 572042 245608
rect 580166 245596 580172 245608
rect 572036 245568 580172 245596
rect 572036 245556 572042 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 398466 243176 398472 243228
rect 398524 243216 398530 243228
rect 401410 243216 401416 243228
rect 398524 243188 401416 243216
rect 398524 243176 398530 243188
rect 401410 243176 401416 243188
rect 401468 243176 401474 243228
rect 3878 241408 3884 241460
rect 3936 241448 3942 241460
rect 4982 241448 4988 241460
rect 3936 241420 4988 241448
rect 3936 241408 3942 241420
rect 4982 241408 4988 241420
rect 5040 241408 5046 241460
rect 422294 240796 422300 240848
rect 422352 240836 422358 240848
rect 428458 240836 428464 240848
rect 422352 240808 428464 240836
rect 422352 240796 422358 240808
rect 428458 240796 428464 240808
rect 428516 240796 428522 240848
rect 435358 240728 435364 240780
rect 435416 240768 435422 240780
rect 447778 240768 447784 240780
rect 435416 240740 447784 240768
rect 435416 240728 435422 240740
rect 447778 240728 447784 240740
rect 447836 240728 447842 240780
rect 361758 238688 361764 238740
rect 361816 238728 361822 238740
rect 439590 238728 439596 238740
rect 361816 238700 439596 238728
rect 361816 238688 361822 238700
rect 439590 238688 439596 238700
rect 439648 238688 439654 238740
rect 414658 238008 414664 238060
rect 414716 238048 414722 238060
rect 422294 238048 422300 238060
rect 414716 238020 422300 238048
rect 414716 238008 414722 238020
rect 422294 238008 422300 238020
rect 422352 238008 422358 238060
rect 386414 235220 386420 235272
rect 386472 235260 386478 235272
rect 398466 235260 398472 235272
rect 386472 235232 398472 235260
rect 386472 235220 386478 235232
rect 398466 235220 398472 235232
rect 398524 235220 398530 235272
rect 570598 233180 570604 233232
rect 570656 233220 570662 233232
rect 579982 233220 579988 233232
rect 570656 233192 579988 233220
rect 570656 233180 570662 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 427078 232500 427084 232552
rect 427136 232540 427142 232552
rect 435358 232540 435364 232552
rect 427136 232512 435364 232540
rect 427136 232500 427142 232512
rect 435358 232500 435364 232512
rect 435416 232500 435422 232552
rect 384666 232024 384672 232076
rect 384724 232064 384730 232076
rect 386414 232064 386420 232076
rect 384724 232036 386420 232064
rect 384724 232024 384730 232036
rect 386414 232024 386420 232036
rect 386472 232024 386478 232076
rect 361758 227672 361764 227724
rect 361816 227712 361822 227724
rect 442258 227712 442264 227724
rect 361816 227684 442264 227712
rect 361816 227672 361822 227684
rect 442258 227672 442264 227684
rect 442316 227672 442322 227724
rect 455230 222096 455236 222148
rect 455288 222136 455294 222148
rect 456794 222136 456800 222148
rect 455288 222108 456800 222136
rect 455288 222096 455294 222108
rect 456794 222096 456800 222108
rect 456852 222096 456858 222148
rect 394694 221416 394700 221468
rect 394752 221456 394758 221468
rect 414658 221456 414664 221468
rect 394752 221428 414664 221456
rect 394752 221416 394758 221428
rect 414658 221416 414664 221428
rect 414716 221416 414722 221468
rect 428458 221416 428464 221468
rect 428516 221456 428522 221468
rect 435450 221456 435456 221468
rect 428516 221428 435456 221456
rect 428516 221416 428522 221428
rect 435450 221416 435456 221428
rect 435508 221416 435514 221468
rect 559558 219376 559564 219428
rect 559616 219416 559622 219428
rect 580166 219416 580172 219428
rect 559616 219388 580172 219416
rect 559616 219376 559622 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 391934 218016 391940 218068
rect 391992 218056 391998 218068
rect 394694 218056 394700 218068
rect 391992 218028 394700 218056
rect 391992 218016 391998 218028
rect 394694 218016 394700 218028
rect 394752 218016 394758 218068
rect 361574 216316 361580 216368
rect 361632 216356 361638 216368
rect 363598 216356 363604 216368
rect 361632 216328 363604 216356
rect 361632 216316 361638 216328
rect 363598 216316 363604 216328
rect 363656 216316 363662 216368
rect 387610 215296 387616 215348
rect 387668 215336 387674 215348
rect 391934 215336 391940 215348
rect 387668 215308 391940 215336
rect 387668 215296 387674 215308
rect 391934 215296 391940 215308
rect 391992 215296 391998 215348
rect 3786 214752 3792 214804
rect 3844 214792 3850 214804
rect 5074 214792 5080 214804
rect 3844 214764 5080 214792
rect 3844 214752 3850 214764
rect 5074 214752 5080 214764
rect 5132 214752 5138 214804
rect 411898 213188 411904 213240
rect 411956 213228 411962 213240
rect 427078 213228 427084 213240
rect 411956 213200 427084 213228
rect 411956 213188 411962 213200
rect 427078 213188 427084 213200
rect 427136 213188 427142 213240
rect 379330 212984 379336 213036
rect 379388 213024 379394 213036
rect 384666 213024 384672 213036
rect 379388 212996 384672 213024
rect 379388 212984 379394 212996
rect 384666 212984 384672 212996
rect 384724 212984 384730 213036
rect 448330 207612 448336 207664
rect 448388 207652 448394 207664
rect 454034 207652 454040 207664
rect 448388 207624 454040 207652
rect 448388 207612 448394 207624
rect 454034 207612 454040 207624
rect 454092 207652 454098 207664
rect 456886 207652 456892 207664
rect 454092 207624 456892 207652
rect 454092 207612 454098 207624
rect 456886 207612 456892 207624
rect 456944 207612 456950 207664
rect 418062 207272 418068 207324
rect 418120 207312 418126 207324
rect 422938 207312 422944 207324
rect 418120 207284 422944 207312
rect 418120 207272 418126 207284
rect 422938 207272 422944 207284
rect 422996 207272 423002 207324
rect 404078 205640 404084 205692
rect 404136 205680 404142 205692
rect 411898 205680 411904 205692
rect 404136 205652 411904 205680
rect 404136 205640 404142 205652
rect 411898 205640 411904 205652
rect 411956 205640 411962 205692
rect 361758 205572 361764 205624
rect 361816 205612 361822 205624
rect 439498 205612 439504 205624
rect 361816 205584 439504 205612
rect 361816 205572 361822 205584
rect 439498 205572 439504 205584
rect 439556 205572 439562 205624
rect 362310 204892 362316 204944
rect 362368 204932 362374 204944
rect 379330 204932 379336 204944
rect 362368 204904 379336 204932
rect 362368 204892 362374 204904
rect 379330 204892 379336 204904
rect 379388 204892 379394 204944
rect 3970 204212 3976 204264
rect 4028 204252 4034 204264
rect 5166 204252 5172 204264
rect 4028 204224 5172 204252
rect 4028 204212 4034 204224
rect 5166 204212 5172 204224
rect 5224 204212 5230 204264
rect 414658 201016 414664 201068
rect 414716 201056 414722 201068
rect 418062 201056 418068 201068
rect 414716 201028 418068 201056
rect 414716 201016 414722 201028
rect 418062 201016 418068 201028
rect 418120 201016 418126 201068
rect 458726 200744 458732 200796
rect 458784 200784 458790 200796
rect 481634 200784 481640 200796
rect 458784 200756 481640 200784
rect 458784 200744 458790 200756
rect 481634 200744 481640 200756
rect 481692 200744 481698 200796
rect 379330 199384 379336 199436
rect 379388 199424 379394 199436
rect 387610 199424 387616 199436
rect 379388 199396 387616 199424
rect 379388 199384 379394 199396
rect 387610 199384 387616 199396
rect 387668 199384 387674 199436
rect 456794 197956 456800 198008
rect 456852 197996 456858 198008
rect 485774 197996 485780 198008
rect 456852 197968 485780 197996
rect 456852 197956 456858 197968
rect 485774 197956 485780 197968
rect 485832 197956 485838 198008
rect 361666 194488 361672 194540
rect 361724 194528 361730 194540
rect 443638 194528 443644 194540
rect 361724 194500 443644 194528
rect 361724 194488 361730 194500
rect 443638 194488 443644 194500
rect 443696 194488 443702 194540
rect 551278 193128 551284 193180
rect 551336 193168 551342 193180
rect 580166 193168 580172 193180
rect 551336 193140 580172 193168
rect 551336 193128 551342 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 372614 189728 372620 189780
rect 372672 189768 372678 189780
rect 379330 189768 379336 189780
rect 372672 189740 379336 189768
rect 372672 189728 372678 189740
rect 379330 189728 379336 189740
rect 379388 189728 379394 189780
rect 361206 186940 361212 186992
rect 361264 186980 361270 186992
rect 372614 186980 372620 186992
rect 361264 186952 372620 186980
rect 361264 186940 361270 186952
rect 372614 186940 372620 186952
rect 372672 186940 372678 186992
rect 361666 183472 361672 183524
rect 361724 183512 361730 183524
rect 436738 183512 436744 183524
rect 361724 183484 436744 183512
rect 361724 183472 361730 183484
rect 436738 183472 436744 183484
rect 436796 183472 436802 183524
rect 555418 179324 555424 179376
rect 555476 179364 555482 179376
rect 580166 179364 580172 179376
rect 555476 179336 580172 179364
rect 555476 179324 555482 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 425054 178032 425060 178084
rect 425112 178072 425118 178084
rect 428458 178072 428464 178084
rect 425112 178044 428464 178072
rect 425112 178032 425118 178044
rect 428458 178032 428464 178044
rect 428516 178032 428522 178084
rect 399570 176808 399576 176860
rect 399628 176848 399634 176860
rect 404078 176848 404084 176860
rect 399628 176820 404084 176848
rect 399628 176808 399634 176820
rect 404078 176808 404084 176820
rect 404136 176808 404142 176860
rect 411254 171844 411260 171896
rect 411312 171884 411318 171896
rect 425054 171884 425060 171896
rect 411312 171856 425060 171884
rect 411312 171844 411318 171856
rect 425054 171844 425060 171856
rect 425112 171844 425118 171896
rect 361758 171776 361764 171828
rect 361816 171816 361822 171828
rect 440878 171816 440884 171828
rect 361816 171788 440884 171816
rect 361816 171776 361822 171788
rect 440878 171776 440884 171788
rect 440936 171816 440942 171828
rect 524414 171816 524420 171828
rect 440936 171788 524420 171816
rect 440936 171776 440942 171788
rect 524414 171776 524420 171788
rect 524472 171776 524478 171828
rect 404078 168376 404084 168428
rect 404136 168416 404142 168428
rect 411254 168416 411260 168428
rect 404136 168388 411260 168416
rect 404136 168376 404142 168388
rect 411254 168376 411260 168388
rect 411312 168376 411318 168428
rect 537478 166948 537484 167000
rect 537536 166988 537542 167000
rect 580166 166988 580172 167000
rect 537536 166960 580172 166988
rect 537536 166948 537542 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 411898 164840 411904 164892
rect 411956 164880 411962 164892
rect 454034 164880 454040 164892
rect 411956 164852 454040 164880
rect 411956 164840 411962 164852
rect 454034 164840 454040 164852
rect 454092 164840 454098 164892
rect 402974 163480 402980 163532
rect 403032 163520 403038 163532
rect 414658 163520 414664 163532
rect 403032 163492 414664 163520
rect 403032 163480 403038 163492
rect 414658 163480 414664 163492
rect 414716 163480 414722 163532
rect 448422 163480 448428 163532
rect 448480 163520 448486 163532
rect 528554 163520 528560 163532
rect 448480 163492 528560 163520
rect 448480 163480 448486 163492
rect 528554 163480 528560 163492
rect 528612 163480 528618 163532
rect 445202 163072 445208 163124
rect 445260 163112 445266 163124
rect 449986 163112 449992 163124
rect 445260 163084 449992 163112
rect 445260 163072 445266 163084
rect 449986 163072 449992 163084
rect 450044 163072 450050 163124
rect 418706 162188 418712 162240
rect 418764 162228 418770 162240
rect 458082 162228 458088 162240
rect 418764 162200 458088 162228
rect 418764 162188 418770 162200
rect 458082 162188 458088 162200
rect 458140 162228 458146 162240
rect 458140 162200 460934 162228
rect 458140 162188 458146 162200
rect 414750 162120 414756 162172
rect 414808 162160 414814 162172
rect 456794 162160 456800 162172
rect 414808 162132 456800 162160
rect 414808 162120 414814 162132
rect 456794 162120 456800 162132
rect 456852 162120 456858 162172
rect 460906 162160 460934 162200
rect 489914 162160 489920 162172
rect 460906 162132 489920 162160
rect 489914 162120 489920 162132
rect 489972 162120 489978 162172
rect 426158 161780 426164 161832
rect 426216 161820 426222 161832
rect 496814 161820 496820 161832
rect 426216 161792 496820 161820
rect 426216 161780 426222 161792
rect 496814 161780 496820 161792
rect 496872 161780 496878 161832
rect 428642 161712 428648 161764
rect 428700 161752 428706 161764
rect 500954 161752 500960 161764
rect 428700 161724 500960 161752
rect 428700 161712 428706 161724
rect 500954 161712 500960 161724
rect 501012 161712 501018 161764
rect 421374 161644 421380 161696
rect 421432 161684 421438 161696
rect 494054 161684 494060 161696
rect 421432 161656 494060 161684
rect 421432 161644 421438 161656
rect 494054 161644 494060 161656
rect 494112 161644 494118 161696
rect 431862 161576 431868 161628
rect 431920 161616 431926 161628
rect 505094 161616 505100 161628
rect 431920 161588 505100 161616
rect 431920 161576 431926 161588
rect 505094 161576 505100 161588
rect 505152 161576 505158 161628
rect 438762 161508 438768 161560
rect 438820 161548 438826 161560
rect 513374 161548 513380 161560
rect 438820 161520 513380 161548
rect 438820 161508 438826 161520
rect 513374 161508 513380 161520
rect 513432 161508 513438 161560
rect 362402 161440 362408 161492
rect 362460 161480 362466 161492
rect 441614 161480 441620 161492
rect 362460 161452 441620 161480
rect 362460 161440 362466 161452
rect 441614 161440 441620 161452
rect 441672 161480 441678 161492
rect 442902 161480 442908 161492
rect 441672 161452 442908 161480
rect 441672 161440 441678 161452
rect 442902 161440 442908 161452
rect 442960 161480 442966 161492
rect 517514 161480 517520 161492
rect 442960 161452 517520 161480
rect 442960 161440 442966 161452
rect 517514 161440 517520 161452
rect 517572 161440 517578 161492
rect 361758 161372 361764 161424
rect 361816 161412 361822 161424
rect 444282 161412 444288 161424
rect 361816 161384 444288 161412
rect 361816 161372 361822 161384
rect 444282 161372 444288 161384
rect 444340 161372 444346 161424
rect 391934 160692 391940 160744
rect 391992 160732 391998 160744
rect 402974 160732 402980 160744
rect 391992 160704 402980 160732
rect 391992 160692 391998 160704
rect 402974 160692 402980 160704
rect 403032 160692 403038 160744
rect 444282 160692 444288 160744
rect 444340 160732 444346 160744
rect 521654 160732 521660 160744
rect 444340 160704 521660 160732
rect 444340 160692 444346 160704
rect 521654 160692 521660 160704
rect 521712 160692 521718 160744
rect 406838 160556 406844 160608
rect 406896 160596 406902 160608
rect 414750 160596 414756 160608
rect 406896 160568 414756 160596
rect 406896 160556 406902 160568
rect 414750 160556 414756 160568
rect 414808 160556 414814 160608
rect 404170 160488 404176 160540
rect 404228 160528 404234 160540
rect 411622 160528 411628 160540
rect 404228 160500 411628 160528
rect 404228 160488 404234 160500
rect 411622 160488 411628 160500
rect 411680 160488 411686 160540
rect 410518 160420 410524 160472
rect 410576 160460 410582 160472
rect 418154 160460 418160 160472
rect 410576 160432 418160 160460
rect 410576 160420 410582 160432
rect 418154 160420 418160 160432
rect 418212 160420 418218 160472
rect 410610 160352 410616 160404
rect 410668 160392 410674 160404
rect 425146 160392 425152 160404
rect 410668 160364 425152 160392
rect 410668 160352 410674 160364
rect 425146 160352 425152 160364
rect 425204 160392 425210 160404
rect 426158 160392 426164 160404
rect 425204 160364 426164 160392
rect 425204 160352 425210 160364
rect 426158 160352 426164 160364
rect 426216 160352 426222 160404
rect 407850 160284 407856 160336
rect 407908 160324 407914 160336
rect 407908 160296 411576 160324
rect 407908 160284 407914 160296
rect 407758 160216 407764 160268
rect 407816 160256 407822 160268
rect 411438 160256 411444 160268
rect 407816 160228 411444 160256
rect 407816 160216 407822 160228
rect 411438 160216 411444 160228
rect 411496 160216 411502 160268
rect 411548 160256 411576 160296
rect 411622 160284 411628 160336
rect 411680 160324 411686 160336
rect 421374 160324 421380 160336
rect 411680 160296 421380 160324
rect 411680 160284 411686 160296
rect 421374 160284 421380 160296
rect 421432 160284 421438 160336
rect 427998 160256 428004 160268
rect 411548 160228 428004 160256
rect 427998 160216 428004 160228
rect 428056 160216 428062 160268
rect 409322 160148 409328 160200
rect 409380 160188 409386 160200
rect 431310 160188 431316 160200
rect 409380 160160 431316 160188
rect 409380 160148 409386 160160
rect 431310 160148 431316 160160
rect 431368 160148 431374 160200
rect 435266 160148 435272 160200
rect 435324 160188 435330 160200
rect 436002 160188 436008 160200
rect 435324 160160 436008 160188
rect 435324 160148 435330 160160
rect 436002 160148 436008 160160
rect 436060 160188 436066 160200
rect 451182 160188 451188 160200
rect 436060 160160 451188 160188
rect 436060 160148 436066 160160
rect 451182 160148 451188 160160
rect 451240 160148 451246 160200
rect 410702 160080 410708 160132
rect 410760 160120 410766 160132
rect 438256 160120 438262 160132
rect 410760 160092 438262 160120
rect 410760 160080 410766 160092
rect 438256 160080 438262 160092
rect 438314 160080 438320 160132
rect 444880 160080 444886 160132
rect 444938 160120 444944 160132
rect 445202 160120 445208 160132
rect 444938 160092 445208 160120
rect 444938 160080 444944 160092
rect 445202 160080 445208 160092
rect 445260 160120 445266 160132
rect 483658 160120 483664 160132
rect 445260 160092 483664 160120
rect 445260 160080 445266 160092
rect 483658 160080 483664 160092
rect 483716 160080 483722 160132
rect 434806 159372 434812 159384
rect 431926 159344 434812 159372
rect 363598 158720 363604 158772
rect 363656 158760 363662 158772
rect 431926 158760 431954 159344
rect 434806 159332 434812 159344
rect 434864 159332 434870 159384
rect 363656 158732 431954 158760
rect 363656 158720 363662 158732
rect 451734 158380 451740 158432
rect 451792 158420 451798 158432
rect 456702 158420 456708 158432
rect 451792 158392 456708 158420
rect 451792 158380 451798 158392
rect 456702 158380 456708 158392
rect 456760 158380 456766 158432
rect 452562 156884 452568 156936
rect 452620 156924 452626 156936
rect 456610 156924 456616 156936
rect 452620 156896 456616 156924
rect 452620 156884 452626 156896
rect 456610 156884 456616 156896
rect 456668 156884 456674 156936
rect 382090 155184 382096 155236
rect 382148 155224 382154 155236
rect 391934 155224 391940 155236
rect 382148 155196 391940 155224
rect 382148 155184 382154 155196
rect 391934 155184 391940 155196
rect 391992 155184 391998 155236
rect 547138 153144 547144 153196
rect 547196 153184 547202 153196
rect 580166 153184 580172 153196
rect 547196 153156 580172 153184
rect 547196 153144 547202 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 452102 152940 452108 152992
rect 452160 152980 452166 152992
rect 460474 152980 460480 152992
rect 452160 152952 460480 152980
rect 452160 152940 452166 152952
rect 460474 152940 460480 152952
rect 460532 152940 460538 152992
rect 452562 151444 452568 151496
rect 452620 151484 452626 151496
rect 457806 151484 457812 151496
rect 452620 151456 457812 151484
rect 452620 151444 452626 151456
rect 457806 151444 457812 151456
rect 457864 151444 457870 151496
rect 393958 149064 393964 149116
rect 394016 149104 394022 149116
rect 399570 149104 399576 149116
rect 394016 149076 399576 149104
rect 394016 149064 394022 149076
rect 399570 149064 399576 149076
rect 399628 149064 399634 149116
rect 452562 147364 452568 147416
rect 452620 147404 452626 147416
rect 459462 147404 459468 147416
rect 452620 147376 459468 147404
rect 452620 147364 452626 147376
rect 459462 147364 459468 147376
rect 459520 147364 459526 147416
rect 452562 146140 452568 146192
rect 452620 146180 452626 146192
rect 457530 146180 457536 146192
rect 452620 146152 457536 146180
rect 452620 146140 452626 146152
rect 457530 146140 457536 146152
rect 457588 146140 457594 146192
rect 452562 144644 452568 144696
rect 452620 144684 452626 144696
rect 455046 144684 455052 144696
rect 452620 144656 455052 144684
rect 452620 144644 452626 144656
rect 455046 144644 455052 144656
rect 455104 144644 455110 144696
rect 452562 143284 452568 143336
rect 452620 143324 452626 143336
rect 459370 143324 459376 143336
rect 452620 143296 459376 143324
rect 452620 143284 452626 143296
rect 459370 143284 459376 143296
rect 459428 143284 459434 143336
rect 483658 142876 483664 142928
rect 483716 142916 483722 142928
rect 533982 142916 533988 142928
rect 483716 142888 533988 142916
rect 483716 142876 483722 142888
rect 533982 142876 533988 142888
rect 534040 142876 534046 142928
rect 451182 142808 451188 142860
rect 451240 142848 451246 142860
rect 509602 142848 509608 142860
rect 451240 142820 509608 142848
rect 451240 142808 451246 142820
rect 509602 142808 509608 142820
rect 509660 142808 509666 142860
rect 533982 142128 533988 142180
rect 534040 142168 534046 142180
rect 539778 142168 539784 142180
rect 534040 142140 539784 142168
rect 534040 142128 534046 142140
rect 539778 142128 539784 142140
rect 539836 142128 539842 142180
rect 452562 141924 452568 141976
rect 452620 141964 452626 141976
rect 457622 141964 457628 141976
rect 452620 141936 457628 141964
rect 452620 141924 452626 141936
rect 457622 141924 457628 141936
rect 457680 141924 457686 141976
rect 388346 140768 388352 140820
rect 388404 140808 388410 140820
rect 393958 140808 393964 140820
rect 388404 140780 393964 140808
rect 388404 140768 388410 140780
rect 393958 140768 393964 140780
rect 394016 140768 394022 140820
rect 452102 140632 452108 140684
rect 452160 140672 452166 140684
rect 455138 140672 455144 140684
rect 452160 140644 455144 140672
rect 452160 140632 452166 140644
rect 455138 140632 455144 140644
rect 455196 140632 455202 140684
rect 530670 140088 530676 140140
rect 530728 140128 530734 140140
rect 542538 140128 542544 140140
rect 530728 140100 542544 140128
rect 530728 140088 530734 140100
rect 542538 140088 542544 140100
rect 542596 140088 542602 140140
rect 530578 140020 530584 140072
rect 530636 140060 530642 140072
rect 542446 140060 542452 140072
rect 530636 140032 542452 140060
rect 530636 140020 530642 140032
rect 542446 140020 542452 140032
rect 542504 140020 542510 140072
rect 379330 139408 379336 139460
rect 379388 139448 379394 139460
rect 382090 139448 382096 139460
rect 379388 139420 382096 139448
rect 379388 139408 379394 139420
rect 382090 139408 382096 139420
rect 382148 139408 382154 139460
rect 361758 139340 361764 139392
rect 361816 139380 361822 139392
rect 410702 139380 410708 139392
rect 361816 139352 410708 139380
rect 361816 139340 361822 139352
rect 410702 139340 410708 139352
rect 410760 139340 410766 139392
rect 452562 139340 452568 139392
rect 452620 139380 452626 139392
rect 459278 139380 459284 139392
rect 452620 139352 459284 139380
rect 452620 139340 452626 139352
rect 459278 139340 459284 139352
rect 459336 139340 459342 139392
rect 554038 139340 554044 139392
rect 554096 139380 554102 139392
rect 580166 139380 580172 139392
rect 554096 139352 580172 139380
rect 554096 139340 554102 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 538858 139204 538864 139256
rect 538916 139244 538922 139256
rect 543182 139244 543188 139256
rect 538916 139216 543188 139244
rect 538916 139204 538922 139216
rect 543182 139204 543188 139216
rect 543240 139204 543246 139256
rect 452562 137844 452568 137896
rect 452620 137884 452626 137896
rect 457714 137884 457720 137896
rect 452620 137856 457720 137884
rect 452620 137844 452626 137856
rect 457714 137844 457720 137856
rect 457772 137844 457778 137896
rect 538950 136552 538956 136604
rect 539008 136592 539014 136604
rect 539502 136592 539508 136604
rect 539008 136564 539508 136592
rect 539008 136552 539014 136564
rect 539502 136552 539508 136564
rect 539560 136552 539566 136604
rect 452562 136484 452568 136536
rect 452620 136524 452626 136536
rect 454770 136524 454776 136536
rect 452620 136496 454776 136524
rect 452620 136484 452626 136496
rect 454770 136484 454776 136496
rect 454828 136484 454834 136536
rect 363690 135872 363696 135924
rect 363748 135912 363754 135924
rect 388346 135912 388352 135924
rect 363748 135884 388352 135912
rect 363748 135872 363754 135884
rect 388346 135872 388352 135884
rect 388404 135872 388410 135924
rect 452562 135124 452568 135176
rect 452620 135164 452626 135176
rect 459186 135164 459192 135176
rect 452620 135136 459192 135164
rect 452620 135124 452626 135136
rect 459186 135124 459192 135136
rect 459244 135124 459250 135176
rect 452470 133764 452476 133816
rect 452528 133804 452534 133816
rect 453758 133804 453764 133816
rect 452528 133776 453764 133804
rect 452528 133764 452534 133776
rect 453758 133764 453764 133776
rect 453816 133764 453822 133816
rect 452102 132404 452108 132456
rect 452160 132444 452166 132456
rect 453666 132444 453672 132456
rect 452160 132416 453672 132444
rect 452160 132404 452166 132416
rect 453666 132404 453672 132416
rect 453724 132404 453730 132456
rect 361298 131112 361304 131164
rect 361356 131152 361362 131164
rect 363690 131152 363696 131164
rect 361356 131124 363696 131152
rect 361356 131112 361362 131124
rect 363690 131112 363696 131124
rect 363748 131112 363754 131164
rect 452562 131044 452568 131096
rect 452620 131084 452626 131096
rect 453942 131084 453948 131096
rect 452620 131056 453948 131084
rect 452620 131044 452626 131056
rect 453942 131044 453948 131056
rect 454000 131044 454006 131096
rect 373626 129004 373632 129056
rect 373684 129044 373690 129056
rect 379330 129044 379336 129056
rect 373684 129016 379336 129044
rect 373684 129004 373690 129016
rect 379330 129004 379336 129016
rect 379388 129004 379394 129056
rect 361574 128188 361580 128240
rect 361632 128228 361638 128240
rect 363598 128228 363604 128240
rect 361632 128200 363604 128228
rect 361632 128188 361638 128200
rect 363598 128188 363604 128200
rect 363656 128188 363662 128240
rect 452194 126896 452200 126948
rect 452252 126936 452258 126948
rect 453206 126936 453212 126948
rect 452252 126908 453212 126936
rect 452252 126896 452258 126908
rect 453206 126896 453212 126908
rect 453264 126896 453270 126948
rect 576118 126896 576124 126948
rect 576176 126936 576182 126948
rect 580166 126936 580172 126948
rect 576176 126908 580172 126936
rect 576176 126896 576182 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 451734 124720 451740 124772
rect 451792 124760 451798 124772
rect 453850 124760 453856 124772
rect 451792 124732 453856 124760
rect 451792 124720 451798 124732
rect 453850 124720 453856 124732
rect 453908 124720 453914 124772
rect 451734 123088 451740 123140
rect 451792 123128 451798 123140
rect 454862 123128 454868 123140
rect 451792 123100 454868 123128
rect 451792 123088 451798 123100
rect 454862 123088 454868 123100
rect 454920 123088 454926 123140
rect 451734 121592 451740 121644
rect 451792 121632 451798 121644
rect 454954 121632 454960 121644
rect 451792 121604 454960 121632
rect 451792 121592 451798 121604
rect 454954 121592 454960 121604
rect 455012 121592 455018 121644
rect 369026 120232 369032 120284
rect 369084 120272 369090 120284
rect 373626 120272 373632 120284
rect 369084 120244 373632 120272
rect 369084 120232 369090 120244
rect 373626 120232 373632 120244
rect 373684 120232 373690 120284
rect 362402 117920 362408 117972
rect 362460 117960 362466 117972
rect 369026 117960 369032 117972
rect 362460 117932 369032 117960
rect 362460 117920 362466 117932
rect 369026 117920 369032 117932
rect 369084 117920 369090 117972
rect 361574 117240 361580 117292
rect 361632 117280 361638 117292
rect 409322 117280 409328 117292
rect 361632 117252 409328 117280
rect 361632 117240 361638 117252
rect 409322 117240 409328 117252
rect 409380 117240 409386 117292
rect 573358 113092 573364 113144
rect 573416 113132 573422 113144
rect 579798 113132 579804 113144
rect 573416 113104 579804 113132
rect 573416 113092 573422 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 359642 106904 359648 106956
rect 359700 106944 359706 106956
rect 362402 106944 362408 106956
rect 359700 106916 362408 106944
rect 359700 106904 359706 106916
rect 362402 106904 362408 106916
rect 362460 106904 362466 106956
rect 361574 106224 361580 106276
rect 361632 106264 361638 106276
rect 407850 106264 407856 106276
rect 361632 106236 407856 106264
rect 361632 106224 361638 106236
rect 407850 106224 407856 106236
rect 407908 106224 407914 106276
rect 569218 100648 569224 100700
rect 569276 100688 569282 100700
rect 580166 100688 580172 100700
rect 569276 100660 580172 100688
rect 569276 100648 569282 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 361758 95140 361764 95192
rect 361816 95180 361822 95192
rect 410610 95180 410616 95192
rect 361816 95152 410616 95180
rect 361816 95140 361822 95152
rect 410610 95140 410616 95152
rect 410668 95140 410674 95192
rect 394602 88952 394608 89004
rect 394660 88992 394666 89004
rect 404078 88992 404084 89004
rect 394660 88964 404084 88992
rect 394660 88952 394666 88964
rect 404078 88952 404084 88964
rect 404136 88952 404142 89004
rect 574738 86912 574744 86964
rect 574796 86952 574802 86964
rect 580166 86952 580172 86964
rect 574796 86924 580172 86952
rect 574796 86912 574802 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3418 86232 3424 86284
rect 3476 86272 3482 86284
rect 20898 86272 20904 86284
rect 3476 86244 20904 86272
rect 3476 86232 3482 86244
rect 20898 86232 20904 86244
rect 20956 86232 20962 86284
rect 388438 85552 388444 85604
rect 388496 85592 388502 85604
rect 394602 85592 394608 85604
rect 388496 85564 394608 85592
rect 388496 85552 388502 85564
rect 394602 85552 394608 85564
rect 394660 85552 394666 85604
rect 361758 84124 361764 84176
rect 361816 84164 361822 84176
rect 404170 84164 404176 84176
rect 361816 84136 404176 84164
rect 361816 84124 361822 84136
rect 404170 84124 404176 84136
rect 404228 84124 404234 84176
rect 361758 73108 361764 73160
rect 361816 73148 361822 73160
rect 410518 73148 410524 73160
rect 361816 73120 410524 73148
rect 361816 73108 361822 73120
rect 410518 73108 410524 73120
rect 410576 73108 410582 73160
rect 548518 73108 548524 73160
rect 548576 73148 548582 73160
rect 580166 73148 580172 73160
rect 548576 73120 580172 73148
rect 548576 73108 548582 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 4798 68960 4804 69012
rect 4856 69000 4862 69012
rect 7374 69000 7380 69012
rect 4856 68972 7380 69000
rect 4856 68960 4862 68972
rect 7374 68960 7380 68972
rect 7432 68960 7438 69012
rect 7374 67464 7380 67516
rect 7432 67504 7438 67516
rect 8662 67504 8668 67516
rect 7432 67476 8668 67504
rect 7432 67464 7438 67476
rect 8662 67464 8668 67476
rect 8720 67464 8726 67516
rect 4982 66172 4988 66224
rect 5040 66212 5046 66224
rect 5810 66212 5816 66224
rect 5040 66184 5816 66212
rect 5040 66172 5046 66184
rect 5810 66172 5816 66184
rect 5868 66172 5874 66224
rect 359734 63520 359740 63572
rect 359792 63560 359798 63572
rect 362310 63560 362316 63572
rect 359792 63532 362316 63560
rect 359792 63520 359798 63532
rect 362310 63520 362316 63532
rect 362368 63520 362374 63572
rect 449894 62772 449900 62824
rect 449952 62812 449958 62824
rect 537478 62812 537484 62824
rect 449952 62784 537484 62812
rect 449952 62772 449958 62784
rect 537478 62772 537484 62784
rect 537536 62772 537542 62824
rect 5810 62092 5816 62144
rect 5868 62132 5874 62144
rect 5868 62104 6914 62132
rect 5868 62092 5874 62104
rect 6886 62064 6914 62104
rect 9582 62064 9588 62076
rect 6886 62036 9588 62064
rect 9582 62024 9588 62036
rect 9640 62024 9646 62076
rect 361758 62024 361764 62076
rect 361816 62064 361822 62076
rect 406838 62064 406844 62076
rect 361816 62036 406844 62064
rect 361816 62024 361822 62036
rect 406838 62024 406844 62036
rect 406896 62024 406902 62076
rect 5074 61276 5080 61328
rect 5132 61316 5138 61328
rect 5534 61316 5540 61328
rect 5132 61288 5540 61316
rect 5132 61276 5138 61288
rect 5534 61276 5540 61288
rect 5592 61276 5598 61328
rect 385678 61208 385684 61260
rect 385736 61248 385742 61260
rect 388438 61248 388444 61260
rect 385736 61220 388444 61248
rect 385736 61208 385742 61220
rect 388438 61208 388444 61220
rect 388496 61208 388502 61260
rect 544378 60664 544384 60716
rect 544436 60704 544442 60716
rect 580166 60704 580172 60716
rect 544436 60676 580172 60704
rect 544436 60664 544442 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3602 59984 3608 60036
rect 3660 60024 3666 60036
rect 20898 60024 20904 60036
rect 3660 59996 20904 60024
rect 3660 59984 3666 59996
rect 20898 59984 20904 59996
rect 20956 59984 20962 60036
rect 8662 59304 8668 59356
rect 8720 59344 8726 59356
rect 10318 59344 10324 59356
rect 8720 59316 10324 59344
rect 8720 59304 8726 59316
rect 10318 59304 10324 59316
rect 10376 59304 10382 59356
rect 372614 58624 372620 58676
rect 372672 58664 372678 58676
rect 385678 58664 385684 58676
rect 372672 58636 385684 58664
rect 372672 58624 372678 58636
rect 385678 58624 385684 58636
rect 385736 58624 385742 58676
rect 9674 57944 9680 57996
rect 9732 57984 9738 57996
rect 9732 57956 11100 57984
rect 9732 57944 9738 57956
rect 4890 57876 4896 57928
rect 4948 57916 4954 57928
rect 6086 57916 6092 57928
rect 4948 57888 6092 57916
rect 4948 57876 4954 57888
rect 6086 57876 6092 57888
rect 6144 57876 6150 57928
rect 11072 57916 11100 57956
rect 13722 57916 13728 57928
rect 11072 57888 13728 57916
rect 13722 57876 13728 57888
rect 13780 57876 13786 57928
rect 5534 57196 5540 57248
rect 5592 57236 5598 57248
rect 15194 57236 15200 57248
rect 5592 57208 15200 57236
rect 5592 57196 5598 57208
rect 15194 57196 15200 57208
rect 15252 57196 15258 57248
rect 368290 56312 368296 56364
rect 368348 56352 368354 56364
rect 372614 56352 372620 56364
rect 368348 56324 372620 56352
rect 368348 56312 368354 56324
rect 372614 56312 372620 56324
rect 372672 56312 372678 56364
rect 6086 54476 6092 54528
rect 6144 54516 6150 54528
rect 8202 54516 8208 54528
rect 6144 54488 8208 54516
rect 6144 54476 6150 54488
rect 8202 54476 8208 54488
rect 8260 54476 8266 54528
rect 15194 54476 15200 54528
rect 15252 54516 15258 54528
rect 20898 54516 20904 54528
rect 15252 54488 20904 54516
rect 15252 54476 15258 54488
rect 20898 54476 20904 54488
rect 20956 54476 20962 54528
rect 5166 53796 5172 53848
rect 5224 53836 5230 53848
rect 5224 53808 6914 53836
rect 5224 53796 5230 53808
rect 6886 53768 6914 53808
rect 7374 53768 7380 53780
rect 6886 53740 7380 53768
rect 7374 53728 7380 53740
rect 7432 53728 7438 53780
rect 13722 53728 13728 53780
rect 13780 53768 13786 53780
rect 19242 53768 19248 53780
rect 13780 53740 19248 53768
rect 13780 53728 13786 53740
rect 19242 53728 19248 53740
rect 19300 53728 19306 53780
rect 361758 52368 361764 52420
rect 361816 52408 361822 52420
rect 407758 52408 407764 52420
rect 361816 52380 407764 52408
rect 361816 52368 361822 52380
rect 407758 52368 407764 52380
rect 407816 52368 407822 52420
rect 10318 51756 10324 51808
rect 10376 51796 10382 51808
rect 11238 51796 11244 51808
rect 10376 51768 11244 51796
rect 10376 51756 10382 51768
rect 11238 51756 11244 51768
rect 11296 51756 11302 51808
rect 540606 51076 540612 51128
rect 540664 51116 540670 51128
rect 543734 51116 543740 51128
rect 540664 51088 543740 51116
rect 540664 51076 540670 51088
rect 543734 51076 543740 51088
rect 543792 51076 543798 51128
rect 7374 50804 7380 50856
rect 7432 50844 7438 50856
rect 11330 50844 11336 50856
rect 7432 50816 11336 50844
rect 7432 50804 7438 50816
rect 11330 50804 11336 50816
rect 11388 50804 11394 50856
rect 8294 48288 8300 48340
rect 8352 48328 8358 48340
rect 8352 48300 9720 48328
rect 8352 48288 8358 48300
rect 9692 48260 9720 48300
rect 11238 48288 11244 48340
rect 11296 48328 11302 48340
rect 11296 48300 12480 48328
rect 11296 48288 11302 48300
rect 11422 48260 11428 48272
rect 9692 48232 11428 48260
rect 11422 48220 11428 48232
rect 11480 48220 11486 48272
rect 12452 48260 12480 48300
rect 16482 48260 16488 48272
rect 12452 48232 16488 48260
rect 16482 48220 16488 48232
rect 16540 48220 16546 48272
rect 11330 48152 11336 48204
rect 11388 48192 11394 48204
rect 15194 48192 15200 48204
rect 11388 48164 15200 48192
rect 11388 48152 11394 48164
rect 15194 48152 15200 48164
rect 15252 48152 15258 48204
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 456518 47036 456524 47048
rect 3292 47008 456524 47036
rect 3292 46996 3298 47008
rect 456518 46996 456524 47008
rect 456576 46996 456582 47048
rect 3418 46860 3424 46912
rect 3476 46900 3482 46912
rect 460290 46900 460296 46912
rect 3476 46872 460296 46900
rect 3476 46860 3482 46872
rect 460290 46860 460296 46872
rect 460348 46860 460354 46912
rect 563698 46860 563704 46912
rect 563756 46900 563762 46912
rect 580166 46900 580172 46912
rect 563756 46872 580172 46900
rect 563756 46860 563762 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3602 46792 3608 46844
rect 3660 46832 3666 46844
rect 460382 46832 460388 46844
rect 3660 46804 460388 46832
rect 3660 46792 3666 46804
rect 460382 46792 460388 46804
rect 460440 46792 460446 46844
rect 4062 46724 4068 46776
rect 4120 46764 4126 46776
rect 459002 46764 459008 46776
rect 4120 46736 459008 46764
rect 4120 46724 4126 46736
rect 459002 46724 459008 46736
rect 459060 46724 459066 46776
rect 3326 46656 3332 46708
rect 3384 46696 3390 46708
rect 456334 46696 456340 46708
rect 3384 46668 456340 46696
rect 3384 46656 3390 46668
rect 456334 46656 456340 46668
rect 456392 46656 456398 46708
rect 3786 46588 3792 46640
rect 3844 46628 3850 46640
rect 456426 46628 456432 46640
rect 3844 46600 456432 46628
rect 3844 46588 3850 46600
rect 456426 46588 456432 46600
rect 456484 46588 456490 46640
rect 3694 46520 3700 46572
rect 3752 46560 3758 46572
rect 453574 46560 453580 46572
rect 3752 46532 453580 46560
rect 3752 46520 3758 46532
rect 453574 46520 453580 46532
rect 453632 46520 453638 46572
rect 3878 46452 3884 46504
rect 3936 46492 3942 46504
rect 453482 46492 453488 46504
rect 3936 46464 453488 46492
rect 3936 46452 3942 46464
rect 453482 46452 453488 46464
rect 453540 46452 453546 46504
rect 3510 46384 3516 46436
rect 3568 46424 3574 46436
rect 450906 46424 450912 46436
rect 3568 46396 450912 46424
rect 3568 46384 3574 46396
rect 450906 46384 450912 46396
rect 450964 46384 450970 46436
rect 19978 46316 19984 46368
rect 20036 46356 20042 46368
rect 457438 46356 457444 46368
rect 20036 46328 457444 46356
rect 20036 46316 20042 46328
rect 457438 46316 457444 46328
rect 457496 46316 457502 46368
rect 21450 46248 21456 46300
rect 21508 46288 21514 46300
rect 451090 46288 451096 46300
rect 21508 46260 451096 46288
rect 21508 46248 21514 46260
rect 451090 46248 451096 46260
rect 451148 46248 451154 46300
rect 21358 46180 21364 46232
rect 21416 46220 21422 46232
rect 450998 46220 451004 46232
rect 21416 46192 451004 46220
rect 21416 46180 21422 46192
rect 450998 46180 451004 46192
rect 451056 46180 451062 46232
rect 15194 46112 15200 46164
rect 15252 46152 15258 46164
rect 359734 46152 359740 46164
rect 15252 46124 359740 46152
rect 15252 46112 15258 46124
rect 359734 46112 359740 46124
rect 359792 46112 359798 46164
rect 358722 46044 358728 46096
rect 358780 46084 358786 46096
rect 368290 46084 368296 46096
rect 358780 46056 368296 46084
rect 358780 46044 358786 46056
rect 368290 46044 368296 46056
rect 368348 46044 368354 46096
rect 3970 45500 3976 45552
rect 4028 45540 4034 45552
rect 453390 45540 453396 45552
rect 4028 45512 453396 45540
rect 4028 45500 4034 45512
rect 453390 45500 453396 45512
rect 453448 45500 453454 45552
rect 3418 45432 3424 45484
rect 3476 45472 3482 45484
rect 399478 45472 399484 45484
rect 3476 45444 399484 45472
rect 3476 45432 3482 45444
rect 399478 45432 399484 45444
rect 399536 45432 399542 45484
rect 11422 45364 11428 45416
rect 11480 45404 11486 45416
rect 361298 45404 361304 45416
rect 11480 45376 361304 45404
rect 11480 45364 11486 45376
rect 361298 45364 361304 45376
rect 361356 45364 361362 45416
rect 16574 45296 16580 45348
rect 16632 45336 16638 45348
rect 358722 45336 358728 45348
rect 16632 45308 358728 45336
rect 16632 45296 16638 45308
rect 358722 45296 358728 45308
rect 358780 45296 358786 45348
rect 69014 45228 69020 45280
rect 69072 45268 69078 45280
rect 406654 45268 406660 45280
rect 69072 45240 406660 45268
rect 69072 45228 69078 45240
rect 406654 45228 406660 45240
rect 406712 45228 406718 45280
rect 64874 45160 64880 45212
rect 64932 45200 64938 45212
rect 406378 45200 406384 45212
rect 64932 45172 406384 45200
rect 64932 45160 64938 45172
rect 406378 45160 406384 45172
rect 406436 45160 406442 45212
rect 60734 45092 60740 45144
rect 60792 45132 60798 45144
rect 406562 45132 406568 45144
rect 60792 45104 406568 45132
rect 60792 45092 60798 45104
rect 406562 45092 406568 45104
rect 406620 45092 406626 45144
rect 57974 45024 57980 45076
rect 58032 45064 58038 45076
rect 406470 45064 406476 45076
rect 58032 45036 406476 45064
rect 58032 45024 58038 45036
rect 406470 45024 406476 45036
rect 406528 45024 406534 45076
rect 51074 44956 51080 45008
rect 51132 44996 51138 45008
rect 406746 44996 406752 45008
rect 51132 44968 406752 44996
rect 51132 44956 51138 44968
rect 406746 44956 406752 44968
rect 406804 44956 406810 45008
rect 46934 44888 46940 44940
rect 46992 44928 46998 44940
rect 409138 44928 409144 44940
rect 46992 44900 409144 44928
rect 46992 44888 46998 44900
rect 409138 44888 409144 44900
rect 409196 44888 409202 44940
rect 53834 44820 53840 44872
rect 53892 44860 53898 44872
rect 456242 44860 456248 44872
rect 53892 44832 456248 44860
rect 53892 44820 53898 44832
rect 456242 44820 456248 44832
rect 456300 44820 456306 44872
rect 71774 44752 71780 44804
rect 71832 44792 71838 44804
rect 403986 44792 403992 44804
rect 71832 44764 403992 44792
rect 71832 44752 71838 44764
rect 403986 44752 403992 44764
rect 404044 44752 404050 44804
rect 86954 44684 86960 44736
rect 87012 44724 87018 44736
rect 387518 44724 387524 44736
rect 87012 44696 387524 44724
rect 87012 44684 87018 44696
rect 387518 44684 387524 44696
rect 387576 44684 387582 44736
rect 107654 44616 107660 44668
rect 107712 44656 107718 44668
rect 398374 44656 398380 44668
rect 107712 44628 398380 44656
rect 107712 44616 107718 44628
rect 398374 44616 398380 44628
rect 398432 44616 398438 44668
rect 103514 42712 103520 42764
rect 103572 42752 103578 42764
rect 398282 42752 398288 42764
rect 103572 42724 398288 42752
rect 103572 42712 103578 42724
rect 398282 42712 398288 42724
rect 398340 42712 398346 42764
rect 100754 42644 100760 42696
rect 100812 42684 100818 42696
rect 401134 42684 401140 42696
rect 100812 42656 401140 42684
rect 100812 42644 100818 42656
rect 401134 42644 401140 42656
rect 401192 42644 401198 42696
rect 74534 42576 74540 42628
rect 74592 42616 74598 42628
rect 376478 42616 376484 42628
rect 74592 42588 376484 42616
rect 74592 42576 74598 42588
rect 376478 42576 376484 42588
rect 376536 42576 376542 42628
rect 96614 42508 96620 42560
rect 96672 42548 96678 42560
rect 401042 42548 401048 42560
rect 96672 42520 401048 42548
rect 96672 42508 96678 42520
rect 401042 42508 401048 42520
rect 401100 42508 401106 42560
rect 93854 42440 93860 42492
rect 93912 42480 93918 42492
rect 401226 42480 401232 42492
rect 93912 42452 401232 42480
rect 93912 42440 93918 42452
rect 401226 42440 401232 42452
rect 401284 42440 401290 42492
rect 89714 42372 89720 42424
rect 89772 42412 89778 42424
rect 400950 42412 400956 42424
rect 89772 42384 400956 42412
rect 89772 42372 89778 42384
rect 400950 42372 400956 42384
rect 401008 42372 401014 42424
rect 85574 42304 85580 42356
rect 85632 42344 85638 42356
rect 401318 42344 401324 42356
rect 85632 42316 401324 42344
rect 85632 42304 85638 42316
rect 401318 42304 401324 42316
rect 401376 42304 401382 42356
rect 82814 42236 82820 42288
rect 82872 42276 82878 42288
rect 403802 42276 403808 42288
rect 82872 42248 403808 42276
rect 82872 42236 82878 42248
rect 403802 42236 403808 42248
rect 403860 42236 403866 42288
rect 78674 42168 78680 42220
rect 78732 42208 78738 42220
rect 403710 42208 403716 42220
rect 78732 42180 403716 42208
rect 78732 42168 78738 42180
rect 403710 42168 403716 42180
rect 403768 42168 403774 42220
rect 75914 42100 75920 42152
rect 75972 42140 75978 42152
rect 403618 42140 403624 42152
rect 75972 42112 403624 42140
rect 75972 42100 75978 42112
rect 403618 42100 403624 42112
rect 403676 42100 403682 42152
rect 11054 42032 11060 42084
rect 11112 42072 11118 42084
rect 403894 42072 403900 42084
rect 11112 42044 403900 42072
rect 11112 42032 11118 42044
rect 403894 42032 403900 42044
rect 403952 42032 403958 42084
rect 110414 41964 110420 42016
rect 110472 42004 110478 42016
rect 398190 42004 398196 42016
rect 110472 41976 398196 42004
rect 110472 41964 110478 41976
rect 398190 41964 398196 41976
rect 398248 41964 398254 42016
rect 111794 41896 111800 41948
rect 111852 41936 111858 41948
rect 384574 41936 384580 41948
rect 111852 41908 384580 41936
rect 111852 41896 111858 41908
rect 384574 41896 384580 41908
rect 384632 41896 384638 41948
rect 114554 39992 114560 40044
rect 114612 40032 114618 40044
rect 398098 40032 398104 40044
rect 114612 40004 398104 40032
rect 114612 39992 114618 40004
rect 398098 39992 398104 40004
rect 398156 39992 398162 40044
rect 91094 39924 91100 39976
rect 91152 39964 91158 39976
rect 387334 39964 387340 39976
rect 91152 39936 387340 39964
rect 91152 39924 91158 39936
rect 387334 39924 387340 39936
rect 387392 39924 387398 39976
rect 59354 39856 59360 39908
rect 59412 39896 59418 39908
rect 393038 39896 393044 39908
rect 59412 39868 393044 39896
rect 59412 39856 59418 39868
rect 393038 39856 393044 39868
rect 393096 39856 393102 39908
rect 55214 39788 55220 39840
rect 55272 39828 55278 39840
rect 392946 39828 392952 39840
rect 55272 39800 392952 39828
rect 55272 39788 55278 39800
rect 392946 39788 392952 39800
rect 393004 39788 393010 39840
rect 118694 39720 118700 39772
rect 118752 39760 118758 39772
rect 460198 39760 460204 39772
rect 118752 39732 460204 39760
rect 118752 39720 118758 39732
rect 460198 39720 460204 39732
rect 460256 39720 460262 39772
rect 44174 39652 44180 39704
rect 44232 39692 44238 39704
rect 395614 39692 395620 39704
rect 44232 39664 395620 39692
rect 44232 39652 44238 39664
rect 395614 39652 395620 39664
rect 395672 39652 395678 39704
rect 40034 39584 40040 39636
rect 40092 39624 40098 39636
rect 395430 39624 395436 39636
rect 40092 39596 395436 39624
rect 40092 39584 40098 39596
rect 395430 39584 395436 39596
rect 395488 39584 395494 39636
rect 35894 39516 35900 39568
rect 35952 39556 35958 39568
rect 395798 39556 395804 39568
rect 35952 39528 395804 39556
rect 35952 39516 35958 39528
rect 395798 39516 395804 39528
rect 395856 39516 395862 39568
rect 20714 39448 20720 39500
rect 20772 39488 20778 39500
rect 395522 39488 395528 39500
rect 20772 39460 395528 39488
rect 20772 39448 20778 39460
rect 395522 39448 395528 39460
rect 395580 39448 395586 39500
rect 2774 39380 2780 39432
rect 2832 39420 2838 39432
rect 395706 39420 395712 39432
rect 2832 39392 395712 39420
rect 2832 39380 2838 39392
rect 395706 39380 395712 39392
rect 395764 39380 395770 39432
rect 33134 39312 33140 39364
rect 33192 39352 33198 39364
rect 450814 39352 450820 39364
rect 33192 39324 450820 39352
rect 33192 39312 33198 39324
rect 450814 39312 450820 39324
rect 450872 39312 450878 39364
rect 104894 37204 104900 37256
rect 104952 37244 104958 37256
rect 387426 37244 387432 37256
rect 104952 37216 387432 37244
rect 104952 37204 104958 37216
rect 387426 37204 387432 37216
rect 387484 37204 387490 37256
rect 102134 37136 102140 37188
rect 102192 37176 102198 37188
rect 387150 37176 387156 37188
rect 102192 37148 387156 37176
rect 102192 37136 102198 37148
rect 387150 37136 387156 37148
rect 387208 37136 387214 37188
rect 97994 37068 98000 37120
rect 98052 37108 98058 37120
rect 387058 37108 387064 37120
rect 98052 37080 387064 37108
rect 98052 37068 98058 37080
rect 387058 37068 387064 37080
rect 387116 37068 387122 37120
rect 93946 37000 93952 37052
rect 94004 37040 94010 37052
rect 387242 37040 387248 37052
rect 94004 37012 387248 37040
rect 94004 37000 94010 37012
rect 387242 37000 387248 37012
rect 387300 37000 387306 37052
rect 84194 36932 84200 36984
rect 84252 36972 84258 36984
rect 390094 36972 390100 36984
rect 84252 36944 390100 36972
rect 84252 36932 84258 36944
rect 390094 36932 390100 36944
rect 390152 36932 390158 36984
rect 80054 36864 80060 36916
rect 80112 36904 80118 36916
rect 390278 36904 390284 36916
rect 80112 36876 390284 36904
rect 80112 36864 80118 36876
rect 390278 36864 390284 36876
rect 390336 36864 390342 36916
rect 77294 36796 77300 36848
rect 77352 36836 77358 36848
rect 389910 36836 389916 36848
rect 77352 36808 389916 36836
rect 77352 36796 77358 36808
rect 389910 36796 389916 36808
rect 389968 36796 389974 36848
rect 73154 36728 73160 36780
rect 73212 36768 73218 36780
rect 390002 36768 390008 36780
rect 73212 36740 390008 36768
rect 73212 36728 73218 36740
rect 390002 36728 390008 36740
rect 390060 36728 390066 36780
rect 69106 36660 69112 36712
rect 69164 36700 69170 36712
rect 390186 36700 390192 36712
rect 69164 36672 390192 36700
rect 69164 36660 69170 36672
rect 390186 36660 390192 36672
rect 390244 36660 390250 36712
rect 66254 36592 66260 36644
rect 66312 36632 66318 36644
rect 392854 36632 392860 36644
rect 66312 36604 392860 36632
rect 66312 36592 66318 36604
rect 392854 36592 392860 36604
rect 392912 36592 392918 36644
rect 62114 36524 62120 36576
rect 62172 36564 62178 36576
rect 392762 36564 392768 36576
rect 62172 36536 392768 36564
rect 62172 36524 62178 36536
rect 392762 36524 392768 36536
rect 392820 36524 392826 36576
rect 109034 36456 109040 36508
rect 109092 36496 109098 36508
rect 384482 36496 384488 36508
rect 109092 36468 384488 36496
rect 109092 36456 109098 36468
rect 384482 36456 384488 36468
rect 384540 36456 384546 36508
rect 115934 36388 115940 36440
rect 115992 36428 115998 36440
rect 384390 36428 384396 36440
rect 115992 36400 384396 36428
rect 115992 36388 115998 36400
rect 384390 36388 384396 36400
rect 384448 36388 384454 36440
rect 60826 34416 60832 34468
rect 60884 34456 60890 34468
rect 376386 34456 376392 34468
rect 60884 34428 376392 34456
rect 60884 34416 60890 34428
rect 376386 34416 376392 34428
rect 376444 34416 376450 34468
rect 56594 34348 56600 34400
rect 56652 34388 56658 34400
rect 379146 34388 379152 34400
rect 56652 34360 379152 34388
rect 56652 34348 56658 34360
rect 379146 34348 379152 34360
rect 379204 34348 379210 34400
rect 49694 34280 49700 34332
rect 49752 34320 49758 34332
rect 379238 34320 379244 34332
rect 49752 34292 379244 34320
rect 49752 34280 49758 34292
rect 379238 34280 379244 34292
rect 379296 34280 379302 34332
rect 44266 34212 44272 34264
rect 44324 34252 44330 34264
rect 378870 34252 378876 34264
rect 44324 34224 378876 34252
rect 44324 34212 44330 34224
rect 378870 34212 378876 34224
rect 378928 34212 378934 34264
rect 41414 34144 41420 34196
rect 41472 34184 41478 34196
rect 378962 34184 378968 34196
rect 41472 34156 378968 34184
rect 41472 34144 41478 34156
rect 378962 34144 378968 34156
rect 379020 34144 379026 34196
rect 37274 34076 37280 34128
rect 37332 34116 37338 34128
rect 379054 34116 379060 34128
rect 37332 34088 379060 34116
rect 37332 34076 37338 34088
rect 379054 34076 379060 34088
rect 379112 34076 379118 34128
rect 34514 34008 34520 34060
rect 34572 34048 34578 34060
rect 381998 34048 382004 34060
rect 34572 34020 382004 34048
rect 34572 34008 34578 34020
rect 381998 34008 382004 34020
rect 382056 34008 382062 34060
rect 30374 33940 30380 33992
rect 30432 33980 30438 33992
rect 381814 33980 381820 33992
rect 30432 33952 381820 33980
rect 30432 33940 30438 33952
rect 381814 33940 381820 33952
rect 381872 33940 381878 33992
rect 22094 33872 22100 33924
rect 22152 33912 22158 33924
rect 381906 33912 381912 33924
rect 22152 33884 381912 33912
rect 22152 33872 22158 33884
rect 381906 33872 381912 33884
rect 381964 33872 381970 33924
rect 17954 33804 17960 33856
rect 18012 33844 18018 33856
rect 384298 33844 384304 33856
rect 18012 33816 384304 33844
rect 18012 33804 18018 33816
rect 384298 33804 384304 33816
rect 384356 33804 384362 33856
rect 9674 33736 9680 33788
rect 9732 33776 9738 33788
rect 378778 33776 378784 33788
rect 9732 33748 378784 33776
rect 9732 33736 9738 33748
rect 378778 33736 378784 33748
rect 378836 33736 378842 33788
rect 118786 33668 118792 33720
rect 118844 33708 118850 33720
rect 381722 33708 381728 33720
rect 118844 33680 381728 33708
rect 118844 33668 118850 33680
rect 381722 33668 381728 33680
rect 381780 33668 381786 33720
rect 122834 33600 122840 33652
rect 122892 33640 122898 33652
rect 381538 33640 381544 33652
rect 122892 33612 381544 33640
rect 122892 33600 122898 33612
rect 381538 33600 381544 33612
rect 381596 33600 381602 33652
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 400858 33096 400864 33108
rect 3568 33068 400864 33096
rect 3568 33056 3574 33068
rect 400858 33056 400864 33068
rect 400916 33056 400922 33108
rect 565078 33056 565084 33108
rect 565136 33096 565142 33108
rect 580166 33096 580172 33108
rect 565136 33068 580172 33096
rect 565136 33056 565142 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 113174 31696 113180 31748
rect 113232 31736 113238 31748
rect 370958 31736 370964 31748
rect 113232 31708 370964 31736
rect 113232 31696 113238 31708
rect 370958 31696 370964 31708
rect 371016 31696 371022 31748
rect 106274 31628 106280 31680
rect 106332 31668 106338 31680
rect 370682 31668 370688 31680
rect 106332 31640 370688 31668
rect 106332 31628 106338 31640
rect 370682 31628 370688 31640
rect 370740 31628 370746 31680
rect 99374 31560 99380 31612
rect 99432 31600 99438 31612
rect 370774 31600 370780 31612
rect 99432 31572 370780 31600
rect 99432 31560 99438 31572
rect 370774 31560 370780 31572
rect 370832 31560 370838 31612
rect 95234 31492 95240 31544
rect 95292 31532 95298 31544
rect 373350 31532 373356 31544
rect 95292 31504 373356 31532
rect 95292 31492 95298 31504
rect 373350 31492 373356 31504
rect 373408 31492 373414 31544
rect 88334 31424 88340 31476
rect 88392 31464 88398 31476
rect 373534 31464 373540 31476
rect 88392 31436 373540 31464
rect 88392 31424 88398 31436
rect 373534 31424 373540 31436
rect 373592 31424 373598 31476
rect 85666 31356 85672 31408
rect 85724 31396 85730 31408
rect 373258 31396 373264 31408
rect 85724 31368 373264 31396
rect 85724 31356 85730 31368
rect 373258 31356 373264 31368
rect 373316 31356 373322 31408
rect 77386 31288 77392 31340
rect 77444 31328 77450 31340
rect 373442 31328 373448 31340
rect 77444 31300 373448 31328
rect 77444 31288 77450 31300
rect 373442 31288 373448 31300
rect 373500 31288 373506 31340
rect 70394 31220 70400 31272
rect 70452 31260 70458 31272
rect 376202 31260 376208 31272
rect 70452 31232 376208 31260
rect 70452 31220 70458 31232
rect 376202 31220 376208 31232
rect 376260 31220 376266 31272
rect 67634 31152 67640 31204
rect 67692 31192 67698 31204
rect 376110 31192 376116 31204
rect 67692 31164 376116 31192
rect 67692 31152 67698 31164
rect 376110 31152 376116 31164
rect 376168 31152 376174 31204
rect 63494 31084 63500 31136
rect 63552 31124 63558 31136
rect 376294 31124 376300 31136
rect 63552 31096 376300 31124
rect 63552 31084 63558 31096
rect 376294 31084 376300 31096
rect 376352 31084 376358 31136
rect 19334 31016 19340 31068
rect 19392 31056 19398 31068
rect 370866 31056 370872 31068
rect 19392 31028 370872 31056
rect 19392 31016 19398 31028
rect 370866 31016 370872 31028
rect 370924 31016 370930 31068
rect 117314 30948 117320 31000
rect 117372 30988 117378 31000
rect 370498 30988 370504 31000
rect 117372 30960 370504 30988
rect 117372 30948 117378 30960
rect 370498 30948 370504 30960
rect 370556 30948 370562 31000
rect 120074 30880 120080 30932
rect 120132 30920 120138 30932
rect 370590 30920 370596 30932
rect 120132 30892 370596 30920
rect 120132 30880 120138 30892
rect 370590 30880 370596 30892
rect 370648 30880 370654 30932
rect 45554 28432 45560 28484
rect 45612 28472 45618 28484
rect 368014 28472 368020 28484
rect 45612 28444 368020 28472
rect 45612 28432 45618 28444
rect 368014 28432 368020 28444
rect 368072 28432 368078 28484
rect 42794 28364 42800 28416
rect 42852 28404 42858 28416
rect 367830 28404 367836 28416
rect 42852 28376 367836 28404
rect 42852 28364 42858 28376
rect 367830 28364 367836 28376
rect 367888 28364 367894 28416
rect 38654 28296 38660 28348
rect 38712 28336 38718 28348
rect 367922 28336 367928 28348
rect 38712 28308 367928 28336
rect 38712 28296 38718 28308
rect 367922 28296 367928 28308
rect 367980 28296 367986 28348
rect 31754 28228 31760 28280
rect 31812 28268 31818 28280
rect 368106 28268 368112 28280
rect 31812 28240 368112 28268
rect 31812 28228 31818 28240
rect 368106 28228 368112 28240
rect 368164 28228 368170 28280
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 376018 20652 376024 20664
rect 3476 20624 376024 20652
rect 3476 20612 3482 20624
rect 376018 20612 376024 20624
rect 376076 20612 376082 20664
rect 566458 20612 566464 20664
rect 566516 20652 566522 20664
rect 579982 20652 579988 20664
rect 566516 20624 579988 20652
rect 566516 20612 566522 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 396718 6848 396724 6860
rect 3476 6820 396724 6848
rect 3476 6808 3482 6820
rect 396718 6808 396724 6820
rect 396776 6808 396782 6860
rect 562318 6808 562324 6860
rect 562376 6848 562382 6860
rect 580166 6848 580172 6860
rect 562376 6820 580172 6848
rect 562376 6808 562382 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 52546 4088 52552 4140
rect 52604 4128 52610 4140
rect 359458 4128 359464 4140
rect 52604 4100 359464 4128
rect 52604 4088 52610 4100
rect 359458 4088 359464 4100
rect 359516 4088 359522 4140
rect 35986 4020 35992 4072
rect 36044 4060 36050 4072
rect 360930 4060 360936 4072
rect 36044 4032 360936 4060
rect 36044 4020 36050 4032
rect 360930 4020 360936 4032
rect 360988 4020 360994 4072
rect 124674 3952 124680 4004
rect 124732 3992 124738 4004
rect 458818 3992 458824 4004
rect 124732 3964 458824 3992
rect 124732 3952 124738 3964
rect 458818 3952 458824 3964
rect 458876 3952 458882 4004
rect 48958 3884 48964 3936
rect 49016 3924 49022 3936
rect 392670 3924 392676 3936
rect 49016 3896 392676 3924
rect 49016 3884 49022 3896
rect 392670 3884 392676 3896
rect 392728 3884 392734 3936
rect 14734 3816 14740 3868
rect 14792 3856 14798 3868
rect 359550 3856 359556 3868
rect 14792 3828 359556 3856
rect 14792 3816 14798 3828
rect 359550 3816 359556 3828
rect 359608 3816 359614 3868
rect 27706 3748 27712 3800
rect 27764 3788 27770 3800
rect 381630 3788 381636 3800
rect 27764 3760 381636 3788
rect 27764 3748 27770 3760
rect 381630 3748 381636 3760
rect 381688 3748 381694 3800
rect 82078 3680 82084 3732
rect 82136 3720 82142 3732
rect 456058 3720 456064 3732
rect 82136 3692 456064 3720
rect 82136 3680 82142 3692
rect 456058 3680 456064 3692
rect 456116 3680 456122 3732
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 389818 3652 389824 3664
rect 13596 3624 389824 3652
rect 13596 3612 13602 3624
rect 389818 3612 389824 3624
rect 389876 3612 389882 3664
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 395338 3584 395344 3596
rect 17092 3556 395344 3584
rect 17092 3544 17098 3556
rect 395338 3544 395344 3556
rect 395396 3544 395402 3596
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 404998 3516 405004 3528
rect 24268 3488 405004 3516
rect 24268 3476 24274 3488
rect 404998 3476 405004 3488
rect 405056 3476 405062 3528
rect 53742 3408 53748 3460
rect 53800 3448 53806 3460
rect 450630 3448 450636 3460
rect 53800 3420 450636 3448
rect 53800 3408 53806 3420
rect 450630 3408 450636 3420
rect 450688 3408 450694 3460
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 85574 3340 85580 3392
rect 85632 3380 85638 3392
rect 86494 3380 86500 3392
rect 85632 3352 86500 3380
rect 85632 3340 85638 3352
rect 86494 3340 86500 3352
rect 86552 3340 86558 3392
rect 92750 3340 92756 3392
rect 92808 3380 92814 3392
rect 361114 3380 361120 3392
rect 92808 3352 361120 3380
rect 92808 3340 92814 3352
rect 361114 3340 361120 3352
rect 361172 3340 361178 3392
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 360838 3312 360844 3324
rect 103388 3284 360844 3312
rect 103388 3272 103394 3284
rect 360838 3272 360844 3284
rect 360896 3272 360902 3324
rect 110414 3204 110420 3256
rect 110472 3244 110478 3256
rect 111610 3244 111616 3256
rect 110472 3216 111616 3244
rect 110472 3204 110478 3216
rect 111610 3204 111616 3216
rect 111668 3204 111674 3256
rect 361022 3244 361028 3256
rect 113146 3216 361028 3244
rect 110506 3136 110512 3188
rect 110564 3176 110570 3188
rect 113146 3176 113174 3216
rect 361022 3204 361028 3216
rect 361080 3204 361086 3256
rect 110564 3148 113174 3176
rect 110564 3136 110570 3148
rect 30098 2116 30104 2168
rect 30156 2156 30162 2168
rect 450538 2156 450544 2168
rect 30156 2128 450544 2156
rect 30156 2116 30162 2128
rect 450538 2116 450544 2128
rect 450596 2116 450602 2168
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 453298 2088 453304 2100
rect 2924 2060 453304 2088
rect 2924 2048 2930 2060
rect 453298 2048 453304 2060
rect 453356 2048 453362 2100
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 429844 700748 429896 700800
rect 449164 700748 449216 700800
rect 364984 700680 365036 700732
rect 445024 700680 445076 700732
rect 348792 700612 348844 700664
rect 446404 700612 446456 700664
rect 235172 700544 235224 700596
rect 450544 700544 450596 700596
rect 218980 700476 219032 700528
rect 449256 700476 449308 700528
rect 170312 700408 170364 700460
rect 444288 700408 444340 700460
rect 105452 700340 105504 700392
rect 445116 700340 445168 700392
rect 72976 700272 73028 700324
rect 445208 700272 445260 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 573364 696940 573416 696992
rect 580172 696940 580224 696992
rect 299480 687896 299532 687948
rect 449348 687896 449400 687948
rect 266360 686468 266412 686520
rect 446496 686468 446548 686520
rect 88340 685244 88392 685296
rect 418804 685244 418856 685296
rect 23480 685176 23532 685228
rect 446588 685176 446640 685228
rect 6920 685108 6972 685160
rect 446772 685108 446824 685160
rect 3976 684700 4028 684752
rect 420368 684700 420420 684752
rect 3148 684632 3200 684684
rect 420184 684632 420236 684684
rect 3332 684564 3384 684616
rect 420552 684564 420604 684616
rect 3884 684496 3936 684548
rect 446956 684496 447008 684548
rect 331220 683748 331272 683800
rect 418896 683748 418948 683800
rect 20904 683544 20956 683596
rect 359464 683544 359516 683596
rect 19984 683476 20036 683528
rect 417424 683476 417476 683528
rect 4068 683408 4120 683460
rect 420736 683408 420788 683460
rect 3792 683340 3844 683392
rect 420644 683340 420696 683392
rect 3700 683272 3752 683324
rect 445300 683272 445352 683324
rect 3424 683204 3476 683256
rect 445484 683204 445536 683256
rect 3516 683136 3568 683188
rect 446680 683136 446732 683188
rect 576124 683136 576176 683188
rect 580172 683136 580224 683188
rect 2872 682728 2924 682780
rect 420828 682728 420880 682780
rect 2964 682660 3016 682712
rect 447048 682660 447100 682712
rect 18144 680348 18196 680400
rect 20904 680348 20956 680400
rect 361764 678988 361816 679040
rect 382924 678988 382976 679040
rect 3516 678512 3568 678564
rect 3516 678308 3568 678360
rect 16580 675248 16632 675300
rect 18144 675248 18196 675300
rect 567844 670692 567896 670744
rect 580172 670692 580224 670744
rect 13084 667904 13136 667956
rect 16488 667904 16540 667956
rect 361764 667904 361816 667956
rect 378784 667904 378836 667956
rect 8944 662396 8996 662448
rect 13084 662396 13136 662448
rect 361764 656888 361816 656940
rect 400864 656888 400916 656940
rect 4804 652672 4856 652724
rect 8944 652740 8996 652792
rect 361764 645872 361816 645924
rect 376024 645872 376076 645924
rect 361580 634788 361632 634840
rect 403624 634788 403676 634840
rect 3700 631320 3752 631372
rect 19984 631320 20036 631372
rect 574744 630640 574796 630692
rect 580172 630640 580224 630692
rect 361580 623772 361632 623824
rect 374644 623772 374696 623824
rect 361580 612756 361632 612808
rect 406384 612756 406436 612808
rect 359464 609968 359516 610020
rect 365720 609900 365772 609952
rect 365720 607112 365772 607164
rect 367836 607112 367888 607164
rect 458732 602760 458784 602812
rect 459100 602760 459152 602812
rect 361580 601740 361632 601792
rect 371884 601740 371936 601792
rect 367836 601672 367888 601724
rect 369124 601672 369176 601724
rect 457812 600244 457864 600296
rect 461676 600244 461728 600296
rect 457536 600176 457588 600228
rect 461584 600176 461636 600228
rect 459192 599972 459244 600024
rect 462504 599972 462556 600024
rect 458640 599700 458692 599752
rect 465080 599700 465132 599752
rect 457260 599632 457312 599684
rect 465172 599632 465224 599684
rect 457904 599564 457956 599616
rect 468484 599564 468536 599616
rect 515404 599564 515456 599616
rect 580356 599564 580408 599616
rect 459836 598408 459888 598460
rect 463700 598408 463752 598460
rect 458824 598340 458876 598392
rect 467932 598340 467984 598392
rect 484492 598340 484544 598392
rect 494152 598340 494204 598392
rect 457628 598272 457680 598324
rect 468576 598272 468628 598324
rect 477500 598272 477552 598324
rect 494060 598272 494112 598324
rect 447968 598204 448020 598256
rect 505468 598204 505520 598256
rect 491484 597796 491536 597848
rect 494244 597796 494296 597848
rect 459744 596844 459796 596896
rect 463792 596844 463844 596896
rect 457720 596572 457772 596624
rect 461768 596572 461820 596624
rect 457444 595484 457496 595536
rect 464344 595484 464396 595536
rect 449808 595416 449860 595468
rect 469220 595416 469272 595468
rect 369124 595348 369176 595400
rect 370688 595348 370740 595400
rect 459652 594056 459704 594108
rect 466460 594056 466512 594108
rect 370688 593308 370740 593360
rect 372620 593308 372672 593360
rect 361764 590656 361816 590708
rect 370688 590656 370740 590708
rect 511264 590656 511316 590708
rect 580172 590656 580224 590708
rect 372620 590588 372672 590640
rect 376116 590588 376168 590640
rect 376116 582360 376168 582412
rect 378876 582360 378928 582412
rect 361764 579640 361816 579692
rect 367744 579640 367796 579692
rect 378876 574948 378928 575000
rect 380808 574948 380860 575000
rect 380808 571344 380860 571396
rect 385684 571276 385736 571328
rect 361580 568760 361632 568812
rect 363604 568760 363656 568812
rect 515496 563048 515548 563100
rect 579896 563048 579948 563100
rect 385684 560192 385736 560244
rect 387156 560192 387208 560244
rect 361580 557744 361632 557796
rect 363696 557744 363748 557796
rect 387156 556180 387208 556232
rect 388444 556180 388496 556232
rect 361764 546456 361816 546508
rect 407764 546456 407816 546508
rect 457352 542988 457404 543040
rect 466552 542988 466604 543040
rect 514024 536800 514076 536852
rect 580172 536800 580224 536852
rect 459560 536052 459612 536104
rect 469404 536052 469456 536104
rect 361764 535440 361816 535492
rect 410524 535440 410576 535492
rect 361764 524424 361816 524476
rect 411904 524424 411956 524476
rect 457996 523676 458048 523728
rect 467104 523676 467156 523728
rect 388444 522928 388496 522980
rect 389824 522928 389876 522980
rect 458088 522316 458140 522368
rect 468668 522316 468720 522368
rect 448060 522248 448112 522300
rect 462412 522248 462464 522300
rect 459284 520888 459336 520940
rect 470876 520888 470928 520940
rect 482928 520888 482980 520940
rect 518900 520888 518952 520940
rect 449992 520344 450044 520396
rect 488632 520344 488684 520396
rect 389824 520208 389876 520260
rect 391204 520208 391256 520260
rect 450636 519528 450688 519580
rect 512000 519528 512052 519580
rect 459376 518236 459428 518288
rect 470692 518236 470744 518288
rect 448336 518168 448388 518220
rect 498200 518168 498252 518220
rect 480168 517488 480220 517540
rect 482652 517488 482704 517540
rect 448428 516128 448480 516180
rect 491852 516128 491904 516180
rect 494152 515380 494204 515432
rect 538220 515380 538272 515432
rect 3976 514768 4028 514820
rect 4804 514768 4856 514820
rect 361764 513340 361816 513392
rect 414664 513340 414716 513392
rect 494152 512592 494204 512644
rect 494336 512592 494388 512644
rect 535460 512592 535512 512644
rect 494060 507832 494112 507884
rect 532700 507832 532752 507884
rect 494244 505112 494296 505164
rect 529940 505112 529992 505164
rect 361764 502324 361816 502376
rect 416044 502324 416096 502376
rect 448060 501780 448112 501832
rect 448336 501780 448388 501832
rect 391204 500556 391256 500608
rect 393412 500556 393464 500608
rect 448520 500216 448572 500268
rect 545120 500216 545172 500268
rect 447416 499536 447468 499588
rect 449716 499536 449768 499588
rect 447968 499468 448020 499520
rect 494060 499468 494112 499520
rect 448060 499400 448112 499452
rect 494244 499400 494296 499452
rect 449716 498788 449768 498840
rect 542452 498788 542504 498840
rect 457444 497564 457496 497616
rect 482652 497564 482704 497616
rect 453304 497496 453356 497548
rect 480260 497496 480312 497548
rect 451924 497428 451976 497480
rect 491300 497428 491352 497480
rect 454132 497020 454184 497072
rect 459560 497020 459612 497072
rect 454040 496952 454092 497004
rect 458088 496952 458140 497004
rect 452844 496884 452896 496936
rect 455144 496884 455196 496936
rect 455420 496884 455472 496936
rect 461032 496884 461084 496936
rect 451372 496816 451424 496868
rect 453672 496816 453724 496868
rect 454684 496816 454736 496868
rect 456616 496816 456668 496868
rect 393412 496204 393464 496256
rect 397552 496204 397604 496256
rect 449900 496068 449952 496120
rect 547880 496068 547932 496120
rect 449900 494708 449952 494760
rect 450636 494708 450688 494760
rect 361764 491308 361816 491360
rect 417516 491308 417568 491360
rect 397552 489880 397604 489932
rect 400956 489812 401008 489864
rect 518164 484372 518216 484424
rect 580172 484372 580224 484424
rect 361764 480224 361816 480276
rect 364984 480224 365036 480276
rect 400956 476756 401008 476808
rect 402244 476756 402296 476808
rect 518256 470568 518308 470620
rect 579988 470568 580040 470620
rect 402244 469820 402296 469872
rect 406016 469820 406068 469872
rect 361764 469208 361816 469260
rect 418988 469208 419040 469260
rect 406016 465060 406068 465112
rect 409144 464992 409196 465044
rect 514116 464380 514168 464432
rect 542360 464380 542412 464432
rect 450084 464312 450136 464364
rect 525800 464312 525852 464364
rect 494704 462476 494756 462528
rect 527640 462476 527692 462528
rect 436100 462408 436152 462460
rect 554136 462408 554188 462460
rect 433248 462340 433300 462392
rect 551192 462340 551244 462392
rect 480168 461592 480220 461644
rect 521752 461592 521804 461644
rect 450176 460912 450228 460964
rect 524420 460912 524472 460964
rect 361764 458192 361816 458244
rect 381636 458192 381688 458244
rect 409144 458124 409196 458176
rect 409880 458124 409932 458176
rect 449808 457444 449860 457496
rect 488540 457444 488592 457496
rect 473728 456764 473780 456816
rect 480168 456764 480220 456816
rect 488264 456016 488316 456068
rect 494704 456016 494756 456068
rect 450636 455472 450688 455524
rect 480996 455472 481048 455524
rect 409880 455404 409932 455456
rect 423588 455404 423640 455456
rect 473728 455404 473780 455456
rect 414388 455336 414440 455388
rect 450268 454792 450320 454844
rect 481732 454792 481784 454844
rect 449716 454724 449768 454776
rect 484400 454724 484452 454776
rect 449624 454656 449676 454708
rect 487160 454656 487212 454708
rect 414388 453296 414440 453348
rect 416688 453296 416740 453348
rect 416688 447924 416740 447976
rect 419080 447924 419132 447976
rect 422484 447516 422536 447568
rect 423588 447516 423640 447568
rect 432420 447516 432472 447568
rect 433248 447516 433300 447568
rect 361580 447176 361632 447228
rect 363788 447176 363840 447228
rect 433248 447176 433300 447228
rect 444196 447176 444248 447228
rect 423588 447108 423640 447160
rect 445576 447108 445628 447160
rect 436100 445680 436152 445732
rect 437388 445680 437440 445732
rect 427728 444524 427780 444576
rect 446220 444524 446272 444576
rect 437296 444456 437348 444508
rect 444380 444456 444432 444508
rect 442632 444388 442684 444440
rect 444104 444388 444156 444440
rect 444196 444320 444248 444372
rect 447232 444320 447284 444372
rect 456892 429836 456944 429888
rect 474280 429836 474332 429888
rect 480904 429156 480956 429208
rect 482284 429156 482336 429208
rect 483664 429156 483716 429208
rect 484952 429156 485004 429208
rect 486424 429156 486476 429208
rect 487620 429156 487672 429208
rect 457536 428408 457588 428460
rect 471612 428408 471664 428460
rect 502524 424328 502576 424380
rect 557540 424328 557592 424380
rect 529204 423580 529256 423632
rect 530216 423580 530268 423632
rect 530584 423580 530636 423632
rect 532792 423580 532844 423632
rect 511448 423512 511500 423564
rect 523776 423512 523828 423564
rect 522304 423444 522356 423496
rect 549536 423444 549588 423496
rect 502984 423376 503036 423428
rect 522488 423376 522540 423428
rect 523684 423376 523736 423428
rect 552112 423376 552164 423428
rect 485780 423308 485832 423360
rect 526352 423308 526404 423360
rect 526444 423308 526496 423360
rect 554688 423308 554740 423360
rect 487160 423240 487212 423292
rect 528928 423240 528980 423292
rect 488540 423172 488592 423224
rect 531504 423172 531556 423224
rect 496820 423104 496872 423156
rect 545672 423104 545724 423156
rect 498200 423036 498252 423088
rect 548248 423036 548300 423088
rect 499580 422968 499632 423020
rect 550824 422968 550876 423020
rect 501052 422900 501104 422952
rect 553400 422900 553452 422952
rect 483020 421540 483072 421592
rect 521200 421540 521252 421592
rect 419080 420588 419132 420640
rect 423956 420588 424008 420640
rect 494060 420180 494112 420232
rect 541808 420180 541860 420232
rect 362316 418752 362368 418804
rect 440884 418752 440936 418804
rect 421472 417732 421524 417784
rect 503720 417732 503772 417784
rect 425336 417664 425388 417716
rect 507860 417664 507912 417716
rect 424048 417596 424100 417648
rect 506480 417596 506532 417648
rect 424692 417528 424744 417580
rect 506572 417528 506624 417580
rect 422116 417460 422168 417512
rect 503996 417460 504048 417512
rect 425980 417392 426032 417444
rect 507952 417392 508004 417444
rect 423956 416780 424008 416832
rect 428464 416780 428516 416832
rect 362224 416032 362276 416084
rect 436744 416032 436796 416084
rect 361580 413992 361632 414044
rect 439504 413992 439556 414044
rect 428464 411272 428516 411324
rect 431224 411272 431276 411324
rect 511356 404336 511408 404388
rect 580172 404336 580224 404388
rect 361580 402976 361632 403028
rect 442264 402976 442316 403028
rect 497464 400868 497516 400920
rect 546500 400868 546552 400920
rect 431224 400120 431276 400172
rect 432604 400120 432656 400172
rect 494152 399440 494204 399492
rect 539600 399440 539652 399492
rect 459928 398080 459980 398132
rect 483664 398080 483716 398132
rect 492680 398080 492732 398132
rect 538220 398080 538272 398132
rect 458456 396720 458508 396772
rect 478880 396720 478932 396772
rect 492772 396720 492824 396772
rect 536840 396720 536892 396772
rect 458180 395292 458232 395344
rect 476120 395292 476172 395344
rect 491576 395292 491628 395344
rect 535460 395292 535512 395344
rect 465540 393932 465592 393984
rect 490012 393932 490064 393984
rect 491300 393932 491352 393984
rect 534172 393932 534224 393984
rect 496452 392640 496504 392692
rect 543740 392640 543792 392692
rect 422392 392572 422444 392624
rect 506020 392572 506072 392624
rect 361580 391960 361632 392012
rect 440976 391960 441028 392012
rect 459652 391280 459704 391332
rect 480904 391280 480956 391332
rect 495716 391280 495768 391332
rect 542360 391280 542412 391332
rect 422300 391212 422352 391264
rect 505284 391212 505336 391264
rect 461124 389784 461176 389836
rect 486424 389784 486476 389836
rect 490564 389784 490616 389836
rect 534080 389784 534132 389836
rect 449900 389240 449952 389292
rect 450728 389240 450780 389292
rect 465080 389240 465132 389292
rect 465908 389240 465960 389292
rect 492680 389240 492732 389292
rect 493140 389240 493192 389292
rect 494060 389240 494112 389292
rect 494612 389240 494664 389292
rect 453764 389104 453816 389156
rect 454684 389104 454736 389156
rect 461676 389104 461728 389156
rect 462596 389104 462648 389156
rect 464344 389104 464396 389156
rect 469220 389104 469272 389156
rect 461860 389036 461912 389088
rect 465540 389036 465592 389088
rect 483940 388968 483992 389020
rect 502984 388968 503036 389020
rect 468484 388900 468536 388952
rect 475108 388900 475160 388952
rect 499396 388900 499448 388952
rect 522304 388900 522356 388952
rect 456708 388832 456760 388884
rect 457536 388832 457588 388884
rect 468668 388832 468720 388884
rect 480996 388832 481048 388884
rect 500868 388832 500920 388884
rect 523684 388832 523736 388884
rect 468576 388764 468628 388816
rect 478052 388764 478104 388816
rect 502340 388764 502392 388816
rect 526444 388764 526496 388816
rect 467104 388696 467156 388748
rect 480260 388696 480312 388748
rect 484676 388696 484728 388748
rect 511448 388696 511500 388748
rect 467196 388628 467248 388680
rect 481732 388628 481784 388680
rect 485412 388628 485464 388680
rect 524420 388628 524472 388680
rect 461584 388560 461636 388612
rect 476580 388560 476632 388612
rect 486884 388560 486936 388612
rect 527180 388560 527232 388612
rect 461768 388492 461820 388544
rect 478788 388492 478840 388544
rect 488356 388492 488408 388544
rect 529204 388492 529256 388544
rect 462964 388424 463016 388476
rect 482468 388424 482520 388476
rect 489828 388424 489880 388476
rect 530584 388424 530636 388476
rect 447876 387132 447928 387184
rect 457444 387132 457496 387184
rect 448980 387064 449032 387116
rect 491116 387064 491168 387116
rect 445576 386520 445628 386572
rect 553952 386520 554004 386572
rect 381544 386452 381596 386504
rect 512184 386452 512236 386504
rect 370504 386384 370556 386436
rect 512000 386384 512052 386436
rect 448428 385976 448480 386028
rect 451924 385976 451976 386028
rect 447784 385364 447836 385416
rect 453304 385364 453356 385416
rect 450360 385092 450412 385144
rect 563428 385092 563480 385144
rect 370596 385024 370648 385076
rect 512092 385024 512144 385076
rect 512736 383732 512788 383784
rect 534724 383732 534776 383784
rect 513288 383664 513340 383716
rect 547144 383664 547196 383716
rect 378784 383596 378836 383648
rect 447324 383596 447376 383648
rect 382924 383528 382976 383580
rect 447140 383528 447192 383580
rect 512460 382984 512512 383036
rect 518348 382984 518400 383036
rect 513012 382440 513064 382492
rect 519636 382440 519688 382492
rect 512276 382304 512328 382356
rect 515588 382304 515640 382356
rect 376024 382168 376076 382220
rect 447324 382168 447376 382220
rect 400864 382100 400916 382152
rect 447140 382100 447192 382152
rect 361580 380876 361632 380928
rect 442356 380876 442408 380928
rect 513288 380876 513340 380928
rect 548524 380876 548576 380928
rect 374644 380808 374696 380860
rect 447508 380808 447560 380860
rect 403624 380740 403676 380792
rect 447140 380740 447192 380792
rect 406384 380672 406436 380724
rect 447324 380672 447376 380724
rect 512000 380400 512052 380452
rect 512368 380400 512420 380452
rect 512000 380264 512052 380316
rect 514208 380264 514260 380316
rect 513288 379516 513340 379568
rect 544384 379516 544436 379568
rect 370688 379448 370740 379500
rect 447508 379448 447560 379500
rect 371884 379380 371936 379432
rect 447140 379380 447192 379432
rect 512184 378292 512236 378344
rect 522304 378292 522356 378344
rect 513288 378224 513340 378276
rect 548616 378224 548668 378276
rect 516784 378156 516836 378208
rect 580172 378156 580224 378208
rect 363604 378088 363656 378140
rect 447324 378088 447376 378140
rect 367744 378020 367796 378072
rect 447140 378020 447192 378072
rect 432604 377952 432656 378004
rect 436836 377952 436888 378004
rect 512828 377408 512880 377460
rect 549904 377408 549956 377460
rect 513196 376728 513248 376780
rect 516968 376728 517020 376780
rect 363696 376660 363748 376712
rect 447140 376660 447192 376712
rect 407764 376592 407816 376644
rect 447324 376592 447376 376644
rect 512460 375980 512512 376032
rect 547236 375980 547288 376032
rect 513288 375640 513340 375692
rect 520280 375640 520332 375692
rect 410524 375300 410576 375352
rect 447140 375300 447192 375352
rect 411904 375232 411956 375284
rect 447324 375232 447376 375284
rect 512460 374144 512512 374196
rect 515680 374144 515732 374196
rect 414664 373940 414716 373992
rect 447140 373940 447192 373992
rect 416044 373872 416096 373924
rect 447324 373872 447376 373924
rect 512644 373736 512696 373788
rect 516232 373736 516284 373788
rect 513288 372716 513340 372768
rect 521660 372716 521712 372768
rect 512092 372648 512144 372700
rect 514852 372648 514904 372700
rect 364984 372512 365036 372564
rect 447324 372512 447376 372564
rect 417516 372444 417568 372496
rect 447140 372444 447192 372496
rect 512460 371764 512512 371816
rect 516324 371764 516376 371816
rect 381636 371152 381688 371204
rect 447324 371152 447376 371204
rect 418988 371084 419040 371136
rect 447140 371084 447192 371136
rect 513288 370064 513340 370116
rect 520372 370064 520424 370116
rect 512736 369928 512788 369980
rect 516140 369928 516192 369980
rect 361580 369860 361632 369912
rect 429200 369860 429252 369912
rect 363788 369792 363840 369844
rect 447140 369792 447192 369844
rect 436744 369724 436796 369776
rect 447324 369724 447376 369776
rect 513288 368500 513340 368552
rect 520464 368500 520516 368552
rect 439504 368432 439556 368484
rect 447324 368432 447376 368484
rect 440884 368364 440936 368416
rect 447140 368364 447192 368416
rect 512644 367344 512696 367396
rect 518992 367344 519044 367396
rect 512000 367208 512052 367260
rect 514944 367208 514996 367260
rect 440976 367004 441028 367056
rect 447140 367004 447192 367056
rect 442264 366936 442316 366988
rect 447324 366936 447376 366988
rect 513288 365848 513340 365900
rect 520556 365848 520608 365900
rect 513196 365712 513248 365764
rect 518900 365712 518952 365764
rect 429200 365644 429252 365696
rect 447140 365644 447192 365696
rect 442356 365576 442408 365628
rect 447324 365576 447376 365628
rect 512000 364488 512052 364540
rect 514300 364488 514352 364540
rect 513288 364352 513340 364404
rect 523040 364352 523092 364404
rect 569224 364352 569276 364404
rect 580172 364352 580224 364404
rect 512092 363536 512144 363588
rect 513656 363536 513708 363588
rect 437020 362992 437072 363044
rect 447140 362992 447192 363044
rect 432604 362924 432656 362976
rect 447324 362924 447376 362976
rect 512368 362312 512420 362364
rect 513748 362312 513800 362364
rect 513196 361768 513248 361820
rect 519084 361768 519136 361820
rect 442264 361632 442316 361684
rect 447324 361632 447376 361684
rect 439688 361564 439740 361616
rect 447140 361564 447192 361616
rect 513288 361564 513340 361616
rect 521752 361564 521804 361616
rect 522304 360816 522356 360868
rect 550640 360816 550692 360868
rect 512828 360408 512880 360460
rect 519176 360408 519228 360460
rect 513288 360340 513340 360392
rect 523132 360340 523184 360392
rect 442356 360272 442408 360324
rect 447324 360272 447376 360324
rect 512368 360272 512420 360324
rect 515128 360272 515180 360324
rect 435456 360204 435508 360256
rect 447140 360204 447192 360256
rect 548616 360136 548668 360188
rect 552020 360136 552072 360188
rect 548524 359048 548576 359100
rect 558184 359048 558236 359100
rect 544384 358980 544436 359032
rect 553768 358980 553820 359032
rect 512368 358912 512420 358964
rect 513840 358912 513892 358964
rect 547144 358912 547196 358964
rect 565544 358912 565596 358964
rect 441068 358844 441120 358896
rect 447324 358844 447376 358896
rect 512920 358844 512972 358896
rect 519268 358844 519320 358896
rect 534724 358844 534776 358896
rect 567016 358844 567068 358896
rect 436928 358776 436980 358828
rect 447140 358776 447192 358828
rect 514208 358776 514260 358828
rect 555240 358776 555292 358828
rect 549904 358708 549956 358760
rect 556712 358708 556764 358760
rect 519636 358640 519688 358692
rect 564072 358640 564124 358692
rect 518348 358572 518400 358624
rect 562600 358572 562652 358624
rect 547236 358504 547288 358556
rect 559656 358504 559708 358556
rect 515588 358436 515640 358488
rect 561128 358436 561180 358488
rect 512920 356192 512972 356244
rect 516508 356192 516560 356244
rect 513288 355104 513340 355156
rect 517520 355104 517572 355156
rect 445576 354220 445628 354272
rect 447324 354220 447376 354272
rect 512368 353608 512420 353660
rect 515036 353608 515088 353660
rect 512828 353064 512880 353116
rect 517612 353064 517664 353116
rect 512368 352384 512420 352436
rect 515220 352384 515272 352436
rect 511448 352112 511500 352164
rect 580172 352112 580224 352164
rect 513288 351976 513340 352028
rect 519360 351976 519412 352028
rect 512368 350888 512420 350940
rect 515312 350888 515364 350940
rect 513012 350616 513064 350668
rect 517704 350616 517756 350668
rect 405740 350548 405792 350600
rect 447140 350548 447192 350600
rect 513196 349528 513248 349580
rect 520648 349528 520700 349580
rect 512368 349256 512420 349308
rect 513932 349256 513984 349308
rect 513012 349188 513064 349240
rect 516600 349188 516652 349240
rect 513012 348032 513064 348084
rect 517796 348032 517848 348084
rect 361764 347760 361816 347812
rect 402244 347760 402296 347812
rect 362224 347692 362276 347744
rect 447140 347692 447192 347744
rect 513288 346672 513340 346724
rect 519452 346672 519504 346724
rect 513104 346536 513156 346588
rect 516876 346536 516928 346588
rect 446220 344904 446272 344956
rect 448428 344904 448480 344956
rect 432696 344292 432748 344344
rect 442264 344292 442316 344344
rect 447324 344224 447376 344276
rect 447508 344224 447560 344276
rect 436836 343884 436888 343936
rect 439136 343884 439188 343936
rect 512644 343680 512696 343732
rect 520740 343680 520792 343732
rect 513012 343136 513064 343188
rect 517888 343136 517940 343188
rect 402244 342864 402296 342916
rect 447508 342864 447560 342916
rect 513288 342252 513340 342304
rect 521844 342252 521896 342304
rect 447232 342184 447284 342236
rect 447600 342184 447652 342236
rect 513012 341096 513064 341148
rect 516692 341096 516744 341148
rect 418160 340960 418212 341012
rect 447140 340960 447192 341012
rect 513288 340960 513340 341012
rect 517980 340960 518032 341012
rect 361764 340892 361816 340944
rect 447232 340892 447284 340944
rect 513288 339600 513340 339652
rect 519636 339600 519688 339652
rect 443736 339532 443788 339584
rect 447232 339532 447284 339584
rect 513104 339532 513156 339584
rect 518072 339532 518124 339584
rect 399484 339464 399536 339516
rect 447140 339464 447192 339516
rect 513196 339464 513248 339516
rect 521936 339464 521988 339516
rect 512644 338240 512696 338292
rect 520832 338240 520884 338292
rect 436836 338172 436888 338224
rect 447140 338172 447192 338224
rect 385684 338104 385736 338156
rect 447232 338104 447284 338156
rect 512828 338104 512880 338156
rect 522028 338104 522080 338156
rect 439136 338036 439188 338088
rect 441252 338036 441304 338088
rect 362224 337356 362276 337408
rect 418160 337356 418212 337408
rect 513288 337016 513340 337068
rect 518348 337016 518400 337068
rect 513288 336880 513340 336932
rect 519728 336880 519780 336932
rect 420460 336812 420512 336864
rect 429844 336812 429896 336864
rect 431224 336812 431276 336864
rect 447232 336812 447284 336864
rect 416780 336744 416832 336796
rect 439872 336744 439924 336796
rect 440976 336744 441028 336796
rect 447140 336744 447192 336796
rect 418804 336200 418856 336252
rect 438124 336200 438176 336252
rect 418896 336132 418948 336184
rect 441344 336132 441396 336184
rect 412640 336064 412692 336116
rect 449440 336064 449492 336116
rect 397460 335996 397512 336048
rect 441160 335996 441212 336048
rect 413100 335384 413152 335436
rect 435548 335384 435600 335436
rect 439780 335384 439832 335436
rect 447140 335384 447192 335436
rect 409420 335316 409472 335368
rect 431316 335316 431368 335368
rect 435364 335316 435416 335368
rect 447232 335316 447284 335368
rect 420368 335044 420420 335096
rect 420828 335044 420880 335096
rect 443828 335044 443880 335096
rect 443920 334976 443972 335028
rect 420736 334908 420788 334960
rect 446220 334908 446272 334960
rect 417424 334840 417476 334892
rect 444012 334840 444064 334892
rect 420184 334772 420236 334824
rect 449072 334772 449124 334824
rect 420552 334704 420604 334756
rect 450452 334704 450504 334756
rect 420644 334636 420696 334688
rect 450728 334636 450780 334688
rect 420276 334568 420328 334620
rect 450636 334568 450688 334620
rect 428096 334364 428148 334416
rect 512736 334296 512788 334348
rect 514760 334296 514812 334348
rect 447416 334092 447468 334144
rect 442264 334024 442316 334076
rect 447508 334024 447560 334076
rect 363604 333956 363656 334008
rect 447232 333956 447284 334008
rect 439504 332800 439556 332852
rect 447140 332800 447192 332852
rect 436744 332664 436796 332716
rect 432972 332596 433024 332648
rect 437020 332596 437072 332648
rect 447416 332732 447468 332784
rect 443644 332596 443696 332648
rect 447232 332596 447284 332648
rect 512920 331440 512972 331492
rect 516416 331440 516468 331492
rect 444104 331304 444156 331356
rect 444288 331304 444340 331356
rect 447232 331304 447284 331356
rect 432788 331236 432840 331288
rect 439688 331236 439740 331288
rect 440884 331236 440936 331288
rect 447140 331236 447192 331288
rect 442908 330556 442960 330608
rect 444380 330556 444432 330608
rect 447140 330556 447192 330608
rect 438768 330488 438820 330540
rect 447600 330488 447652 330540
rect 432604 330012 432656 330064
rect 435456 330012 435508 330064
rect 431868 329060 431920 329112
rect 447416 329060 447468 329112
rect 436008 328448 436060 328500
rect 447140 328448 447192 328500
rect 429200 328380 429252 328432
rect 448244 328380 448296 328432
rect 429844 327020 429896 327072
rect 447416 327020 447468 327072
rect 448152 327020 448204 327072
rect 439872 326952 439924 327004
rect 447968 326952 448020 327004
rect 435548 325524 435600 325576
rect 448060 325524 448112 325576
rect 431316 324912 431368 324964
rect 448336 324912 448388 324964
rect 449532 324912 449584 324964
rect 432696 323552 432748 323604
rect 442356 323552 442408 323604
rect 509700 323416 509752 323468
rect 510252 323416 510304 323468
rect 507492 322668 507544 322720
rect 510068 322668 510120 322720
rect 507584 322600 507636 322652
rect 509608 322600 509660 322652
rect 507400 322532 507452 322584
rect 510160 322532 510212 322584
rect 507308 322464 507360 322516
rect 509976 322464 510028 322516
rect 450452 322328 450504 322380
rect 463516 322396 463568 322448
rect 507124 322396 507176 322448
rect 511172 322396 511224 322448
rect 441252 322260 441304 322312
rect 464896 322328 464948 322380
rect 459652 322260 459704 322312
rect 463516 322260 463568 322312
rect 443920 322192 443972 322244
rect 463240 322192 463292 322244
rect 502156 322192 502208 322244
rect 580448 322192 580500 322244
rect 449256 322124 449308 322176
rect 471796 322124 471848 322176
rect 450728 322056 450780 322108
rect 484216 322056 484268 322108
rect 445668 321988 445720 322040
rect 481180 321988 481232 322040
rect 446220 321920 446272 321972
rect 483940 321920 483992 321972
rect 449072 321852 449124 321904
rect 474096 321852 474148 321904
rect 479616 321852 479668 321904
rect 518164 321852 518216 321904
rect 444012 321784 444064 321836
rect 463884 321784 463936 321836
rect 469128 321784 469180 321836
rect 518256 321784 518308 321836
rect 459192 321716 459244 321768
rect 515496 321716 515548 321768
rect 449164 321648 449216 321700
rect 460572 321648 460624 321700
rect 459744 321580 459796 321632
rect 567844 321648 567896 321700
rect 463516 321580 463568 321632
rect 580264 321580 580316 321632
rect 458916 321512 458968 321564
rect 580540 321512 580592 321564
rect 445024 321444 445076 321496
rect 460848 321444 460900 321496
rect 470232 321444 470284 321496
rect 576124 321444 576176 321496
rect 450544 321376 450596 321428
rect 461400 321376 461452 321428
rect 469956 321376 470008 321428
rect 574744 321376 574796 321428
rect 445484 321308 445536 321360
rect 462504 321308 462556 321360
rect 468576 321308 468628 321360
rect 569224 321308 569276 321360
rect 480720 321240 480772 321292
rect 573364 321240 573416 321292
rect 458088 321172 458140 321224
rect 511448 321172 511500 321224
rect 458364 321104 458416 321156
rect 511356 321104 511408 321156
rect 446404 321036 446456 321088
rect 471336 321036 471388 321088
rect 479064 321036 479116 321088
rect 516784 321036 516836 321088
rect 450636 320968 450688 321020
rect 484584 320968 484636 321020
rect 447048 320900 447100 320952
rect 473544 320900 473596 320952
rect 496820 320900 496872 320952
rect 580724 320900 580776 320952
rect 461860 320832 461912 320884
rect 580632 320832 580684 320884
rect 441160 320764 441212 320816
rect 481548 320764 481600 320816
rect 438124 320696 438176 320748
rect 472440 320696 472492 320748
rect 446956 320628 447008 320680
rect 473820 320628 473872 320680
rect 445116 320560 445168 320612
rect 461952 320560 462004 320612
rect 441344 320492 441396 320544
rect 481824 320492 481876 320544
rect 458640 320084 458692 320136
rect 461860 320084 461912 320136
rect 464896 320084 464948 320136
rect 474372 320084 474424 320136
rect 479340 320084 479392 320136
rect 496820 320084 496872 320136
rect 449348 320016 449400 320068
rect 461124 320016 461176 320068
rect 469680 320016 469732 320068
rect 580356 320016 580408 320068
rect 444196 319948 444248 320000
rect 460296 319948 460348 320000
rect 478788 319948 478840 320000
rect 580172 319948 580224 320000
rect 470508 319880 470560 319932
rect 514116 319880 514168 319932
rect 449440 319812 449492 319864
rect 471060 319812 471112 319864
rect 480996 319812 481048 319864
rect 519544 319812 519596 319864
rect 443828 319744 443880 319796
rect 463056 319744 463108 319796
rect 480444 319744 480496 319796
rect 515404 319744 515456 319796
rect 445300 319676 445352 319728
rect 462780 319676 462832 319728
rect 479892 319676 479944 319728
rect 514024 319676 514076 319728
rect 458916 319608 458968 319660
rect 465540 319608 465592 319660
rect 469404 319608 469456 319660
rect 502156 319608 502208 319660
rect 459100 319540 459152 319592
rect 476028 319540 476080 319592
rect 480168 319540 480220 319592
rect 511264 319540 511316 319592
rect 460388 319472 460440 319524
rect 476304 319472 476356 319524
rect 498108 319472 498160 319524
rect 530676 319472 530728 319524
rect 456156 319404 456208 319456
rect 486516 319404 486568 319456
rect 502800 319404 502852 319456
rect 538864 319404 538916 319456
rect 460296 319336 460348 319388
rect 465816 319336 465868 319388
rect 498660 319336 498712 319388
rect 530584 319336 530636 319388
rect 445392 319268 445444 319320
rect 473268 319268 473320 319320
rect 487252 319268 487304 319320
rect 487804 319268 487856 319320
rect 494428 319268 494480 319320
rect 494704 319268 494756 319320
rect 455512 319200 455564 319252
rect 456340 319200 456392 319252
rect 466552 319200 466604 319252
rect 467380 319200 467432 319252
rect 468852 319200 468904 319252
rect 580816 319200 580868 319252
rect 446680 319132 446732 319184
rect 472992 319132 473044 319184
rect 474832 319132 474884 319184
rect 475108 319132 475160 319184
rect 476212 319132 476264 319184
rect 477316 319132 477368 319184
rect 477592 319132 477644 319184
rect 478144 319132 478196 319184
rect 446864 319064 446916 319116
rect 483480 319064 483532 319116
rect 485872 319064 485924 319116
rect 486976 319064 487028 319116
rect 488908 319064 488960 319116
rect 489736 319064 489788 319116
rect 493048 319064 493100 319116
rect 493600 319064 493652 319116
rect 495808 319064 495860 319116
rect 496360 319064 496412 319116
rect 496912 319064 496964 319116
rect 497188 319064 497240 319116
rect 498568 319064 498620 319116
rect 499396 319064 499448 319116
rect 499672 319064 499724 319116
rect 500776 319064 500828 319116
rect 501052 319064 501104 319116
rect 501328 319064 501380 319116
rect 502432 319064 502484 319116
rect 503536 319064 503588 319116
rect 446496 318996 446548 319048
rect 482100 318996 482152 319048
rect 492772 318996 492824 319048
rect 493876 318996 493928 319048
rect 495532 318996 495584 319048
rect 496636 318996 496688 319048
rect 498292 318996 498344 319048
rect 499120 318996 499172 319048
rect 455604 318928 455656 318980
rect 456064 318928 456116 318980
rect 456892 318928 456944 318980
rect 457444 318928 457496 318980
rect 466828 318928 466880 318980
rect 467104 318928 467156 318980
rect 476488 318928 476540 318980
rect 476764 318928 476816 318980
rect 491944 318928 491996 318980
rect 492496 318928 492548 318980
rect 497188 318928 497240 318980
rect 497740 318928 497792 318980
rect 455420 318860 455472 318912
rect 456616 318860 456668 318912
rect 442816 318724 442868 318776
rect 470784 318724 470836 318776
rect 478512 318724 478564 318776
rect 479524 318724 479576 318776
rect 457812 318316 457864 318368
rect 461584 318316 461636 318368
rect 459192 318248 459244 318300
rect 491484 318248 491536 318300
rect 501696 318248 501748 318300
rect 540336 318248 540388 318300
rect 452108 318180 452160 318232
rect 495624 318180 495676 318232
rect 496176 318180 496228 318232
rect 540980 318180 541032 318232
rect 458824 318112 458876 318164
rect 512276 318112 512328 318164
rect 448244 318044 448296 318096
rect 455236 318044 455288 318096
rect 456064 318044 456116 318096
rect 512460 318044 512512 318096
rect 456340 317364 456392 317416
rect 475752 317364 475804 317416
rect 456524 317296 456576 317348
rect 486240 317296 486292 317348
rect 453580 317228 453632 317280
rect 485688 317228 485740 317280
rect 500316 317228 500368 317280
rect 539692 317228 539744 317280
rect 454776 317160 454828 317212
rect 491576 317160 491628 317212
rect 502524 317160 502576 317212
rect 543096 317160 543148 317212
rect 453396 317092 453448 317144
rect 485964 317092 486016 317144
rect 487344 317092 487396 317144
rect 529940 317092 529992 317144
rect 455052 317024 455104 317076
rect 509884 317024 509936 317076
rect 456248 316956 456300 317008
rect 511080 316956 511132 317008
rect 454868 316888 454920 316940
rect 510252 316888 510304 316940
rect 450728 316820 450780 316872
rect 509700 316820 509752 316872
rect 450636 316752 450688 316804
rect 512368 316752 512420 316804
rect 450544 316684 450596 316736
rect 514760 316684 514812 316736
rect 456432 316616 456484 316668
rect 475476 316616 475528 316668
rect 453488 316548 453540 316600
rect 464988 316548 465040 316600
rect 459008 316480 459060 316532
rect 465264 316480 465316 316532
rect 361764 315936 361816 315988
rect 399484 315936 399536 315988
rect 452016 315324 452068 315376
rect 494152 315324 494204 315376
rect 501144 315324 501196 315376
rect 541072 315324 541124 315376
rect 455696 315256 455748 315308
rect 562324 315256 562376 315308
rect 451096 314236 451148 314288
rect 464712 314236 464764 314288
rect 451004 314168 451056 314220
rect 475016 314168 475068 314220
rect 457444 314100 457496 314152
rect 485320 314100 485372 314152
rect 502984 314100 503036 314152
rect 538956 314100 539008 314152
rect 452200 314032 452252 314084
rect 494980 314032 495032 314084
rect 501328 314032 501380 314084
rect 543004 314032 543056 314084
rect 450820 313964 450872 314016
rect 513380 313964 513432 314016
rect 450912 313896 450964 313948
rect 474832 313896 474884 313948
rect 476764 313896 476816 313948
rect 548524 313896 548576 313948
rect 482284 313284 482336 313336
rect 484492 313284 484544 313336
rect 468208 313216 468260 313268
rect 580172 313216 580224 313268
rect 466644 312536 466696 312588
rect 544384 312536 544436 312588
rect 451924 311176 451976 311228
rect 489460 311176 489512 311228
rect 502708 311176 502760 311228
rect 542728 311176 542780 311228
rect 432604 311108 432656 311160
rect 441068 311108 441120 311160
rect 477684 311108 477736 311160
rect 547144 311108 547196 311160
rect 461676 310904 461728 310956
rect 463792 310904 463844 310956
rect 495532 309816 495584 309868
rect 539600 309816 539652 309868
rect 453672 309748 453724 309800
rect 490840 309748 490892 309800
rect 497004 309748 497056 309800
rect 542912 309748 542964 309800
rect 453764 308456 453816 308508
rect 491116 308456 491168 308508
rect 487804 308388 487856 308440
rect 529204 308388 529256 308440
rect 432420 307708 432472 307760
rect 436928 307708 436980 307760
rect 471244 307708 471296 307760
rect 473728 307708 473780 307760
rect 487528 307164 487580 307216
rect 530032 307164 530084 307216
rect 449624 307096 449676 307148
rect 536840 307096 536892 307148
rect 465724 307028 465776 307080
rect 566464 307028 566516 307080
rect 409236 306280 409288 306332
rect 454960 306280 455012 306332
rect 409144 306212 409196 306264
rect 455052 306212 455104 306264
rect 406752 306144 406804 306196
rect 454868 306144 454920 306196
rect 457536 306144 457588 306196
rect 493048 306144 493100 306196
rect 400864 306076 400916 306128
rect 465448 306076 465500 306128
rect 476488 306076 476540 306128
rect 565084 306076 565136 306128
rect 406476 306008 406528 306060
rect 510988 306008 511040 306060
rect 403992 305940 404044 305992
rect 510896 305940 510948 305992
rect 403624 305872 403676 305924
rect 510804 305872 510856 305924
rect 406568 305804 406620 305856
rect 513932 305804 513984 305856
rect 406660 305736 406712 305788
rect 515220 305736 515272 305788
rect 406384 305668 406436 305720
rect 515312 305668 515364 305720
rect 359464 305600 359516 305652
rect 512552 305600 512604 305652
rect 447784 305532 447836 305584
rect 464068 305532 464120 305584
rect 3608 304988 3660 305040
rect 4804 304988 4856 305040
rect 361764 304920 361816 304972
rect 443736 304920 443788 304972
rect 446404 304444 446456 304496
rect 461676 304444 461728 304496
rect 455604 304376 455656 304428
rect 563704 304376 563756 304428
rect 362224 304308 362276 304360
rect 512828 304308 512880 304360
rect 360844 304240 360896 304292
rect 512184 304240 512236 304292
rect 401048 303560 401100 303612
rect 510620 303560 510672 303612
rect 403808 303492 403860 303544
rect 513840 303492 513892 303544
rect 398380 303424 398432 303476
rect 509332 303424 509384 303476
rect 401232 303356 401284 303408
rect 513656 303356 513708 303408
rect 400956 303288 401008 303340
rect 513748 303288 513800 303340
rect 401324 303220 401376 303272
rect 515128 303220 515180 303272
rect 401140 303152 401192 303204
rect 514944 303152 514996 303204
rect 398288 303084 398340 303136
rect 513472 303084 513524 303136
rect 398196 303016 398248 303068
rect 516324 303016 516376 303068
rect 455512 302948 455564 303000
rect 574744 302948 574796 303000
rect 360936 302880 360988 302932
rect 512644 302880 512696 302932
rect 403716 302812 403768 302864
rect 509424 302812 509476 302864
rect 396724 302744 396776 302796
rect 485872 302744 485924 302796
rect 455420 301452 455472 301504
rect 576124 301452 576176 301504
rect 456984 300704 457036 300756
rect 537484 300704 537536 300756
rect 398104 300636 398156 300688
rect 516232 300636 516284 300688
rect 395620 300568 395672 300620
rect 517980 300568 518032 300620
rect 395804 300500 395856 300552
rect 518348 300500 518400 300552
rect 395436 300432 395488 300484
rect 518072 300432 518124 300484
rect 392768 300364 392820 300416
rect 516600 300364 516652 300416
rect 392952 300296 393004 300348
rect 516876 300296 516928 300348
rect 393044 300228 393096 300280
rect 517796 300228 517848 300280
rect 392676 300160 392728 300212
rect 517888 300160 517940 300212
rect 361028 300092 361080 300144
rect 512000 300092 512052 300144
rect 461584 299412 461636 299464
rect 580172 299412 580224 299464
rect 457168 298052 457220 298104
rect 578884 298052 578936 298104
rect 392860 297984 392912 298036
rect 517704 297984 517756 298036
rect 387248 297916 387300 297968
rect 514300 297916 514352 297968
rect 389916 297848 389968 297900
rect 516508 297848 516560 297900
rect 390192 297780 390244 297832
rect 517612 297780 517664 297832
rect 390100 297712 390152 297764
rect 519268 297712 519320 297764
rect 387524 297644 387576 297696
rect 519176 297644 519228 297696
rect 387340 297576 387392 297628
rect 519084 297576 519136 297628
rect 387156 297508 387208 297560
rect 518992 297508 519044 297560
rect 387064 297440 387116 297492
rect 520556 297440 520608 297492
rect 361120 297372 361172 297424
rect 512092 297372 512144 297424
rect 390008 297304 390060 297356
rect 511540 297304 511592 297356
rect 390284 297236 390336 297288
rect 507584 297236 507636 297288
rect 456892 295944 456944 295996
rect 571984 295944 572036 295996
rect 384304 295264 384356 295316
rect 507400 295264 507452 295316
rect 381912 295196 381964 295248
rect 507492 295196 507544 295248
rect 384580 295128 384632 295180
rect 514852 295128 514904 295180
rect 384396 295060 384448 295112
rect 515680 295060 515732 295112
rect 387432 294992 387484 295044
rect 520464 294992 520516 295044
rect 384488 294924 384540 294976
rect 520372 294924 520424 294976
rect 382004 294856 382056 294908
rect 519728 294856 519780 294908
rect 378876 294788 378928 294840
rect 516692 294788 516744 294840
rect 381728 294720 381780 294772
rect 520280 294720 520332 294772
rect 378968 294652 379020 294704
rect 519636 294652 519688 294704
rect 379060 294584 379112 294636
rect 520832 294584 520884 294636
rect 476212 294516 476264 294568
rect 573364 294516 573416 294568
rect 361764 293904 361816 293956
rect 385684 293904 385736 293956
rect 467104 293224 467156 293276
rect 559564 293224 559616 293276
rect 3608 292544 3660 292596
rect 19984 292544 20036 292596
rect 373448 292476 373500 292528
rect 513564 292476 513616 292528
rect 379152 292408 379204 292460
rect 519452 292408 519504 292460
rect 376484 292340 376536 292392
rect 517520 292340 517572 292392
rect 379244 292272 379296 292324
rect 520740 292272 520792 292324
rect 376116 292204 376168 292256
rect 519360 292204 519412 292256
rect 376300 292136 376352 292188
rect 520648 292136 520700 292188
rect 370688 292068 370740 292120
rect 516140 292068 516192 292120
rect 370780 292000 370832 292052
rect 518900 292000 518952 292052
rect 373540 291932 373592 291984
rect 521752 291932 521804 291984
rect 373356 291864 373408 291916
rect 523040 291864 523092 291916
rect 373264 291796 373316 291848
rect 523132 291796 523184 291848
rect 376208 291728 376260 291780
rect 515036 291728 515088 291780
rect 466920 291660 466972 291712
rect 569224 291660 569276 291712
rect 399484 291592 399536 291644
rect 486148 291592 486200 291644
rect 477868 290436 477920 290488
rect 551284 290436 551336 290488
rect 439688 289620 439740 289672
rect 446404 289620 446456 289672
rect 477592 289620 477644 289672
rect 570604 289620 570656 289672
rect 405004 289552 405056 289604
rect 516416 289552 516468 289604
rect 368112 289484 368164 289536
rect 507124 289484 507176 289536
rect 368204 289416 368256 289468
rect 507308 289416 507360 289468
rect 367744 289348 367796 289400
rect 507216 289348 507268 289400
rect 370964 289280 371016 289332
rect 521660 289280 521712 289332
rect 368020 289212 368072 289264
rect 521844 289212 521896 289264
rect 367928 289144 367980 289196
rect 522028 289144 522080 289196
rect 367836 289076 367888 289128
rect 521936 289076 521988 289128
rect 465724 288396 465776 288448
rect 471244 288396 471296 288448
rect 476764 288396 476816 288448
rect 482284 288396 482336 288448
rect 445024 288328 445076 288380
rect 447784 288328 447836 288380
rect 487252 287648 487304 287700
rect 531320 287648 531372 287700
rect 453856 284996 453908 285048
rect 489184 284996 489236 285048
rect 376024 284928 376076 284980
rect 476580 284928 476632 284980
rect 498384 284928 498436 284980
rect 539876 284928 539928 284980
rect 452476 283568 452528 283620
rect 494520 283568 494572 283620
rect 361764 282820 361816 282872
rect 436836 282820 436888 282872
rect 455052 282208 455104 282260
rect 493324 282208 493376 282260
rect 466828 282140 466880 282192
rect 554044 282140 554096 282192
rect 457628 280780 457680 280832
rect 492864 280780 492916 280832
rect 502432 280780 502484 280832
rect 539048 280780 539100 280832
rect 459284 279488 459336 279540
rect 492220 279488 492272 279540
rect 453948 279420 454000 279472
rect 490564 279420 490616 279472
rect 500224 279420 500276 279472
rect 540152 279420 540204 279472
rect 460480 277992 460532 278044
rect 494704 277992 494756 278044
rect 499948 277992 500000 278044
rect 541440 277992 541492 278044
rect 454868 276632 454920 276684
rect 489000 276632 489052 276684
rect 499764 276632 499816 276684
rect 539968 276632 540020 276684
rect 459468 275340 459520 275392
rect 492772 275340 492824 275392
rect 452292 275272 452344 275324
rect 490012 275272 490064 275324
rect 498844 275272 498896 275324
rect 541256 275272 541308 275324
rect 460572 274048 460624 274100
rect 465724 274048 465776 274100
rect 455144 273980 455196 274032
rect 491944 273980 491996 274032
rect 498568 273980 498620 274032
rect 541348 273980 541400 274032
rect 456616 273912 456668 273964
rect 495900 273912 495952 273964
rect 497464 273912 497516 273964
rect 541164 273912 541216 273964
rect 479524 273164 479576 273216
rect 580172 273164 580224 273216
rect 457720 272552 457772 272604
rect 491668 272552 491720 272604
rect 457812 272484 457864 272536
rect 494428 272484 494480 272536
rect 501052 272484 501104 272536
rect 540244 272484 540296 272536
rect 361764 271804 361816 271856
rect 431224 271804 431276 271856
rect 459376 271260 459428 271312
rect 493140 271260 493192 271312
rect 454960 271192 455012 271244
rect 488632 271192 488684 271244
rect 498292 271192 498344 271244
rect 540060 271192 540112 271244
rect 453212 271124 453264 271176
rect 488908 271124 488960 271176
rect 499672 271124 499724 271176
rect 541532 271124 541584 271176
rect 503812 269968 503864 270020
rect 543740 269968 543792 270020
rect 456708 269900 456760 269952
rect 488080 269900 488132 269952
rect 497188 269900 497240 269952
rect 542820 269900 542872 269952
rect 467932 269832 467984 269884
rect 580264 269832 580316 269884
rect 359556 269764 359608 269816
rect 512736 269764 512788 269816
rect 481088 269288 481140 269340
rect 484768 269288 484820 269340
rect 445668 268540 445720 268592
rect 476764 268540 476816 268592
rect 447784 268472 447836 268524
rect 481088 268472 481140 268524
rect 452384 268404 452436 268456
rect 490288 268404 490340 268456
rect 496912 268404 496964 268456
rect 542636 268404 542688 268456
rect 466552 268336 466604 268388
rect 555424 268336 555476 268388
rect 435456 266976 435508 267028
rect 460572 266976 460624 267028
rect 3516 266364 3568 266416
rect 4896 266364 4948 266416
rect 447968 265616 448020 265668
rect 457904 265616 457956 265668
rect 420920 264256 420972 264308
rect 439688 264256 439740 264308
rect 422944 264188 422996 264240
rect 445668 264188 445720 264240
rect 449716 263508 449768 263560
rect 456800 263508 456852 263560
rect 431224 262828 431276 262880
rect 445024 262828 445076 262880
rect 411904 261468 411956 261520
rect 420920 261468 420972 261520
rect 361764 260788 361816 260840
rect 440976 260788 441028 260840
rect 401416 255960 401468 256012
rect 411904 255960 411956 256012
rect 428464 253920 428516 253972
rect 431224 253920 431276 253972
rect 361764 249704 361816 249756
rect 435364 249704 435416 249756
rect 449808 249704 449860 249756
rect 449992 249704 450044 249756
rect 449992 248412 450044 248464
rect 456800 248412 456852 248464
rect 571984 245556 572036 245608
rect 580172 245556 580224 245608
rect 398472 243176 398524 243228
rect 401416 243176 401468 243228
rect 3884 241408 3936 241460
rect 4988 241408 5040 241460
rect 422300 240796 422352 240848
rect 428464 240796 428516 240848
rect 435364 240728 435416 240780
rect 447784 240728 447836 240780
rect 361764 238688 361816 238740
rect 439596 238688 439648 238740
rect 414664 238008 414716 238060
rect 422300 238008 422352 238060
rect 386420 235220 386472 235272
rect 398472 235220 398524 235272
rect 570604 233180 570656 233232
rect 579988 233180 580040 233232
rect 427084 232500 427136 232552
rect 435364 232500 435416 232552
rect 384672 232024 384724 232076
rect 386420 232024 386472 232076
rect 361764 227672 361816 227724
rect 442264 227672 442316 227724
rect 455236 222096 455288 222148
rect 456800 222096 456852 222148
rect 394700 221416 394752 221468
rect 414664 221416 414716 221468
rect 428464 221416 428516 221468
rect 435456 221416 435508 221468
rect 559564 219376 559616 219428
rect 580172 219376 580224 219428
rect 391940 218016 391992 218068
rect 394700 218016 394752 218068
rect 361580 216316 361632 216368
rect 363604 216316 363656 216368
rect 387616 215296 387668 215348
rect 391940 215296 391992 215348
rect 3792 214752 3844 214804
rect 5080 214752 5132 214804
rect 411904 213188 411956 213240
rect 427084 213188 427136 213240
rect 379336 212984 379388 213036
rect 384672 212984 384724 213036
rect 448336 207612 448388 207664
rect 454040 207612 454092 207664
rect 456892 207612 456944 207664
rect 418068 207272 418120 207324
rect 422944 207272 422996 207324
rect 404084 205640 404136 205692
rect 411904 205640 411956 205692
rect 361764 205572 361816 205624
rect 439504 205572 439556 205624
rect 362316 204892 362368 204944
rect 379336 204892 379388 204944
rect 3976 204212 4028 204264
rect 5172 204212 5224 204264
rect 414664 201016 414716 201068
rect 418068 201016 418120 201068
rect 458732 200744 458784 200796
rect 481640 200744 481692 200796
rect 379336 199384 379388 199436
rect 387616 199384 387668 199436
rect 456800 197956 456852 198008
rect 485780 197956 485832 198008
rect 361672 194488 361724 194540
rect 443644 194488 443696 194540
rect 551284 193128 551336 193180
rect 580172 193128 580224 193180
rect 372620 189728 372672 189780
rect 379336 189728 379388 189780
rect 361212 186940 361264 186992
rect 372620 186940 372672 186992
rect 361672 183472 361724 183524
rect 436744 183472 436796 183524
rect 555424 179324 555476 179376
rect 580172 179324 580224 179376
rect 425060 178032 425112 178084
rect 428464 178032 428516 178084
rect 399576 176808 399628 176860
rect 404084 176808 404136 176860
rect 411260 171844 411312 171896
rect 425060 171844 425112 171896
rect 361764 171776 361816 171828
rect 440884 171776 440936 171828
rect 524420 171776 524472 171828
rect 404084 168376 404136 168428
rect 411260 168376 411312 168428
rect 537484 166948 537536 167000
rect 580172 166948 580224 167000
rect 411904 164840 411956 164892
rect 454040 164840 454092 164892
rect 402980 163480 403032 163532
rect 414664 163480 414716 163532
rect 448428 163480 448480 163532
rect 528560 163480 528612 163532
rect 445208 163072 445260 163124
rect 449992 163072 450044 163124
rect 418712 162188 418764 162240
rect 458088 162188 458140 162240
rect 414756 162120 414808 162172
rect 456800 162120 456852 162172
rect 489920 162120 489972 162172
rect 426164 161780 426216 161832
rect 496820 161780 496872 161832
rect 428648 161712 428700 161764
rect 500960 161712 501012 161764
rect 421380 161644 421432 161696
rect 494060 161644 494112 161696
rect 431868 161576 431920 161628
rect 505100 161576 505152 161628
rect 438768 161508 438820 161560
rect 513380 161508 513432 161560
rect 362408 161440 362460 161492
rect 441620 161440 441672 161492
rect 442908 161440 442960 161492
rect 517520 161440 517572 161492
rect 361764 161372 361816 161424
rect 444288 161372 444340 161424
rect 391940 160692 391992 160744
rect 402980 160692 403032 160744
rect 444288 160692 444340 160744
rect 521660 160692 521712 160744
rect 406844 160556 406896 160608
rect 414756 160556 414808 160608
rect 404176 160488 404228 160540
rect 411628 160488 411680 160540
rect 410524 160420 410576 160472
rect 418160 160420 418212 160472
rect 410616 160352 410668 160404
rect 425152 160352 425204 160404
rect 426164 160352 426216 160404
rect 407856 160284 407908 160336
rect 407764 160216 407816 160268
rect 411444 160216 411496 160268
rect 411628 160284 411680 160336
rect 421380 160284 421432 160336
rect 428004 160216 428056 160268
rect 409328 160148 409380 160200
rect 431316 160148 431368 160200
rect 435272 160148 435324 160200
rect 436008 160148 436060 160200
rect 451188 160148 451240 160200
rect 410708 160080 410760 160132
rect 438262 160080 438314 160132
rect 444886 160080 444938 160132
rect 445208 160080 445260 160132
rect 483664 160080 483716 160132
rect 363604 158720 363656 158772
rect 434812 159332 434864 159384
rect 451740 158380 451792 158432
rect 456708 158380 456760 158432
rect 452568 156884 452620 156936
rect 456616 156884 456668 156936
rect 382096 155184 382148 155236
rect 391940 155184 391992 155236
rect 547144 153144 547196 153196
rect 580172 153144 580224 153196
rect 452108 152940 452160 152992
rect 460480 152940 460532 152992
rect 452568 151444 452620 151496
rect 457812 151444 457864 151496
rect 393964 149064 394016 149116
rect 399576 149064 399628 149116
rect 452568 147364 452620 147416
rect 459468 147364 459520 147416
rect 452568 146140 452620 146192
rect 457536 146140 457588 146192
rect 452568 144644 452620 144696
rect 455052 144644 455104 144696
rect 452568 143284 452620 143336
rect 459376 143284 459428 143336
rect 483664 142876 483716 142928
rect 533988 142876 534040 142928
rect 451188 142808 451240 142860
rect 509608 142808 509660 142860
rect 533988 142128 534040 142180
rect 539784 142128 539836 142180
rect 452568 141924 452620 141976
rect 457628 141924 457680 141976
rect 388352 140768 388404 140820
rect 393964 140768 394016 140820
rect 452108 140632 452160 140684
rect 455144 140632 455196 140684
rect 530676 140088 530728 140140
rect 542544 140088 542596 140140
rect 530584 140020 530636 140072
rect 542452 140020 542504 140072
rect 379336 139408 379388 139460
rect 382096 139408 382148 139460
rect 361764 139340 361816 139392
rect 410708 139340 410760 139392
rect 452568 139340 452620 139392
rect 459284 139340 459336 139392
rect 554044 139340 554096 139392
rect 580172 139340 580224 139392
rect 538864 139204 538916 139256
rect 543188 139204 543240 139256
rect 452568 137844 452620 137896
rect 457720 137844 457772 137896
rect 538956 136552 539008 136604
rect 539508 136552 539560 136604
rect 452568 136484 452620 136536
rect 454776 136484 454828 136536
rect 363696 135872 363748 135924
rect 388352 135872 388404 135924
rect 452568 135124 452620 135176
rect 459192 135124 459244 135176
rect 452476 133764 452528 133816
rect 453764 133764 453816 133816
rect 452108 132404 452160 132456
rect 453672 132404 453724 132456
rect 361304 131112 361356 131164
rect 363696 131112 363748 131164
rect 452568 131044 452620 131096
rect 453948 131044 454000 131096
rect 373632 129004 373684 129056
rect 379336 129004 379388 129056
rect 361580 128188 361632 128240
rect 363604 128188 363656 128240
rect 452200 126896 452252 126948
rect 453212 126896 453264 126948
rect 576124 126896 576176 126948
rect 580172 126896 580224 126948
rect 451740 124720 451792 124772
rect 453856 124720 453908 124772
rect 451740 123088 451792 123140
rect 454868 123088 454920 123140
rect 451740 121592 451792 121644
rect 454960 121592 455012 121644
rect 369032 120232 369084 120284
rect 373632 120232 373684 120284
rect 362408 117920 362460 117972
rect 369032 117920 369084 117972
rect 361580 117240 361632 117292
rect 409328 117240 409380 117292
rect 573364 113092 573416 113144
rect 579804 113092 579856 113144
rect 359648 106904 359700 106956
rect 362408 106904 362460 106956
rect 361580 106224 361632 106276
rect 407856 106224 407908 106276
rect 569224 100648 569276 100700
rect 580172 100648 580224 100700
rect 361764 95140 361816 95192
rect 410616 95140 410668 95192
rect 394608 88952 394660 89004
rect 404084 88952 404136 89004
rect 574744 86912 574796 86964
rect 580172 86912 580224 86964
rect 3424 86232 3476 86284
rect 20904 86232 20956 86284
rect 388444 85552 388496 85604
rect 394608 85552 394660 85604
rect 361764 84124 361816 84176
rect 404176 84124 404228 84176
rect 361764 73108 361816 73160
rect 410524 73108 410576 73160
rect 548524 73108 548576 73160
rect 580172 73108 580224 73160
rect 4804 68960 4856 69012
rect 7380 68960 7432 69012
rect 7380 67464 7432 67516
rect 8668 67464 8720 67516
rect 4988 66172 5040 66224
rect 5816 66172 5868 66224
rect 359740 63520 359792 63572
rect 362316 63520 362368 63572
rect 449900 62772 449952 62824
rect 537484 62772 537536 62824
rect 5816 62092 5868 62144
rect 9588 62024 9640 62076
rect 361764 62024 361816 62076
rect 406844 62024 406896 62076
rect 5080 61276 5132 61328
rect 5540 61276 5592 61328
rect 385684 61208 385736 61260
rect 388444 61208 388496 61260
rect 544384 60664 544436 60716
rect 580172 60664 580224 60716
rect 3608 59984 3660 60036
rect 20904 59984 20956 60036
rect 8668 59304 8720 59356
rect 10324 59304 10376 59356
rect 372620 58624 372672 58676
rect 385684 58624 385736 58676
rect 9680 57944 9732 57996
rect 4896 57876 4948 57928
rect 6092 57876 6144 57928
rect 13728 57876 13780 57928
rect 5540 57196 5592 57248
rect 15200 57196 15252 57248
rect 368296 56312 368348 56364
rect 372620 56312 372672 56364
rect 6092 54476 6144 54528
rect 8208 54476 8260 54528
rect 15200 54476 15252 54528
rect 20904 54476 20956 54528
rect 5172 53796 5224 53848
rect 7380 53728 7432 53780
rect 13728 53728 13780 53780
rect 19248 53728 19300 53780
rect 361764 52368 361816 52420
rect 407764 52368 407816 52420
rect 10324 51756 10376 51808
rect 11244 51756 11296 51808
rect 540612 51076 540664 51128
rect 543740 51076 543792 51128
rect 7380 50804 7432 50856
rect 11336 50804 11388 50856
rect 8300 48288 8352 48340
rect 11244 48288 11296 48340
rect 11428 48220 11480 48272
rect 16488 48220 16540 48272
rect 11336 48152 11388 48204
rect 15200 48152 15252 48204
rect 3240 46996 3292 47048
rect 456524 46996 456576 47048
rect 3424 46860 3476 46912
rect 460296 46860 460348 46912
rect 563704 46860 563756 46912
rect 580172 46860 580224 46912
rect 3608 46792 3660 46844
rect 460388 46792 460440 46844
rect 4068 46724 4120 46776
rect 459008 46724 459060 46776
rect 3332 46656 3384 46708
rect 456340 46656 456392 46708
rect 3792 46588 3844 46640
rect 456432 46588 456484 46640
rect 3700 46520 3752 46572
rect 453580 46520 453632 46572
rect 3884 46452 3936 46504
rect 453488 46452 453540 46504
rect 3516 46384 3568 46436
rect 450912 46384 450964 46436
rect 19984 46316 20036 46368
rect 457444 46316 457496 46368
rect 21456 46248 21508 46300
rect 451096 46248 451148 46300
rect 21364 46180 21416 46232
rect 451004 46180 451056 46232
rect 15200 46112 15252 46164
rect 359740 46112 359792 46164
rect 358728 46044 358780 46096
rect 368296 46044 368348 46096
rect 3976 45500 4028 45552
rect 453396 45500 453448 45552
rect 3424 45432 3476 45484
rect 399484 45432 399536 45484
rect 11428 45364 11480 45416
rect 361304 45364 361356 45416
rect 16580 45296 16632 45348
rect 358728 45296 358780 45348
rect 69020 45228 69072 45280
rect 406660 45228 406712 45280
rect 64880 45160 64932 45212
rect 406384 45160 406436 45212
rect 60740 45092 60792 45144
rect 406568 45092 406620 45144
rect 57980 45024 58032 45076
rect 406476 45024 406528 45076
rect 51080 44956 51132 45008
rect 406752 44956 406804 45008
rect 46940 44888 46992 44940
rect 409144 44888 409196 44940
rect 53840 44820 53892 44872
rect 456248 44820 456300 44872
rect 71780 44752 71832 44804
rect 403992 44752 404044 44804
rect 86960 44684 87012 44736
rect 387524 44684 387576 44736
rect 107660 44616 107712 44668
rect 398380 44616 398432 44668
rect 103520 42712 103572 42764
rect 398288 42712 398340 42764
rect 100760 42644 100812 42696
rect 401140 42644 401192 42696
rect 74540 42576 74592 42628
rect 376484 42576 376536 42628
rect 96620 42508 96672 42560
rect 401048 42508 401100 42560
rect 93860 42440 93912 42492
rect 401232 42440 401284 42492
rect 89720 42372 89772 42424
rect 400956 42372 401008 42424
rect 85580 42304 85632 42356
rect 401324 42304 401376 42356
rect 82820 42236 82872 42288
rect 403808 42236 403860 42288
rect 78680 42168 78732 42220
rect 403716 42168 403768 42220
rect 75920 42100 75972 42152
rect 403624 42100 403676 42152
rect 11060 42032 11112 42084
rect 403900 42032 403952 42084
rect 110420 41964 110472 42016
rect 398196 41964 398248 42016
rect 111800 41896 111852 41948
rect 384580 41896 384632 41948
rect 114560 39992 114612 40044
rect 398104 39992 398156 40044
rect 91100 39924 91152 39976
rect 387340 39924 387392 39976
rect 59360 39856 59412 39908
rect 393044 39856 393096 39908
rect 55220 39788 55272 39840
rect 392952 39788 393004 39840
rect 118700 39720 118752 39772
rect 460204 39720 460256 39772
rect 44180 39652 44232 39704
rect 395620 39652 395672 39704
rect 40040 39584 40092 39636
rect 395436 39584 395488 39636
rect 35900 39516 35952 39568
rect 395804 39516 395856 39568
rect 20720 39448 20772 39500
rect 395528 39448 395580 39500
rect 2780 39380 2832 39432
rect 395712 39380 395764 39432
rect 33140 39312 33192 39364
rect 450820 39312 450872 39364
rect 104900 37204 104952 37256
rect 387432 37204 387484 37256
rect 102140 37136 102192 37188
rect 387156 37136 387208 37188
rect 98000 37068 98052 37120
rect 387064 37068 387116 37120
rect 93952 37000 94004 37052
rect 387248 37000 387300 37052
rect 84200 36932 84252 36984
rect 390100 36932 390152 36984
rect 80060 36864 80112 36916
rect 390284 36864 390336 36916
rect 77300 36796 77352 36848
rect 389916 36796 389968 36848
rect 73160 36728 73212 36780
rect 390008 36728 390060 36780
rect 69112 36660 69164 36712
rect 390192 36660 390244 36712
rect 66260 36592 66312 36644
rect 392860 36592 392912 36644
rect 62120 36524 62172 36576
rect 392768 36524 392820 36576
rect 109040 36456 109092 36508
rect 384488 36456 384540 36508
rect 115940 36388 115992 36440
rect 384396 36388 384448 36440
rect 60832 34416 60884 34468
rect 376392 34416 376444 34468
rect 56600 34348 56652 34400
rect 379152 34348 379204 34400
rect 49700 34280 49752 34332
rect 379244 34280 379296 34332
rect 44272 34212 44324 34264
rect 378876 34212 378928 34264
rect 41420 34144 41472 34196
rect 378968 34144 379020 34196
rect 37280 34076 37332 34128
rect 379060 34076 379112 34128
rect 34520 34008 34572 34060
rect 382004 34008 382056 34060
rect 30380 33940 30432 33992
rect 381820 33940 381872 33992
rect 22100 33872 22152 33924
rect 381912 33872 381964 33924
rect 17960 33804 18012 33856
rect 384304 33804 384356 33856
rect 9680 33736 9732 33788
rect 378784 33736 378836 33788
rect 118792 33668 118844 33720
rect 381728 33668 381780 33720
rect 122840 33600 122892 33652
rect 381544 33600 381596 33652
rect 3516 33056 3568 33108
rect 400864 33056 400916 33108
rect 565084 33056 565136 33108
rect 580172 33056 580224 33108
rect 113180 31696 113232 31748
rect 370964 31696 371016 31748
rect 106280 31628 106332 31680
rect 370688 31628 370740 31680
rect 99380 31560 99432 31612
rect 370780 31560 370832 31612
rect 95240 31492 95292 31544
rect 373356 31492 373408 31544
rect 88340 31424 88392 31476
rect 373540 31424 373592 31476
rect 85672 31356 85724 31408
rect 373264 31356 373316 31408
rect 77392 31288 77444 31340
rect 373448 31288 373500 31340
rect 70400 31220 70452 31272
rect 376208 31220 376260 31272
rect 67640 31152 67692 31204
rect 376116 31152 376168 31204
rect 63500 31084 63552 31136
rect 376300 31084 376352 31136
rect 19340 31016 19392 31068
rect 370872 31016 370924 31068
rect 117320 30948 117372 31000
rect 370504 30948 370556 31000
rect 120080 30880 120132 30932
rect 370596 30880 370648 30932
rect 45560 28432 45612 28484
rect 368020 28432 368072 28484
rect 42800 28364 42852 28416
rect 367836 28364 367888 28416
rect 38660 28296 38712 28348
rect 367928 28296 367980 28348
rect 31760 28228 31812 28280
rect 368112 28228 368164 28280
rect 3424 20612 3476 20664
rect 376024 20612 376076 20664
rect 566464 20612 566516 20664
rect 579988 20612 580040 20664
rect 3424 6808 3476 6860
rect 396724 6808 396776 6860
rect 562324 6808 562376 6860
rect 580172 6808 580224 6860
rect 52552 4088 52604 4140
rect 359464 4088 359516 4140
rect 35992 4020 36044 4072
rect 360936 4020 360988 4072
rect 124680 3952 124732 4004
rect 458824 3952 458876 4004
rect 48964 3884 49016 3936
rect 392676 3884 392728 3936
rect 14740 3816 14792 3868
rect 359556 3816 359608 3868
rect 27712 3748 27764 3800
rect 381636 3748 381688 3800
rect 82084 3680 82136 3732
rect 456064 3680 456116 3732
rect 13544 3612 13596 3664
rect 389824 3612 389876 3664
rect 17040 3544 17092 3596
rect 395344 3544 395396 3596
rect 24216 3476 24268 3528
rect 405004 3476 405056 3528
rect 53748 3408 53800 3460
rect 450636 3408 450688 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 85580 3340 85632 3392
rect 86500 3340 86552 3392
rect 92756 3340 92808 3392
rect 361120 3340 361172 3392
rect 103336 3272 103388 3324
rect 360844 3272 360896 3324
rect 110420 3204 110472 3256
rect 111616 3204 111668 3256
rect 110512 3136 110564 3188
rect 361028 3204 361080 3256
rect 30104 2116 30156 2168
rect 450544 2116 450596 2168
rect 2872 2048 2924 2100
rect 453304 2048 453356 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 6932 685166 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 23492 685234 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40512 700369 40540 703520
rect 40498 700360 40554 700369
rect 72988 700330 73016 703520
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 40498 700295 40554 700304
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 88352 685302 88380 702406
rect 105464 700398 105492 703520
rect 105452 700392 105504 700398
rect 105452 700334 105504 700340
rect 136652 689353 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 153212 692073 153240 702406
rect 170324 700466 170352 703520
rect 202800 700505 202828 703520
rect 218992 700534 219020 703520
rect 235184 700602 235212 703520
rect 235172 700596 235224 700602
rect 235172 700538 235224 700544
rect 218980 700528 219032 700534
rect 202786 700496 202842 700505
rect 170312 700460 170364 700466
rect 218980 700470 219032 700476
rect 202786 700431 202842 700440
rect 170312 700402 170364 700408
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 153198 692064 153254 692073
rect 153198 691999 153254 692008
rect 136638 689344 136694 689353
rect 136638 689279 136694 689288
rect 266372 686526 266400 697546
rect 282932 690713 282960 702406
rect 282918 690704 282974 690713
rect 282918 690639 282974 690648
rect 299492 687954 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 299480 687948 299532 687954
rect 299480 687890 299532 687896
rect 266360 686520 266412 686526
rect 266360 686462 266412 686468
rect 88340 685296 88392 685302
rect 88340 685238 88392 685244
rect 23480 685228 23532 685234
rect 23480 685170 23532 685176
rect 6920 685160 6972 685166
rect 6920 685102 6972 685108
rect 3976 684752 4028 684758
rect 3976 684694 4028 684700
rect 3148 684684 3200 684690
rect 3148 684626 3200 684632
rect 2872 682780 2924 682786
rect 2872 682722 2924 682728
rect 2884 673454 2912 682722
rect 2964 682712 3016 682718
rect 2964 682654 3016 682660
rect 2976 677770 3004 682654
rect 3160 677906 3188 684626
rect 3332 684616 3384 684622
rect 3332 684558 3384 684564
rect 3344 683114 3372 684558
rect 3884 684548 3936 684554
rect 3884 684490 3936 684496
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3792 683392 3844 683398
rect 3792 683334 3844 683340
rect 3700 683324 3752 683330
rect 3700 683266 3752 683272
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3516 683188 3568 683194
rect 3516 683130 3568 683136
rect 3344 683086 3464 683114
rect 3436 678450 3464 683086
rect 3528 678570 3556 683130
rect 3516 678564 3568 678570
rect 3516 678506 3568 678512
rect 3436 678422 3648 678450
rect 3516 678360 3568 678366
rect 3516 678302 3568 678308
rect 3160 677878 3464 677906
rect 2976 677742 3372 677770
rect 2884 673426 3280 673454
rect 3252 580009 3280 673426
rect 3238 580000 3294 580009
rect 3238 579935 3294 579944
rect 3344 566953 3372 677742
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 3436 462641 3464 677878
rect 3528 671265 3556 678302
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3514 669896 3570 669905
rect 3514 669831 3570 669840
rect 3422 462632 3478 462641
rect 3422 462567 3478 462576
rect 3528 449585 3556 669831
rect 3620 475697 3648 678422
rect 3712 632097 3740 683266
rect 3698 632088 3754 632097
rect 3698 632023 3754 632032
rect 3700 631372 3752 631378
rect 3700 631314 3752 631320
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3514 449576 3570 449585
rect 3514 449511 3570 449520
rect 3712 423609 3740 631314
rect 3804 501809 3832 683334
rect 3896 514865 3924 684490
rect 3988 527921 4016 684694
rect 331232 683806 331260 702986
rect 348804 700670 348832 703520
rect 364996 700738 365024 703520
rect 364984 700732 365036 700738
rect 364984 700674 365036 700680
rect 348792 700664 348844 700670
rect 348792 700606 348844 700612
rect 331220 683800 331272 683806
rect 331220 683742 331272 683748
rect 20904 683596 20956 683602
rect 20904 683538 20956 683544
rect 359464 683596 359516 683602
rect 359464 683538 359516 683544
rect 19984 683528 20036 683534
rect 19984 683470 20036 683476
rect 4068 683460 4120 683466
rect 4068 683402 4120 683408
rect 4080 553897 4108 683402
rect 18144 680400 18196 680406
rect 18144 680342 18196 680348
rect 18156 675306 18184 680342
rect 16580 675300 16632 675306
rect 16580 675242 16632 675248
rect 18144 675300 18196 675306
rect 18144 675242 18196 675248
rect 16592 670698 16620 675242
rect 16500 670670 16620 670698
rect 16500 667962 16528 670670
rect 13084 667956 13136 667962
rect 13084 667898 13136 667904
rect 16488 667956 16540 667962
rect 16488 667898 16540 667904
rect 13096 662454 13124 667898
rect 8944 662448 8996 662454
rect 8944 662390 8996 662396
rect 13084 662448 13136 662454
rect 13084 662390 13136 662396
rect 8956 652798 8984 662390
rect 8944 652792 8996 652798
rect 8944 652734 8996 652740
rect 4804 652724 4856 652730
rect 4804 652666 4856 652672
rect 4066 553888 4122 553897
rect 4066 553823 4122 553832
rect 3974 527912 4030 527921
rect 3974 527847 4030 527856
rect 3882 514856 3938 514865
rect 4816 514826 4844 652666
rect 19996 631378 20024 683470
rect 20916 680406 20944 683538
rect 20904 680400 20956 680406
rect 20904 680342 20956 680348
rect 19984 631372 20036 631378
rect 19984 631314 20036 631320
rect 359476 610026 359504 683538
rect 361764 679040 361816 679046
rect 361762 679008 361764 679017
rect 382924 679040 382976 679046
rect 361816 679008 361818 679017
rect 382924 678982 382976 678988
rect 361762 678943 361818 678952
rect 361762 667992 361818 668001
rect 361762 667927 361764 667936
rect 361816 667927 361818 667936
rect 378784 667956 378836 667962
rect 361764 667898 361816 667904
rect 378784 667898 378836 667904
rect 361762 656976 361818 656985
rect 361762 656911 361764 656920
rect 361816 656911 361818 656920
rect 361764 656882 361816 656888
rect 361762 645960 361818 645969
rect 361762 645895 361764 645904
rect 361816 645895 361818 645904
rect 376024 645924 376076 645930
rect 361764 645866 361816 645872
rect 376024 645866 376076 645872
rect 361578 634944 361634 634953
rect 361578 634879 361634 634888
rect 361592 634846 361620 634879
rect 361580 634840 361632 634846
rect 361580 634782 361632 634788
rect 361578 623928 361634 623937
rect 361578 623863 361634 623872
rect 361592 623830 361620 623863
rect 361580 623824 361632 623830
rect 361580 623766 361632 623772
rect 374644 623824 374696 623830
rect 374644 623766 374696 623772
rect 361578 612912 361634 612921
rect 361578 612847 361634 612856
rect 361592 612814 361620 612847
rect 361580 612808 361632 612814
rect 361580 612750 361632 612756
rect 359464 610020 359516 610026
rect 359464 609962 359516 609968
rect 365720 609952 365772 609958
rect 365720 609894 365772 609900
rect 365732 607170 365760 609894
rect 365720 607164 365772 607170
rect 365720 607106 365772 607112
rect 367836 607164 367888 607170
rect 367836 607106 367888 607112
rect 361578 601896 361634 601905
rect 361578 601831 361634 601840
rect 361592 601798 361620 601831
rect 361580 601792 361632 601798
rect 361580 601734 361632 601740
rect 367848 601730 367876 607106
rect 371884 601792 371936 601798
rect 371884 601734 371936 601740
rect 367836 601724 367888 601730
rect 367836 601666 367888 601672
rect 369124 601724 369176 601730
rect 369124 601666 369176 601672
rect 369136 595406 369164 601666
rect 369124 595400 369176 595406
rect 369124 595342 369176 595348
rect 370688 595400 370740 595406
rect 370688 595342 370740 595348
rect 370700 593366 370728 595342
rect 370688 593360 370740 593366
rect 370688 593302 370740 593308
rect 361762 590880 361818 590889
rect 361762 590815 361818 590824
rect 361776 590714 361804 590815
rect 361764 590708 361816 590714
rect 361764 590650 361816 590656
rect 370688 590708 370740 590714
rect 370688 590650 370740 590656
rect 361762 579864 361818 579873
rect 361762 579799 361818 579808
rect 361776 579698 361804 579799
rect 361764 579692 361816 579698
rect 361764 579634 361816 579640
rect 367744 579692 367796 579698
rect 367744 579634 367796 579640
rect 361578 568848 361634 568857
rect 361578 568783 361580 568792
rect 361632 568783 361634 568792
rect 363604 568812 363656 568818
rect 361580 568754 361632 568760
rect 363604 568754 363656 568760
rect 361578 557832 361634 557841
rect 361578 557767 361580 557776
rect 361632 557767 361634 557776
rect 361580 557738 361632 557744
rect 361762 546816 361818 546825
rect 361762 546751 361818 546760
rect 361776 546514 361804 546751
rect 361764 546508 361816 546514
rect 361764 546450 361816 546456
rect 361762 535800 361818 535809
rect 361762 535735 361818 535744
rect 361776 535498 361804 535735
rect 361764 535492 361816 535498
rect 361764 535434 361816 535440
rect 361762 524784 361818 524793
rect 361762 524719 361818 524728
rect 361776 524482 361804 524719
rect 361764 524476 361816 524482
rect 361764 524418 361816 524424
rect 3882 514791 3938 514800
rect 3976 514820 4028 514826
rect 3976 514762 4028 514768
rect 4804 514820 4856 514826
rect 4804 514762 4856 514768
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3698 423600 3754 423609
rect 3698 423535 3754 423544
rect 3988 410553 4016 514762
rect 361762 513768 361818 513777
rect 361762 513703 361818 513712
rect 361776 513398 361804 513703
rect 361764 513392 361816 513398
rect 361764 513334 361816 513340
rect 361762 502752 361818 502761
rect 361762 502687 361818 502696
rect 361776 502382 361804 502687
rect 361764 502376 361816 502382
rect 361764 502318 361816 502324
rect 361762 491736 361818 491745
rect 361762 491671 361818 491680
rect 361776 491366 361804 491671
rect 361764 491360 361816 491366
rect 361764 491302 361816 491308
rect 361762 480720 361818 480729
rect 361762 480655 361818 480664
rect 361776 480282 361804 480655
rect 361764 480276 361816 480282
rect 361764 480218 361816 480224
rect 361762 469704 361818 469713
rect 361762 469639 361818 469648
rect 361776 469266 361804 469639
rect 361764 469260 361816 469266
rect 361764 469202 361816 469208
rect 361762 458688 361818 458697
rect 361762 458623 361818 458632
rect 361776 458250 361804 458623
rect 361764 458244 361816 458250
rect 361764 458186 361816 458192
rect 361578 447672 361634 447681
rect 361578 447607 361634 447616
rect 361592 447234 361620 447607
rect 361580 447228 361632 447234
rect 361580 447170 361632 447176
rect 362222 436656 362278 436665
rect 362222 436591 362278 436600
rect 362236 416090 362264 436591
rect 362314 425640 362370 425649
rect 362314 425575 362370 425584
rect 362328 418810 362356 425575
rect 362316 418804 362368 418810
rect 362316 418746 362368 418752
rect 362224 416084 362276 416090
rect 362224 416026 362276 416032
rect 361578 414624 361634 414633
rect 361578 414559 361634 414568
rect 361592 414050 361620 414559
rect 361580 414044 361632 414050
rect 361580 413986 361632 413992
rect 3974 410544 4030 410553
rect 3974 410479 4030 410488
rect 361578 403608 361634 403617
rect 361578 403543 361634 403552
rect 361592 403034 361620 403543
rect 361580 403028 361632 403034
rect 361580 402970 361632 402976
rect 3790 397488 3846 397497
rect 3790 397423 3846 397432
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3514 345400 3570 345409
rect 3514 345335 3570 345344
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3252 47054 3280 136711
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3344 46714 3372 149767
rect 3436 86290 3464 306167
rect 3528 266422 3556 345335
rect 3620 305046 3648 358391
rect 3608 305040 3660 305046
rect 3608 304982 3660 304988
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3620 292602 3648 293111
rect 3608 292596 3660 292602
rect 3608 292538 3660 292544
rect 3606 267200 3662 267209
rect 3606 267135 3662 267144
rect 3516 266416 3568 266422
rect 3516 266358 3568 266364
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3424 86284 3476 86290
rect 3424 86226 3476 86232
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3436 46918 3464 71567
rect 3424 46912 3476 46918
rect 3424 46854 3476 46860
rect 3332 46708 3384 46714
rect 3332 46650 3384 46656
rect 3528 46442 3556 254079
rect 3620 60042 3648 267135
rect 3698 241088 3754 241097
rect 3698 241023 3754 241032
rect 3608 60036 3660 60042
rect 3608 59978 3660 59984
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3620 46850 3648 58511
rect 3608 46844 3660 46850
rect 3608 46786 3660 46792
rect 3712 46578 3740 241023
rect 3804 214810 3832 397423
rect 361578 392592 361634 392601
rect 361578 392527 361634 392536
rect 361592 392018 361620 392527
rect 361580 392012 361632 392018
rect 361580 391954 361632 391960
rect 361578 381576 361634 381585
rect 361578 381511 361634 381520
rect 361592 380934 361620 381511
rect 361580 380928 361632 380934
rect 361580 380870 361632 380876
rect 363616 378146 363644 568754
rect 363696 557796 363748 557802
rect 363696 557738 363748 557744
rect 363604 378140 363656 378146
rect 363604 378082 363656 378088
rect 363708 376718 363736 557738
rect 364984 480276 365036 480282
rect 364984 480218 365036 480224
rect 363788 447228 363840 447234
rect 363788 447170 363840 447176
rect 363696 376712 363748 376718
rect 363696 376654 363748 376660
rect 3974 371376 4030 371385
rect 3974 371311 4030 371320
rect 3882 319288 3938 319297
rect 3882 319223 3938 319232
rect 3896 241466 3924 319223
rect 3884 241460 3936 241466
rect 3884 241402 3936 241408
rect 3882 214976 3938 214985
rect 3882 214911 3938 214920
rect 3792 214804 3844 214810
rect 3792 214746 3844 214752
rect 3790 201920 3846 201929
rect 3790 201855 3846 201864
rect 3804 46646 3832 201855
rect 3792 46640 3844 46646
rect 3792 46582 3844 46588
rect 3700 46572 3752 46578
rect 3700 46514 3752 46520
rect 3896 46510 3924 214911
rect 3988 204270 4016 371311
rect 361578 370560 361634 370569
rect 361578 370495 361634 370504
rect 361592 369918 361620 370495
rect 361580 369912 361632 369918
rect 361580 369854 361632 369860
rect 363800 369850 363828 447170
rect 364996 372570 365024 480218
rect 367756 378078 367784 579634
rect 370504 386436 370556 386442
rect 370504 386378 370556 386384
rect 367744 378072 367796 378078
rect 367744 378014 367796 378020
rect 364984 372564 365036 372570
rect 364984 372506 365036 372512
rect 363788 369844 363840 369850
rect 363788 369786 363840 369792
rect 362222 359544 362278 359553
rect 362222 359479 362278 359488
rect 361762 348528 361818 348537
rect 361762 348463 361818 348472
rect 361776 347818 361804 348463
rect 361764 347812 361816 347818
rect 361764 347754 361816 347760
rect 362236 347750 362264 359479
rect 362224 347744 362276 347750
rect 362224 347686 362276 347692
rect 361764 340944 361816 340950
rect 361764 340886 361816 340892
rect 361776 337521 361804 340886
rect 361762 337512 361818 337521
rect 361762 337447 361818 337456
rect 362224 337408 362276 337414
rect 362224 337350 362276 337356
rect 362236 326505 362264 337350
rect 363604 334008 363656 334014
rect 363604 333950 363656 333956
rect 362222 326496 362278 326505
rect 362222 326431 362278 326440
rect 361764 315988 361816 315994
rect 361764 315930 361816 315936
rect 361776 315489 361804 315930
rect 361762 315480 361818 315489
rect 361762 315415 361818 315424
rect 359464 305652 359516 305658
rect 359464 305594 359516 305600
rect 4804 305040 4856 305046
rect 4804 304982 4856 304988
rect 3976 204264 4028 204270
rect 3976 204206 4028 204212
rect 3974 188864 4030 188873
rect 3974 188799 4030 188808
rect 3884 46504 3936 46510
rect 3884 46446 3936 46452
rect 3516 46436 3568 46442
rect 3516 46378 3568 46384
rect 3988 45558 4016 188799
rect 4066 162888 4122 162897
rect 4066 162823 4122 162832
rect 4080 46782 4108 162823
rect 4816 69018 4844 304982
rect 19984 292596 20036 292602
rect 19984 292538 20036 292544
rect 4896 266416 4948 266422
rect 4896 266358 4948 266364
rect 4804 69012 4856 69018
rect 4804 68954 4856 68960
rect 4908 57934 4936 266358
rect 4988 241460 5040 241466
rect 4988 241402 5040 241408
rect 5000 66230 5028 241402
rect 5080 214804 5132 214810
rect 5080 214746 5132 214752
rect 4988 66224 5040 66230
rect 4988 66166 5040 66172
rect 5092 61334 5120 214746
rect 5172 204264 5224 204270
rect 5172 204206 5224 204212
rect 5080 61328 5132 61334
rect 5080 61270 5132 61276
rect 4896 57928 4948 57934
rect 4896 57870 4948 57876
rect 5184 53854 5212 204206
rect 7380 69012 7432 69018
rect 7380 68954 7432 68960
rect 7392 67522 7420 68954
rect 7380 67516 7432 67522
rect 7380 67458 7432 67464
rect 8668 67516 8720 67522
rect 8668 67458 8720 67464
rect 5816 66224 5868 66230
rect 5816 66166 5868 66172
rect 5828 62150 5856 66166
rect 5816 62144 5868 62150
rect 5816 62086 5868 62092
rect 5540 61328 5592 61334
rect 5540 61270 5592 61276
rect 5552 57254 5580 61270
rect 8680 59362 8708 67458
rect 9588 62076 9640 62082
rect 9588 62018 9640 62024
rect 9600 60602 9628 62018
rect 9600 60574 9720 60602
rect 8668 59356 8720 59362
rect 8668 59298 8720 59304
rect 9692 58002 9720 60574
rect 10324 59356 10376 59362
rect 10324 59298 10376 59304
rect 9680 57996 9732 58002
rect 9680 57938 9732 57944
rect 6092 57928 6144 57934
rect 6092 57870 6144 57876
rect 5540 57248 5592 57254
rect 5540 57190 5592 57196
rect 6104 54534 6132 57870
rect 6092 54528 6144 54534
rect 6092 54470 6144 54476
rect 8208 54528 8260 54534
rect 8208 54470 8260 54476
rect 5172 53848 5224 53854
rect 5172 53790 5224 53796
rect 7380 53780 7432 53786
rect 7380 53722 7432 53728
rect 7392 50862 7420 53722
rect 8220 52442 8248 54470
rect 8220 52414 8340 52442
rect 7380 50856 7432 50862
rect 7380 50798 7432 50804
rect 8312 48346 8340 52414
rect 10336 51814 10364 59298
rect 13728 57928 13780 57934
rect 13728 57870 13780 57876
rect 13740 53786 13768 57870
rect 15200 57248 15252 57254
rect 15200 57190 15252 57196
rect 15212 54534 15240 57190
rect 15200 54528 15252 54534
rect 15200 54470 15252 54476
rect 13728 53780 13780 53786
rect 13728 53722 13780 53728
rect 19248 53780 19300 53786
rect 19248 53722 19300 53728
rect 10324 51808 10376 51814
rect 10324 51750 10376 51756
rect 11244 51808 11296 51814
rect 11244 51750 11296 51756
rect 11256 48346 11284 51750
rect 19260 50946 19288 53722
rect 19260 50918 19380 50946
rect 11336 50856 11388 50862
rect 11336 50798 11388 50804
rect 8300 48340 8352 48346
rect 8300 48282 8352 48288
rect 11244 48340 11296 48346
rect 11244 48282 11296 48288
rect 11348 48210 11376 50798
rect 19352 49609 19380 50918
rect 19338 49600 19394 49609
rect 19338 49535 19394 49544
rect 11428 48272 11480 48278
rect 11428 48214 11480 48220
rect 16488 48272 16540 48278
rect 16488 48214 16540 48220
rect 11336 48204 11388 48210
rect 11336 48146 11388 48152
rect 4068 46776 4120 46782
rect 4068 46718 4120 46724
rect 3976 45552 4028 45558
rect 3422 45520 3478 45529
rect 3976 45494 4028 45500
rect 3422 45455 3424 45464
rect 3476 45455 3478 45464
rect 3424 45426 3476 45432
rect 11440 45422 11468 48214
rect 15200 48204 15252 48210
rect 15200 48146 15252 48152
rect 15212 46170 15240 48146
rect 16500 46866 16528 48214
rect 16500 46838 16620 46866
rect 15200 46164 15252 46170
rect 15200 46106 15252 46112
rect 11428 45416 11480 45422
rect 11428 45358 11480 45364
rect 16592 45354 16620 46838
rect 19996 46374 20024 292538
rect 20904 86284 20956 86290
rect 20904 86226 20956 86232
rect 20916 84194 20944 86226
rect 20916 84166 21404 84194
rect 21376 64874 21404 84166
rect 21284 64846 21404 64874
rect 20904 60036 20956 60042
rect 20904 59978 20956 59984
rect 20916 59945 20944 59978
rect 20902 59936 20958 59945
rect 20902 59871 20958 59880
rect 21284 55298 21312 64846
rect 21454 59936 21510 59945
rect 21454 59871 21510 59880
rect 21284 55270 21404 55298
rect 20904 54528 20956 54534
rect 20904 54470 20956 54476
rect 20916 49473 20944 54470
rect 20902 49464 20958 49473
rect 20902 49399 20958 49408
rect 19984 46368 20036 46374
rect 19984 46310 20036 46316
rect 21376 46238 21404 55270
rect 21468 46306 21496 59871
rect 21456 46300 21508 46306
rect 21456 46242 21508 46248
rect 21364 46232 21416 46238
rect 21364 46174 21416 46180
rect 358728 46096 358780 46102
rect 358728 46038 358780 46044
rect 358740 45354 358768 46038
rect 16580 45348 16632 45354
rect 16580 45290 16632 45296
rect 358728 45348 358780 45354
rect 358728 45290 358780 45296
rect 69020 45280 69072 45286
rect 69020 45222 69072 45228
rect 64880 45212 64932 45218
rect 64880 45154 64932 45160
rect 60740 45144 60792 45150
rect 60740 45086 60792 45092
rect 57980 45076 58032 45082
rect 57980 45018 58032 45024
rect 51080 45008 51132 45014
rect 27618 44976 27674 44985
rect 51080 44950 51132 44956
rect 27618 44911 27674 44920
rect 46940 44940 46992 44946
rect 6918 44840 6974 44849
rect 6918 44775 6974 44784
rect 2780 39432 2832 39438
rect 2780 39374 2832 39380
rect 2792 16574 2820 39374
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 6932 16574 6960 44775
rect 11060 42084 11112 42090
rect 11060 42026 11112 42032
rect 9680 33788 9732 33794
rect 9680 33730 9732 33736
rect 2792 16546 3648 16574
rect 6932 16546 7696 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3431
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2884 480 2912 2042
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3620 354 3648 16546
rect 5262 3904 5318 3913
rect 5262 3839 5318 3848
rect 5276 480 5304 3839
rect 6458 3768 6514 3777
rect 6458 3703 6514 3712
rect 6472 480 6500 3703
rect 7668 480 7696 16546
rect 8758 3632 8814 3641
rect 8758 3567 8814 3576
rect 8772 480 8800 3567
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 33730
rect 11072 16574 11100 42026
rect 20720 39500 20772 39506
rect 20720 39442 20772 39448
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 11072 16546 11928 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 14740 3868 14792 3874
rect 14740 3810 14792 3816
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13556 480 13584 3606
rect 14752 480 14780 3810
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17052 480 17080 3538
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 33798
rect 19340 31068 19392 31074
rect 19340 31010 19392 31016
rect 19352 16574 19380 31010
rect 20732 16574 20760 39442
rect 26238 39264 26294 39273
rect 26238 39199 26294 39208
rect 22100 33924 22152 33930
rect 22100 33866 22152 33872
rect 22112 16574 22140 33866
rect 19352 16546 19472 16574
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 19444 480 19472 16546
rect 21836 480 21864 16546
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 480 24256 3470
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 39199
rect 27632 16574 27660 44911
rect 46940 44882 46992 44888
rect 44180 39704 44232 39710
rect 44180 39646 44232 39652
rect 40040 39636 40092 39642
rect 40040 39578 40092 39584
rect 35900 39568 35952 39574
rect 35900 39510 35952 39516
rect 33140 39364 33192 39370
rect 33140 39306 33192 39312
rect 30380 33992 30432 33998
rect 30380 33934 30432 33940
rect 30392 16574 30420 33934
rect 31760 28280 31812 28286
rect 31760 28222 31812 28228
rect 31772 16574 31800 28222
rect 33152 16574 33180 39306
rect 34520 34060 34572 34066
rect 34520 34002 34572 34008
rect 27632 16546 28488 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 27712 3800 27764 3806
rect 27712 3742 27764 3748
rect 27724 480 27752 3742
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 16546
rect 30104 2168 30156 2174
rect 30104 2110 30156 2116
rect 30116 480 30144 2110
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 34002
rect 35912 16574 35940 39510
rect 37280 34128 37332 34134
rect 37280 34070 37332 34076
rect 37292 16574 37320 34070
rect 38660 28348 38712 28354
rect 38660 28290 38712 28296
rect 38672 16574 38700 28290
rect 40052 16574 40080 39578
rect 41420 34196 41472 34202
rect 41420 34138 41472 34144
rect 41432 16574 41460 34138
rect 42800 28416 42852 28422
rect 42800 28358 42852 28364
rect 35912 16546 36768 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35992 4072 36044 4078
rect 35992 4014 36044 4020
rect 36004 480 36032 4014
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 28358
rect 44192 6914 44220 39646
rect 44272 34264 44324 34270
rect 44272 34206 44324 34212
rect 44284 16574 44312 34206
rect 45560 28484 45612 28490
rect 45560 28426 45612 28432
rect 45572 16574 45600 28426
rect 46952 16574 46980 44882
rect 49700 34332 49752 34338
rect 49700 34274 49752 34280
rect 49712 16574 49740 34274
rect 44284 16546 45048 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 44192 6886 44312 6914
rect 44284 480 44312 6886
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45020 354 45048 16546
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45020 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 3936 49016 3942
rect 48964 3878 49016 3884
rect 48976 480 49004 3878
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 44950
rect 53840 44872 53892 44878
rect 53840 44814 53892 44820
rect 53852 16574 53880 44814
rect 55220 39840 55272 39846
rect 55220 39782 55272 39788
rect 55232 16574 55260 39782
rect 56600 34400 56652 34406
rect 56600 34342 56652 34348
rect 56612 16574 56640 34342
rect 57992 16574 58020 45018
rect 59360 39908 59412 39914
rect 59360 39850 59412 39856
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52552 4140 52604 4146
rect 52552 4082 52604 4088
rect 52564 480 52592 4082
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 53760 480 53788 3402
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 39850
rect 60752 3398 60780 45086
rect 62120 36576 62172 36582
rect 62120 36518 62172 36524
rect 60832 34468 60884 34474
rect 60832 34410 60884 34416
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 34410
rect 62132 16574 62160 36518
rect 63500 31136 63552 31142
rect 63500 31078 63552 31084
rect 63512 16574 63540 31078
rect 64892 16574 64920 45154
rect 66260 36644 66312 36650
rect 66260 36586 66312 36592
rect 66272 16574 66300 36586
rect 67640 31204 67692 31210
rect 67640 31146 67692 31152
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 31146
rect 69032 6914 69060 45222
rect 71780 44804 71832 44810
rect 71780 44746 71832 44752
rect 69112 36712 69164 36718
rect 69112 36654 69164 36660
rect 69124 16574 69152 36654
rect 70400 31272 70452 31278
rect 70400 31214 70452 31220
rect 70412 16574 70440 31214
rect 71792 16574 71820 44746
rect 86960 44736 87012 44742
rect 86960 44678 87012 44684
rect 74540 42628 74592 42634
rect 74540 42570 74592 42576
rect 73160 36780 73212 36786
rect 73160 36722 73212 36728
rect 73172 16574 73200 36722
rect 74552 16574 74580 42570
rect 85580 42356 85632 42362
rect 85580 42298 85632 42304
rect 82820 42288 82872 42294
rect 82820 42230 82872 42236
rect 78680 42220 78732 42226
rect 78680 42162 78732 42168
rect 75920 42152 75972 42158
rect 75920 42094 75972 42100
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 42094
rect 77300 36848 77352 36854
rect 77300 36790 77352 36796
rect 77312 6914 77340 36790
rect 77392 31340 77444 31346
rect 77392 31282 77444 31288
rect 77404 16574 77432 31282
rect 78692 16574 78720 42162
rect 80060 36916 80112 36922
rect 80060 36858 80112 36864
rect 80072 16574 80100 36858
rect 82832 16574 82860 42230
rect 84200 36984 84252 36990
rect 84200 36926 84252 36932
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 82832 16546 83320 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 82084 3732 82136 3738
rect 82084 3674 82136 3680
rect 82096 480 82124 3674
rect 83292 480 83320 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 36926
rect 85592 3398 85620 42298
rect 85672 31408 85724 31414
rect 85672 31350 85724 31356
rect 85580 3392 85632 3398
rect 85580 3334 85632 3340
rect 85684 480 85712 31350
rect 86972 16574 87000 44678
rect 107660 44668 107712 44674
rect 107660 44610 107712 44616
rect 103520 42764 103572 42770
rect 103520 42706 103572 42712
rect 100760 42696 100812 42702
rect 100760 42638 100812 42644
rect 96620 42560 96672 42566
rect 96620 42502 96672 42508
rect 93860 42492 93912 42498
rect 93860 42434 93912 42440
rect 89720 42424 89772 42430
rect 89720 42366 89772 42372
rect 88340 31476 88392 31482
rect 88340 31418 88392 31424
rect 88352 16574 88380 31418
rect 89732 16574 89760 42366
rect 91100 39976 91152 39982
rect 91100 39918 91152 39924
rect 91112 16574 91140 39918
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 86500 3392 86552 3398
rect 86500 3334 86552 3340
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3334
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 93872 6914 93900 42434
rect 93952 37052 94004 37058
rect 93952 36994 94004 37000
rect 93964 16574 93992 36994
rect 95240 31544 95292 31550
rect 95240 31486 95292 31492
rect 95252 16574 95280 31486
rect 96632 16574 96660 42502
rect 98000 37120 98052 37126
rect 98000 37062 98052 37068
rect 98012 16574 98040 37062
rect 99380 31612 99432 31618
rect 99380 31554 99432 31560
rect 99392 16574 99420 31554
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 92756 3392 92808 3398
rect 92756 3334 92808 3340
rect 92768 480 92796 3334
rect 93964 480 93992 6886
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 42638
rect 102140 37188 102192 37194
rect 102140 37130 102192 37136
rect 102152 16574 102180 37130
rect 103532 16574 103560 42706
rect 104900 37256 104952 37262
rect 104900 37198 104952 37204
rect 104912 16574 104940 37198
rect 106280 31680 106332 31686
rect 106280 31622 106332 31628
rect 106292 16574 106320 31622
rect 107672 16574 107700 44610
rect 110420 42016 110472 42022
rect 110420 41958 110472 41964
rect 109040 36508 109092 36514
rect 109040 36450 109092 36456
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102244 480 102272 16546
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 103348 480 103376 3266
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 36450
rect 110432 3262 110460 41958
rect 111800 41948 111852 41954
rect 111800 41890 111852 41896
rect 111812 16574 111840 41890
rect 114560 40044 114612 40050
rect 114560 39986 114612 39992
rect 113180 31748 113232 31754
rect 113180 31690 113232 31696
rect 113192 16574 113220 31690
rect 114572 16574 114600 39986
rect 118700 39772 118752 39778
rect 118700 39714 118752 39720
rect 115940 36440 115992 36446
rect 115940 36382 115992 36388
rect 115952 16574 115980 36382
rect 117320 31000 117372 31006
rect 117320 30942 117372 30948
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110420 3256 110472 3262
rect 110420 3198 110472 3204
rect 111616 3256 111668 3262
rect 111616 3198 111668 3204
rect 110512 3188 110564 3194
rect 110512 3130 110564 3136
rect 110524 480 110552 3130
rect 111628 480 111656 3198
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 30942
rect 118712 6914 118740 39714
rect 121458 39400 121514 39409
rect 121458 39335 121514 39344
rect 118792 33720 118844 33726
rect 118792 33662 118844 33668
rect 118804 16574 118832 33662
rect 120080 30932 120132 30938
rect 120080 30874 120132 30880
rect 120092 16574 120120 30874
rect 121472 16574 121500 39335
rect 122840 33652 122892 33658
rect 122840 33594 122892 33600
rect 122852 16574 122880 33594
rect 118804 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 359476 4146 359504 305594
rect 361764 304972 361816 304978
rect 361764 304914 361816 304920
rect 361776 304473 361804 304914
rect 361762 304464 361818 304473
rect 361762 304399 361818 304408
rect 362224 304360 362276 304366
rect 362224 304302 362276 304308
rect 360844 304292 360896 304298
rect 360844 304234 360896 304240
rect 359556 269816 359608 269822
rect 359556 269758 359608 269764
rect 359464 4140 359516 4146
rect 359464 4082 359516 4088
rect 124680 4004 124732 4010
rect 124680 3946 124732 3952
rect 124692 480 124720 3946
rect 359568 3874 359596 269758
rect 359648 106956 359700 106962
rect 359648 106898 359700 106904
rect 359660 46345 359688 106898
rect 359740 63572 359792 63578
rect 359740 63514 359792 63520
rect 359646 46336 359702 46345
rect 359646 46271 359702 46280
rect 359752 46170 359780 63514
rect 359740 46164 359792 46170
rect 359740 46106 359792 46112
rect 359556 3868 359608 3874
rect 359556 3810 359608 3816
rect 360856 3330 360884 304234
rect 360936 302932 360988 302938
rect 360936 302874 360988 302880
rect 360948 4078 360976 302874
rect 361028 300144 361080 300150
rect 361028 300086 361080 300092
rect 360936 4072 360988 4078
rect 360936 4014 360988 4020
rect 360844 3324 360896 3330
rect 360844 3266 360896 3272
rect 361040 3262 361068 300086
rect 361120 297424 361172 297430
rect 361120 297366 361172 297372
rect 361132 3398 361160 297366
rect 361764 293956 361816 293962
rect 361764 293898 361816 293904
rect 361776 293457 361804 293898
rect 361762 293448 361818 293457
rect 361762 293383 361818 293392
rect 361764 282872 361816 282878
rect 361764 282814 361816 282820
rect 361776 282441 361804 282814
rect 361762 282432 361818 282441
rect 361762 282367 361818 282376
rect 361764 271856 361816 271862
rect 361764 271798 361816 271804
rect 361776 271425 361804 271798
rect 361762 271416 361818 271425
rect 361762 271351 361818 271360
rect 361764 260840 361816 260846
rect 361764 260782 361816 260788
rect 361776 260409 361804 260782
rect 361762 260400 361818 260409
rect 361762 260335 361818 260344
rect 361764 249756 361816 249762
rect 361764 249698 361816 249704
rect 361776 249393 361804 249698
rect 361762 249384 361818 249393
rect 361762 249319 361818 249328
rect 361764 238740 361816 238746
rect 361764 238682 361816 238688
rect 361776 238377 361804 238682
rect 361762 238368 361818 238377
rect 361762 238303 361818 238312
rect 361764 227724 361816 227730
rect 361764 227666 361816 227672
rect 361776 227361 361804 227666
rect 361762 227352 361818 227361
rect 361762 227287 361818 227296
rect 361580 216368 361632 216374
rect 361578 216336 361580 216345
rect 361632 216336 361634 216345
rect 361578 216271 361634 216280
rect 361764 205624 361816 205630
rect 361764 205566 361816 205572
rect 361776 205329 361804 205566
rect 361762 205320 361818 205329
rect 361762 205255 361818 205264
rect 361672 194540 361724 194546
rect 361672 194482 361724 194488
rect 361684 194313 361712 194482
rect 361670 194304 361726 194313
rect 361670 194239 361726 194248
rect 361212 186992 361264 186998
rect 361212 186934 361264 186940
rect 361224 46481 361252 186934
rect 361672 183524 361724 183530
rect 361672 183466 361724 183472
rect 361684 183297 361712 183466
rect 361670 183288 361726 183297
rect 361670 183223 361726 183232
rect 361762 172272 361818 172281
rect 361762 172207 361818 172216
rect 361776 171834 361804 172207
rect 361764 171828 361816 171834
rect 361764 171770 361816 171776
rect 361764 161424 361816 161430
rect 361764 161366 361816 161372
rect 361776 161265 361804 161366
rect 361762 161256 361818 161265
rect 361762 161191 361818 161200
rect 361764 139392 361816 139398
rect 361764 139334 361816 139340
rect 361776 139233 361804 139334
rect 361762 139224 361818 139233
rect 361762 139159 361818 139168
rect 361304 131164 361356 131170
rect 361304 131106 361356 131112
rect 361210 46472 361266 46481
rect 361210 46407 361266 46416
rect 361316 45422 361344 131106
rect 361580 128240 361632 128246
rect 361578 128208 361580 128217
rect 361632 128208 361634 128217
rect 361578 128143 361634 128152
rect 361580 117292 361632 117298
rect 361580 117234 361632 117240
rect 361592 117201 361620 117234
rect 361578 117192 361634 117201
rect 361578 117127 361634 117136
rect 361580 106276 361632 106282
rect 361580 106218 361632 106224
rect 361592 106185 361620 106218
rect 361578 106176 361634 106185
rect 361578 106111 361634 106120
rect 361764 95192 361816 95198
rect 361762 95160 361764 95169
rect 361816 95160 361818 95169
rect 361762 95095 361818 95104
rect 361764 84176 361816 84182
rect 361762 84144 361764 84153
rect 361816 84144 361818 84153
rect 361762 84079 361818 84088
rect 361764 73160 361816 73166
rect 361762 73128 361764 73137
rect 361816 73128 361818 73137
rect 361762 73063 361818 73072
rect 361762 62112 361818 62121
rect 361762 62047 361764 62056
rect 361816 62047 361818 62056
rect 361764 62018 361816 62024
rect 361764 52420 361816 52426
rect 361764 52362 361816 52368
rect 361776 51105 361804 52362
rect 361762 51096 361818 51105
rect 361762 51031 361818 51040
rect 361304 45416 361356 45422
rect 361304 45358 361356 45364
rect 362236 3913 362264 304302
rect 363616 216374 363644 333950
rect 368112 289536 368164 289542
rect 368112 289478 368164 289484
rect 367744 289400 367796 289406
rect 367744 289342 367796 289348
rect 363604 216368 363656 216374
rect 363604 216310 363656 216316
rect 362316 204944 362368 204950
rect 362316 204886 362368 204892
rect 362328 63578 362356 204886
rect 362408 161492 362460 161498
rect 362408 161434 362460 161440
rect 362420 150249 362448 161434
rect 363604 158772 363656 158778
rect 363604 158714 363656 158720
rect 362406 150240 362462 150249
rect 362406 150175 362462 150184
rect 363616 128246 363644 158714
rect 363696 135924 363748 135930
rect 363696 135866 363748 135872
rect 363708 131170 363736 135866
rect 363696 131164 363748 131170
rect 363696 131106 363748 131112
rect 363604 128240 363656 128246
rect 363604 128182 363656 128188
rect 362408 117972 362460 117978
rect 362408 117914 362460 117920
rect 362420 106962 362448 117914
rect 362408 106956 362460 106962
rect 362408 106898 362460 106904
rect 362316 63572 362368 63578
rect 362316 63514 362368 63520
rect 362222 3904 362278 3913
rect 362222 3839 362278 3848
rect 367756 3777 367784 289342
rect 368020 289264 368072 289270
rect 368020 289206 368072 289212
rect 367928 289196 367980 289202
rect 367928 289138 367980 289144
rect 367836 289128 367888 289134
rect 367836 289070 367888 289076
rect 367848 28422 367876 289070
rect 367836 28416 367888 28422
rect 367836 28358 367888 28364
rect 367940 28354 367968 289138
rect 368032 28490 368060 289206
rect 368020 28484 368072 28490
rect 368020 28426 368072 28432
rect 367928 28348 367980 28354
rect 367928 28290 367980 28296
rect 368124 28286 368152 289478
rect 368204 289468 368256 289474
rect 368204 289410 368256 289416
rect 368216 44985 368244 289410
rect 369032 120284 369084 120290
rect 369032 120226 369084 120232
rect 369044 117978 369072 120226
rect 369032 117972 369084 117978
rect 369032 117914 369084 117920
rect 368296 56364 368348 56370
rect 368296 56306 368348 56312
rect 368308 46102 368336 56306
rect 368296 46096 368348 46102
rect 368296 46038 368348 46044
rect 368202 44976 368258 44985
rect 368202 44911 368258 44920
rect 370516 31006 370544 386378
rect 370596 385076 370648 385082
rect 370596 385018 370648 385024
rect 370504 31000 370556 31006
rect 370504 30942 370556 30948
rect 370608 30938 370636 385018
rect 370700 379506 370728 590650
rect 370688 379500 370740 379506
rect 370688 379442 370740 379448
rect 371896 379438 371924 601734
rect 372620 593360 372672 593366
rect 372620 593302 372672 593308
rect 372632 590646 372660 593302
rect 372620 590640 372672 590646
rect 372620 590582 372672 590588
rect 374656 380866 374684 623766
rect 376036 382226 376064 645866
rect 376116 590640 376168 590646
rect 376116 590582 376168 590588
rect 376128 582418 376156 590582
rect 376116 582412 376168 582418
rect 376116 582354 376168 582360
rect 378796 383654 378824 667898
rect 378876 582412 378928 582418
rect 378876 582354 378928 582360
rect 378888 575006 378916 582354
rect 378876 575000 378928 575006
rect 378876 574942 378928 574948
rect 380808 575000 380860 575006
rect 380808 574942 380860 574948
rect 380820 571402 380848 574942
rect 380808 571396 380860 571402
rect 380808 571338 380860 571344
rect 381636 458244 381688 458250
rect 381636 458186 381688 458192
rect 381544 386504 381596 386510
rect 381544 386446 381596 386452
rect 378784 383648 378836 383654
rect 378784 383590 378836 383596
rect 376024 382220 376076 382226
rect 376024 382162 376076 382168
rect 374644 380860 374696 380866
rect 374644 380802 374696 380808
rect 371884 379432 371936 379438
rect 371884 379374 371936 379380
rect 378876 294840 378928 294846
rect 378876 294782 378928 294788
rect 378782 294536 378838 294545
rect 378782 294471 378838 294480
rect 373448 292528 373500 292534
rect 373448 292470 373500 292476
rect 370688 292120 370740 292126
rect 370688 292062 370740 292068
rect 370700 31686 370728 292062
rect 370780 292052 370832 292058
rect 370780 291994 370832 292000
rect 370688 31680 370740 31686
rect 370688 31622 370740 31628
rect 370792 31618 370820 291994
rect 373356 291916 373408 291922
rect 373356 291858 373408 291864
rect 373264 291848 373316 291854
rect 373264 291790 373316 291796
rect 370964 289332 371016 289338
rect 370964 289274 371016 289280
rect 370870 289096 370926 289105
rect 370870 289031 370926 289040
rect 370780 31612 370832 31618
rect 370780 31554 370832 31560
rect 370884 31074 370912 289031
rect 370976 31754 371004 289274
rect 372620 189780 372672 189786
rect 372620 189722 372672 189728
rect 372632 186998 372660 189722
rect 372620 186992 372672 186998
rect 372620 186934 372672 186940
rect 372620 58676 372672 58682
rect 372620 58618 372672 58624
rect 372632 56370 372660 58618
rect 372620 56364 372672 56370
rect 372620 56306 372672 56312
rect 370964 31748 371016 31754
rect 370964 31690 371016 31696
rect 373276 31414 373304 291790
rect 373368 31550 373396 291858
rect 373356 31544 373408 31550
rect 373356 31486 373408 31492
rect 373264 31408 373316 31414
rect 373264 31350 373316 31356
rect 373460 31346 373488 292470
rect 376484 292392 376536 292398
rect 376484 292334 376536 292340
rect 376116 292256 376168 292262
rect 376116 292198 376168 292204
rect 373540 291984 373592 291990
rect 373540 291926 373592 291932
rect 373552 31482 373580 291926
rect 376024 284980 376076 284986
rect 376024 284922 376076 284928
rect 373632 129056 373684 129062
rect 373632 128998 373684 129004
rect 373644 120290 373672 128998
rect 373632 120284 373684 120290
rect 373632 120226 373684 120232
rect 373540 31476 373592 31482
rect 373540 31418 373592 31424
rect 373448 31340 373500 31346
rect 373448 31282 373500 31288
rect 370872 31068 370924 31074
rect 370872 31010 370924 31016
rect 370596 30932 370648 30938
rect 370596 30874 370648 30880
rect 368112 28280 368164 28286
rect 368112 28222 368164 28228
rect 376036 20670 376064 284922
rect 376128 31210 376156 292198
rect 376300 292188 376352 292194
rect 376300 292130 376352 292136
rect 376208 291780 376260 291786
rect 376208 291722 376260 291728
rect 376220 31278 376248 291722
rect 376208 31272 376260 31278
rect 376208 31214 376260 31220
rect 376116 31204 376168 31210
rect 376116 31146 376168 31152
rect 376312 31142 376340 292130
rect 376390 291816 376446 291825
rect 376390 291751 376446 291760
rect 376404 34474 376432 291751
rect 376496 42634 376524 292334
rect 376484 42628 376536 42634
rect 376484 42570 376536 42576
rect 376392 34468 376444 34474
rect 376392 34410 376444 34416
rect 378796 33794 378824 294471
rect 378888 34270 378916 294782
rect 378968 294704 379020 294710
rect 378968 294646 379020 294652
rect 378876 34264 378928 34270
rect 378876 34206 378928 34212
rect 378980 34202 379008 294646
rect 379060 294636 379112 294642
rect 379060 294578 379112 294584
rect 378968 34196 379020 34202
rect 378968 34138 379020 34144
rect 379072 34134 379100 294578
rect 379152 292460 379204 292466
rect 379152 292402 379204 292408
rect 379164 34406 379192 292402
rect 379244 292324 379296 292330
rect 379244 292266 379296 292272
rect 379152 34400 379204 34406
rect 379152 34342 379204 34348
rect 379256 34338 379284 292266
rect 379336 213036 379388 213042
rect 379336 212978 379388 212984
rect 379348 204950 379376 212978
rect 379336 204944 379388 204950
rect 379336 204886 379388 204892
rect 379336 199436 379388 199442
rect 379336 199378 379388 199384
rect 379348 189786 379376 199378
rect 379336 189780 379388 189786
rect 379336 189722 379388 189728
rect 379336 139460 379388 139466
rect 379336 139402 379388 139408
rect 379348 129062 379376 139402
rect 379336 129056 379388 129062
rect 379336 128998 379388 129004
rect 379244 34332 379296 34338
rect 379244 34274 379296 34280
rect 379060 34128 379112 34134
rect 379060 34070 379112 34076
rect 378784 33788 378836 33794
rect 378784 33730 378836 33736
rect 381556 33658 381584 386446
rect 381648 371210 381676 458186
rect 382936 383586 382964 678982
rect 385684 571328 385736 571334
rect 385684 571270 385736 571276
rect 385696 560250 385724 571270
rect 385684 560244 385736 560250
rect 385684 560186 385736 560192
rect 387156 560244 387208 560250
rect 387156 560186 387208 560192
rect 387168 556238 387196 560186
rect 387156 556232 387208 556238
rect 387156 556174 387208 556180
rect 388444 556232 388496 556238
rect 388444 556174 388496 556180
rect 388456 522986 388484 556174
rect 388444 522980 388496 522986
rect 388444 522922 388496 522928
rect 389824 522980 389876 522986
rect 389824 522922 389876 522928
rect 389836 520266 389864 522922
rect 389824 520260 389876 520266
rect 389824 520202 389876 520208
rect 391204 520260 391256 520266
rect 391204 520202 391256 520208
rect 391216 500614 391244 520202
rect 391204 500608 391256 500614
rect 391204 500550 391256 500556
rect 393412 500608 393464 500614
rect 393412 500550 393464 500556
rect 393424 496262 393452 500550
rect 393412 496256 393464 496262
rect 393412 496198 393464 496204
rect 382924 383580 382976 383586
rect 382924 383522 382976 383528
rect 381636 371204 381688 371210
rect 381636 371146 381688 371152
rect 385684 338156 385736 338162
rect 385684 338098 385736 338104
rect 384304 295316 384356 295322
rect 384304 295258 384356 295264
rect 381912 295248 381964 295254
rect 381912 295190 381964 295196
rect 381634 294808 381690 294817
rect 381634 294743 381690 294752
rect 381728 294772 381780 294778
rect 381544 33652 381596 33658
rect 381544 33594 381596 33600
rect 376300 31136 376352 31142
rect 376300 31078 376352 31084
rect 376024 20664 376076 20670
rect 376024 20606 376076 20612
rect 381648 3806 381676 294743
rect 381728 294714 381780 294720
rect 381740 33726 381768 294714
rect 381818 294672 381874 294681
rect 381818 294607 381874 294616
rect 381832 33998 381860 294607
rect 381820 33992 381872 33998
rect 381820 33934 381872 33940
rect 381924 33930 381952 295190
rect 382004 294908 382056 294914
rect 382004 294850 382056 294856
rect 382016 34066 382044 294850
rect 382096 155236 382148 155242
rect 382096 155178 382148 155184
rect 382108 139466 382136 155178
rect 382096 139460 382148 139466
rect 382096 139402 382148 139408
rect 382004 34060 382056 34066
rect 382004 34002 382056 34008
rect 381912 33924 381964 33930
rect 381912 33866 381964 33872
rect 384316 33862 384344 295258
rect 384580 295180 384632 295186
rect 384580 295122 384632 295128
rect 384396 295112 384448 295118
rect 384396 295054 384448 295060
rect 384408 36446 384436 295054
rect 384488 294976 384540 294982
rect 384488 294918 384540 294924
rect 384500 36514 384528 294918
rect 384592 41954 384620 295122
rect 385696 293962 385724 338098
rect 397472 336054 397500 703520
rect 400864 656940 400916 656946
rect 400864 656882 400916 656888
rect 397552 496256 397604 496262
rect 397552 496198 397604 496204
rect 397564 489938 397592 496198
rect 397552 489932 397604 489938
rect 397552 489874 397604 489880
rect 400876 382158 400904 656882
rect 403624 634840 403676 634846
rect 403624 634782 403676 634788
rect 400956 489864 401008 489870
rect 400956 489806 401008 489812
rect 400968 476814 400996 489806
rect 400956 476808 401008 476814
rect 400956 476750 401008 476756
rect 402244 476808 402296 476814
rect 402244 476750 402296 476756
rect 402256 469878 402284 476750
rect 402244 469872 402296 469878
rect 402244 469814 402296 469820
rect 400864 382152 400916 382158
rect 400864 382094 400916 382100
rect 403636 380798 403664 634782
rect 406384 612808 406436 612814
rect 406384 612750 406436 612756
rect 406016 469872 406068 469878
rect 406016 469814 406068 469820
rect 406028 465118 406056 469814
rect 406016 465112 406068 465118
rect 406016 465054 406068 465060
rect 403624 380792 403676 380798
rect 403624 380734 403676 380740
rect 406396 380730 406424 612750
rect 407764 546508 407816 546514
rect 407764 546450 407816 546456
rect 406384 380724 406436 380730
rect 406384 380666 406436 380672
rect 407776 376650 407804 546450
rect 410524 535492 410576 535498
rect 410524 535434 410576 535440
rect 409144 465044 409196 465050
rect 409144 464986 409196 464992
rect 409156 458182 409184 464986
rect 409144 458176 409196 458182
rect 409144 458118 409196 458124
rect 409880 458176 409932 458182
rect 409880 458118 409932 458124
rect 409892 455462 409920 458118
rect 409880 455456 409932 455462
rect 409880 455398 409932 455404
rect 407764 376644 407816 376650
rect 407764 376586 407816 376592
rect 410536 375358 410564 535434
rect 411904 524476 411956 524482
rect 411904 524418 411956 524424
rect 410524 375352 410576 375358
rect 410524 375294 410576 375300
rect 411916 375290 411944 524418
rect 411904 375284 411956 375290
rect 411904 375226 411956 375232
rect 405740 350600 405792 350606
rect 405740 350542 405792 350548
rect 402244 347812 402296 347818
rect 402244 347754 402296 347760
rect 402256 342922 402284 347754
rect 402244 342916 402296 342922
rect 402244 342858 402296 342864
rect 399484 339516 399536 339522
rect 399484 339458 399536 339464
rect 397460 336048 397512 336054
rect 397460 335990 397512 335996
rect 399496 315994 399524 339458
rect 402256 334914 402284 342858
rect 402086 334886 402284 334914
rect 405752 334900 405780 350542
rect 412652 336122 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 700806 429884 703520
rect 429844 700800 429896 700806
rect 429844 700742 429896 700748
rect 449164 700800 449216 700806
rect 449164 700742 449216 700748
rect 445024 700732 445076 700738
rect 445024 700674 445076 700680
rect 444288 700460 444340 700466
rect 444288 700402 444340 700408
rect 418804 685296 418856 685302
rect 418804 685238 418856 685244
rect 417424 683528 417476 683534
rect 417424 683470 417476 683476
rect 414664 513392 414716 513398
rect 414664 513334 414716 513340
rect 414388 455388 414440 455394
rect 414388 455330 414440 455336
rect 414400 453354 414428 455330
rect 414388 453348 414440 453354
rect 414388 453290 414440 453296
rect 414676 373998 414704 513334
rect 416044 502376 416096 502382
rect 416044 502318 416096 502324
rect 414664 373992 414716 373998
rect 414664 373934 414716 373940
rect 416056 373930 416084 502318
rect 416688 453348 416740 453354
rect 416688 453290 416740 453296
rect 416700 447982 416728 453290
rect 416688 447976 416740 447982
rect 416688 447918 416740 447924
rect 416044 373924 416096 373930
rect 416044 373866 416096 373872
rect 416780 336796 416832 336802
rect 416780 336738 416832 336744
rect 412640 336116 412692 336122
rect 412640 336058 412692 336064
rect 413100 335436 413152 335442
rect 413100 335378 413152 335384
rect 409420 335368 409472 335374
rect 409420 335310 409472 335316
rect 409432 334900 409460 335310
rect 413112 334900 413140 335378
rect 416792 334900 416820 336738
rect 417436 334898 417464 683470
rect 417516 491360 417568 491366
rect 417516 491302 417568 491308
rect 417528 372502 417556 491302
rect 417516 372496 417568 372502
rect 417516 372438 417568 372444
rect 418160 341012 418212 341018
rect 418160 340954 418212 340960
rect 418172 337414 418200 340954
rect 418160 337408 418212 337414
rect 418160 337350 418212 337356
rect 418816 336258 418844 685238
rect 420368 684752 420420 684758
rect 420368 684694 420420 684700
rect 420184 684684 420236 684690
rect 420184 684626 420236 684632
rect 418896 683800 418948 683806
rect 418896 683742 418948 683748
rect 418804 336252 418856 336258
rect 418804 336194 418856 336200
rect 418908 336190 418936 683742
rect 418988 469260 419040 469266
rect 418988 469202 419040 469208
rect 419000 371142 419028 469202
rect 419080 447976 419132 447982
rect 419080 447918 419132 447924
rect 419092 420646 419120 447918
rect 419080 420640 419132 420646
rect 419080 420582 419132 420588
rect 418988 371136 419040 371142
rect 418988 371078 419040 371084
rect 418896 336184 418948 336190
rect 418896 336126 418948 336132
rect 417424 334892 417476 334898
rect 417424 334834 417476 334840
rect 420196 334830 420224 684626
rect 420274 684584 420330 684593
rect 420274 684519 420330 684528
rect 420184 334824 420236 334830
rect 420184 334766 420236 334772
rect 420288 334626 420316 684519
rect 420380 335102 420408 684694
rect 420552 684616 420604 684622
rect 420552 684558 420604 684564
rect 420460 336864 420512 336870
rect 420460 336806 420512 336812
rect 420368 335096 420420 335102
rect 420368 335038 420420 335044
rect 420472 334642 420500 336806
rect 420564 334762 420592 684558
rect 420736 683460 420788 683466
rect 420736 683402 420788 683408
rect 420644 683392 420696 683398
rect 420644 683334 420696 683340
rect 420552 334756 420604 334762
rect 420552 334698 420604 334704
rect 420656 334694 420684 683334
rect 420748 334966 420776 683402
rect 420828 682780 420880 682786
rect 420828 682722 420880 682728
rect 420840 335102 420868 682722
rect 436100 462460 436152 462466
rect 436100 462402 436152 462408
rect 433248 462392 433300 462398
rect 433248 462334 433300 462340
rect 423588 455456 423640 455462
rect 423588 455398 423640 455404
rect 423600 447574 423628 455398
rect 433260 447574 433288 462334
rect 422484 447568 422536 447574
rect 422484 447510 422536 447516
rect 423588 447568 423640 447574
rect 423588 447510 423640 447516
rect 432420 447568 432472 447574
rect 432420 447510 432472 447516
rect 433248 447568 433300 447574
rect 433248 447510 433300 447516
rect 422496 444924 422524 447510
rect 423600 447166 423628 447510
rect 423588 447160 423640 447166
rect 423588 447102 423640 447108
rect 432432 444924 432460 447510
rect 433260 447234 433288 447510
rect 433248 447228 433300 447234
rect 433248 447170 433300 447176
rect 436112 445738 436140 462402
rect 444196 447228 444248 447234
rect 444196 447170 444248 447176
rect 436100 445732 436152 445738
rect 436100 445674 436152 445680
rect 437388 445732 437440 445738
rect 437388 445674 437440 445680
rect 437400 444938 437428 445674
rect 437308 444924 437428 444938
rect 437308 444910 437414 444924
rect 427728 444576 427780 444582
rect 427478 444524 427728 444530
rect 427478 444518 427780 444524
rect 427478 444502 427768 444518
rect 437308 444514 437336 444910
rect 437296 444508 437348 444514
rect 437296 444450 437348 444456
rect 442632 444440 442684 444446
rect 442382 444388 442632 444394
rect 442382 444382 442684 444388
rect 444104 444440 444156 444446
rect 444104 444382 444156 444388
rect 442382 444366 442672 444382
rect 423956 420640 424008 420646
rect 423956 420582 424008 420588
rect 421484 417790 421512 420036
rect 421472 417784 421524 417790
rect 421472 417726 421524 417732
rect 422128 417518 422156 420036
rect 422312 420022 422786 420050
rect 422864 420022 423430 420050
rect 422116 417512 422168 417518
rect 422116 417454 422168 417460
rect 422312 391270 422340 420022
rect 422864 412634 422892 420022
rect 423968 416838 423996 420582
rect 442906 420200 442962 420209
rect 442906 420135 442962 420144
rect 424060 417654 424088 420036
rect 424048 417648 424100 417654
rect 424048 417590 424100 417596
rect 424704 417586 424732 420036
rect 425348 417722 425376 420036
rect 425336 417716 425388 417722
rect 425336 417658 425388 417664
rect 424692 417580 424744 417586
rect 424692 417522 424744 417528
rect 425992 417450 426020 420036
rect 440884 418804 440936 418810
rect 440884 418746 440936 418752
rect 425980 417444 426032 417450
rect 425980 417386 426032 417392
rect 423956 416832 424008 416838
rect 423956 416774 424008 416780
rect 428464 416832 428516 416838
rect 428464 416774 428516 416780
rect 422404 412606 422892 412634
rect 422404 392630 422432 412606
rect 428476 411330 428504 416774
rect 436744 416084 436796 416090
rect 436744 416026 436796 416032
rect 428464 411324 428516 411330
rect 428464 411266 428516 411272
rect 431224 411324 431276 411330
rect 431224 411266 431276 411272
rect 431236 400178 431264 411266
rect 431224 400172 431276 400178
rect 431224 400114 431276 400120
rect 432604 400172 432656 400178
rect 432604 400114 432656 400120
rect 422392 392624 422444 392630
rect 422392 392566 422444 392572
rect 422300 391264 422352 391270
rect 422300 391206 422352 391212
rect 432616 378010 432644 400114
rect 432604 378004 432656 378010
rect 432604 377946 432656 377952
rect 429200 369912 429252 369918
rect 429200 369854 429252 369860
rect 429212 365702 429240 369854
rect 436756 369782 436784 416026
rect 439504 414044 439556 414050
rect 439504 413986 439556 413992
rect 436836 378004 436888 378010
rect 436836 377946 436888 377952
rect 436744 369776 436796 369782
rect 436744 369718 436796 369724
rect 429200 365696 429252 365702
rect 429200 365638 429252 365644
rect 432604 362976 432656 362982
rect 432604 362918 432656 362924
rect 429844 336864 429896 336870
rect 429844 336806 429896 336812
rect 431224 336864 431276 336870
rect 431224 336806 431276 336812
rect 424138 335472 424194 335481
rect 424138 335407 424194 335416
rect 420828 335096 420880 335102
rect 420828 335038 420880 335044
rect 420736 334960 420788 334966
rect 420736 334902 420788 334908
rect 424152 334900 424180 335407
rect 420644 334688 420696 334694
rect 420472 334628 420592 334642
rect 420644 334630 420696 334636
rect 420276 334620 420328 334626
rect 420486 334614 420592 334628
rect 420276 334562 420328 334568
rect 420564 334506 420592 334614
rect 420734 334520 420790 334529
rect 420486 334478 420734 334506
rect 428094 334520 428150 334529
rect 427846 334478 428094 334506
rect 420734 334455 420790 334464
rect 428094 334455 428150 334464
rect 428108 334422 428136 334455
rect 428096 334416 428148 334422
rect 428096 334358 428148 334364
rect 429198 333024 429254 333033
rect 429198 332959 429254 332968
rect 429212 328438 429240 332959
rect 429200 328432 429252 328438
rect 429200 328374 429252 328380
rect 429856 327078 429884 336806
rect 429844 327072 429896 327078
rect 429844 327014 429896 327020
rect 399484 315988 399536 315994
rect 399484 315930 399536 315936
rect 409236 306332 409288 306338
rect 409236 306274 409288 306280
rect 409144 306264 409196 306270
rect 409144 306206 409196 306212
rect 406752 306196 406804 306202
rect 406752 306138 406804 306144
rect 400864 306128 400916 306134
rect 400864 306070 400916 306076
rect 398380 303476 398432 303482
rect 398380 303418 398432 303424
rect 398288 303136 398340 303142
rect 398288 303078 398340 303084
rect 398196 303068 398248 303074
rect 398196 303010 398248 303016
rect 396724 302796 396776 302802
rect 396724 302738 396776 302744
rect 395620 300620 395672 300626
rect 395620 300562 395672 300568
rect 395342 300520 395398 300529
rect 395342 300455 395398 300464
rect 395436 300484 395488 300490
rect 392768 300416 392820 300422
rect 392768 300358 392820 300364
rect 392676 300212 392728 300218
rect 392676 300154 392728 300160
rect 392582 300112 392638 300121
rect 392582 300047 392638 300056
rect 387248 297968 387300 297974
rect 387248 297910 387300 297916
rect 387156 297560 387208 297566
rect 387156 297502 387208 297508
rect 387064 297492 387116 297498
rect 387064 297434 387116 297440
rect 385684 293956 385736 293962
rect 385684 293898 385736 293904
rect 386420 235272 386472 235278
rect 386420 235214 386472 235220
rect 386432 232082 386460 235214
rect 384672 232076 384724 232082
rect 384672 232018 384724 232024
rect 386420 232076 386472 232082
rect 386420 232018 386472 232024
rect 384684 213042 384712 232018
rect 384672 213036 384724 213042
rect 384672 212978 384724 212984
rect 385684 61260 385736 61266
rect 385684 61202 385736 61208
rect 385696 58682 385724 61202
rect 385684 58676 385736 58682
rect 385684 58618 385736 58624
rect 384580 41948 384632 41954
rect 384580 41890 384632 41896
rect 387076 37126 387104 297434
rect 387168 37194 387196 297502
rect 387156 37188 387208 37194
rect 387156 37130 387208 37136
rect 387064 37120 387116 37126
rect 387064 37062 387116 37068
rect 387260 37058 387288 297910
rect 389916 297900 389968 297906
rect 389916 297842 389968 297848
rect 387524 297696 387576 297702
rect 387524 297638 387576 297644
rect 387340 297628 387392 297634
rect 387340 297570 387392 297576
rect 387352 39982 387380 297570
rect 387432 295044 387484 295050
rect 387432 294986 387484 294992
rect 387340 39976 387392 39982
rect 387340 39918 387392 39924
rect 387444 37262 387472 294986
rect 387536 44742 387564 297638
rect 389822 297392 389878 297401
rect 389822 297327 389878 297336
rect 387616 215348 387668 215354
rect 387616 215290 387668 215296
rect 387628 199442 387656 215290
rect 387616 199436 387668 199442
rect 387616 199378 387668 199384
rect 388352 140820 388404 140826
rect 388352 140762 388404 140768
rect 388364 135930 388392 140762
rect 388352 135924 388404 135930
rect 388352 135866 388404 135872
rect 388444 85604 388496 85610
rect 388444 85546 388496 85552
rect 388456 61266 388484 85546
rect 388444 61260 388496 61266
rect 388444 61202 388496 61208
rect 387524 44736 387576 44742
rect 387524 44678 387576 44684
rect 387432 37256 387484 37262
rect 387432 37198 387484 37204
rect 387248 37052 387300 37058
rect 387248 36994 387300 37000
rect 384488 36508 384540 36514
rect 384488 36450 384540 36456
rect 384396 36440 384448 36446
rect 384396 36382 384448 36388
rect 384304 33856 384356 33862
rect 384304 33798 384356 33804
rect 381728 33720 381780 33726
rect 381728 33662 381780 33668
rect 381636 3800 381688 3806
rect 367742 3768 367798 3777
rect 381636 3742 381688 3748
rect 367742 3703 367798 3712
rect 389836 3670 389864 297327
rect 389928 36854 389956 297842
rect 390192 297832 390244 297838
rect 390192 297774 390244 297780
rect 390100 297764 390152 297770
rect 390100 297706 390152 297712
rect 390008 297356 390060 297362
rect 390008 297298 390060 297304
rect 389916 36848 389968 36854
rect 389916 36790 389968 36796
rect 390020 36786 390048 297298
rect 390112 36990 390140 297706
rect 390100 36984 390152 36990
rect 390100 36926 390152 36932
rect 390008 36780 390060 36786
rect 390008 36722 390060 36728
rect 390204 36718 390232 297774
rect 390284 297288 390336 297294
rect 390284 297230 390336 297236
rect 390296 36922 390324 297230
rect 391940 218068 391992 218074
rect 391940 218010 391992 218016
rect 391952 215354 391980 218010
rect 391940 215348 391992 215354
rect 391940 215290 391992 215296
rect 391940 160744 391992 160750
rect 391940 160686 391992 160692
rect 391952 155242 391980 160686
rect 391940 155236 391992 155242
rect 391940 155178 391992 155184
rect 390284 36916 390336 36922
rect 390284 36858 390336 36864
rect 390192 36712 390244 36718
rect 390192 36654 390244 36660
rect 389824 3664 389876 3670
rect 392596 3641 392624 300047
rect 392688 3942 392716 300154
rect 392780 36582 392808 300358
rect 392952 300348 393004 300354
rect 392952 300290 393004 300296
rect 392860 298036 392912 298042
rect 392860 297978 392912 297984
rect 392872 36650 392900 297978
rect 392964 39846 392992 300290
rect 393044 300280 393096 300286
rect 393044 300222 393096 300228
rect 393056 39914 393084 300222
rect 394700 221468 394752 221474
rect 394700 221410 394752 221416
rect 394712 218074 394740 221410
rect 394700 218068 394752 218074
rect 394700 218010 394752 218016
rect 393964 149116 394016 149122
rect 393964 149058 394016 149064
rect 393976 140826 394004 149058
rect 393964 140820 394016 140826
rect 393964 140762 394016 140768
rect 394608 89004 394660 89010
rect 394608 88946 394660 88952
rect 394620 85610 394648 88946
rect 394608 85604 394660 85610
rect 394608 85546 394660 85552
rect 393044 39908 393096 39914
rect 393044 39850 393096 39856
rect 392952 39840 393004 39846
rect 392952 39782 393004 39788
rect 392860 36644 392912 36650
rect 392860 36586 392912 36592
rect 392768 36576 392820 36582
rect 392768 36518 392820 36524
rect 392676 3936 392728 3942
rect 392676 3878 392728 3884
rect 389824 3606 389876 3612
rect 392582 3632 392638 3641
rect 395356 3602 395384 300455
rect 395436 300426 395488 300432
rect 395448 39642 395476 300426
rect 395526 300248 395582 300257
rect 395526 300183 395582 300192
rect 395436 39636 395488 39642
rect 395436 39578 395488 39584
rect 395540 39506 395568 300183
rect 395632 39710 395660 300562
rect 395804 300552 395856 300558
rect 395804 300494 395856 300500
rect 395710 300384 395766 300393
rect 395710 300319 395766 300328
rect 395620 39704 395672 39710
rect 395620 39646 395672 39652
rect 395528 39500 395580 39506
rect 395528 39442 395580 39448
rect 395724 39438 395752 300319
rect 395816 39574 395844 300494
rect 395804 39568 395856 39574
rect 395804 39510 395856 39516
rect 395712 39432 395764 39438
rect 395712 39374 395764 39380
rect 396736 6866 396764 302738
rect 398104 300688 398156 300694
rect 398104 300630 398156 300636
rect 398116 40050 398144 300630
rect 398208 42022 398236 303010
rect 398300 42770 398328 303078
rect 398392 44674 398420 303418
rect 399484 291644 399536 291650
rect 399484 291586 399536 291592
rect 398472 243228 398524 243234
rect 398472 243170 398524 243176
rect 398484 235278 398512 243170
rect 398472 235272 398524 235278
rect 398472 235214 398524 235220
rect 399496 45490 399524 291586
rect 399576 176860 399628 176866
rect 399576 176802 399628 176808
rect 399588 149122 399616 176802
rect 399576 149116 399628 149122
rect 399576 149058 399628 149064
rect 399484 45484 399536 45490
rect 399484 45426 399536 45432
rect 398380 44668 398432 44674
rect 398380 44610 398432 44616
rect 398288 42764 398340 42770
rect 398288 42706 398340 42712
rect 398196 42016 398248 42022
rect 398196 41958 398248 41964
rect 398104 40044 398156 40050
rect 398104 39986 398156 39992
rect 400876 33114 400904 306070
rect 406476 306060 406528 306066
rect 406476 306002 406528 306008
rect 403992 305992 404044 305998
rect 403992 305934 404044 305940
rect 403624 305924 403676 305930
rect 403624 305866 403676 305872
rect 401048 303612 401100 303618
rect 401048 303554 401100 303560
rect 400956 303340 401008 303346
rect 400956 303282 401008 303288
rect 400968 42430 400996 303282
rect 401060 42566 401088 303554
rect 401232 303408 401284 303414
rect 401232 303350 401284 303356
rect 401140 303204 401192 303210
rect 401140 303146 401192 303152
rect 401152 42702 401180 303146
rect 401140 42696 401192 42702
rect 401140 42638 401192 42644
rect 401048 42560 401100 42566
rect 401048 42502 401100 42508
rect 401244 42498 401272 303350
rect 401324 303272 401376 303278
rect 401324 303214 401376 303220
rect 401232 42492 401284 42498
rect 401232 42434 401284 42440
rect 400956 42424 401008 42430
rect 400956 42366 401008 42372
rect 401336 42362 401364 303214
rect 401416 256012 401468 256018
rect 401416 255954 401468 255960
rect 401428 243234 401456 255954
rect 401416 243228 401468 243234
rect 401416 243170 401468 243176
rect 402980 163532 403032 163538
rect 402980 163474 403032 163480
rect 402992 160750 403020 163474
rect 402980 160744 403032 160750
rect 402980 160686 403032 160692
rect 401324 42356 401376 42362
rect 401324 42298 401376 42304
rect 403636 42158 403664 305866
rect 403808 303544 403860 303550
rect 403808 303486 403860 303492
rect 403716 302864 403768 302870
rect 403716 302806 403768 302812
rect 403728 42226 403756 302806
rect 403820 42294 403848 303486
rect 403898 302832 403954 302841
rect 403898 302767 403954 302776
rect 403808 42288 403860 42294
rect 403808 42230 403860 42236
rect 403716 42220 403768 42226
rect 403716 42162 403768 42168
rect 403624 42152 403676 42158
rect 403624 42094 403676 42100
rect 403912 42090 403940 302767
rect 404004 44810 404032 305934
rect 406384 305720 406436 305726
rect 406384 305662 406436 305668
rect 405004 289604 405056 289610
rect 405004 289546 405056 289552
rect 404084 205692 404136 205698
rect 404084 205634 404136 205640
rect 404096 176866 404124 205634
rect 404084 176860 404136 176866
rect 404084 176802 404136 176808
rect 404084 168428 404136 168434
rect 404084 168370 404136 168376
rect 404096 89010 404124 168370
rect 404176 160540 404228 160546
rect 404176 160482 404228 160488
rect 404084 89004 404136 89010
rect 404084 88946 404136 88952
rect 404188 84182 404216 160482
rect 404176 84176 404228 84182
rect 404176 84118 404228 84124
rect 403992 44804 404044 44810
rect 403992 44746 404044 44752
rect 403900 42084 403952 42090
rect 403900 42026 403952 42032
rect 400864 33108 400916 33114
rect 400864 33050 400916 33056
rect 396724 6860 396776 6866
rect 396724 6802 396776 6808
rect 392582 3567 392638 3576
rect 395344 3596 395396 3602
rect 395344 3538 395396 3544
rect 405016 3534 405044 289546
rect 406396 45218 406424 305662
rect 406384 45212 406436 45218
rect 406384 45154 406436 45160
rect 406488 45082 406516 306002
rect 406568 305856 406620 305862
rect 406568 305798 406620 305804
rect 406580 45150 406608 305798
rect 406660 305788 406712 305794
rect 406660 305730 406712 305736
rect 406672 45286 406700 305730
rect 406660 45280 406712 45286
rect 406660 45222 406712 45228
rect 406568 45144 406620 45150
rect 406568 45086 406620 45092
rect 406476 45076 406528 45082
rect 406476 45018 406528 45024
rect 406764 45014 406792 306138
rect 406844 160608 406896 160614
rect 406844 160550 406896 160556
rect 406856 62082 406884 160550
rect 407856 160336 407908 160342
rect 407856 160278 407908 160284
rect 407764 160268 407816 160274
rect 407764 160210 407816 160216
rect 406844 62076 406896 62082
rect 406844 62018 406896 62024
rect 407776 52426 407804 160210
rect 407868 106282 407896 160278
rect 407856 106276 407908 106282
rect 407856 106218 407908 106224
rect 407764 52420 407816 52426
rect 407764 52362 407816 52368
rect 406752 45008 406804 45014
rect 406752 44950 406804 44956
rect 409156 44946 409184 306206
rect 409144 44940 409196 44946
rect 409144 44882 409196 44888
rect 409248 44849 409276 306274
rect 431236 271862 431264 336806
rect 431316 335368 431368 335374
rect 431316 335310 431368 335316
rect 431328 324970 431356 335310
rect 432616 332897 432644 362918
rect 435456 360256 435508 360262
rect 435456 360198 435508 360204
rect 432696 344344 432748 344350
rect 432696 344286 432748 344292
rect 432602 332888 432658 332897
rect 432602 332823 432658 332832
rect 432604 330064 432656 330070
rect 432604 330006 432656 330012
rect 431868 329112 431920 329118
rect 431868 329054 431920 329060
rect 431316 324964 431368 324970
rect 431316 324906 431368 324912
rect 431224 271856 431276 271862
rect 431224 271798 431276 271804
rect 420920 264308 420972 264314
rect 420920 264250 420972 264256
rect 420932 261526 420960 264250
rect 422944 264240 422996 264246
rect 422944 264182 422996 264188
rect 411904 261520 411956 261526
rect 411904 261462 411956 261468
rect 420920 261520 420972 261526
rect 420920 261462 420972 261468
rect 411916 256018 411944 261462
rect 411904 256012 411956 256018
rect 411904 255954 411956 255960
rect 422300 240848 422352 240854
rect 422300 240790 422352 240796
rect 422312 238066 422340 240790
rect 414664 238060 414716 238066
rect 414664 238002 414716 238008
rect 422300 238060 422352 238066
rect 422300 238002 422352 238008
rect 414676 221474 414704 238002
rect 414664 221468 414716 221474
rect 414664 221410 414716 221416
rect 411904 213240 411956 213246
rect 411904 213182 411956 213188
rect 411916 205698 411944 213182
rect 422956 207330 422984 264182
rect 431224 262880 431276 262886
rect 431224 262822 431276 262828
rect 431236 253978 431264 262822
rect 428464 253972 428516 253978
rect 428464 253914 428516 253920
rect 431224 253972 431276 253978
rect 431224 253914 431276 253920
rect 428476 240854 428504 253914
rect 428464 240848 428516 240854
rect 428464 240790 428516 240796
rect 427084 232552 427136 232558
rect 427084 232494 427136 232500
rect 427096 213246 427124 232494
rect 428464 221468 428516 221474
rect 428464 221410 428516 221416
rect 427084 213240 427136 213246
rect 427084 213182 427136 213188
rect 418068 207324 418120 207330
rect 418068 207266 418120 207272
rect 422944 207324 422996 207330
rect 422944 207266 422996 207272
rect 411904 205692 411956 205698
rect 411904 205634 411956 205640
rect 418080 201074 418108 207266
rect 414664 201068 414716 201074
rect 414664 201010 414716 201016
rect 418068 201068 418120 201074
rect 418068 201010 418120 201016
rect 411260 171896 411312 171902
rect 411260 171838 411312 171844
rect 411272 168434 411300 171838
rect 411260 168428 411312 168434
rect 411260 168370 411312 168376
rect 411904 164892 411956 164898
rect 411904 164834 411956 164840
rect 411628 160540 411680 160546
rect 411628 160482 411680 160488
rect 410524 160472 410576 160478
rect 410524 160414 410576 160420
rect 409328 160200 409380 160206
rect 409328 160142 409380 160148
rect 409340 117298 409368 160142
rect 409328 117292 409380 117298
rect 409328 117234 409380 117240
rect 410536 73166 410564 160414
rect 410616 160404 410668 160410
rect 410616 160346 410668 160352
rect 410628 95198 410656 160346
rect 411640 160342 411668 160482
rect 411628 160336 411680 160342
rect 411628 160278 411680 160284
rect 411444 160268 411496 160274
rect 411444 160210 411496 160216
rect 410708 160132 410760 160138
rect 410708 160074 410760 160080
rect 410720 139398 410748 160074
rect 411456 159882 411484 160210
rect 411916 159882 411944 164834
rect 414676 163538 414704 201010
rect 428476 178090 428504 221410
rect 425060 178084 425112 178090
rect 425060 178026 425112 178032
rect 428464 178084 428516 178090
rect 428464 178026 428516 178032
rect 425072 171902 425100 178026
rect 425060 171896 425112 171902
rect 425060 171838 425112 171844
rect 414664 163532 414716 163538
rect 414664 163474 414716 163480
rect 421378 162752 421434 162761
rect 421378 162687 421434 162696
rect 426162 162752 426218 162761
rect 426162 162687 426218 162696
rect 428646 162752 428702 162761
rect 428646 162687 428702 162696
rect 418712 162240 418764 162246
rect 418712 162182 418764 162188
rect 414756 162172 414808 162178
rect 414756 162114 414808 162120
rect 414768 160614 414796 162114
rect 414756 160608 414808 160614
rect 414756 160550 414808 160556
rect 411456 159854 411944 159882
rect 414768 159882 414796 160550
rect 418160 160472 418212 160478
rect 418160 160414 418212 160420
rect 418172 159882 418200 160414
rect 418724 159882 418752 162182
rect 421392 161702 421420 162687
rect 426176 161838 426204 162687
rect 426164 161832 426216 161838
rect 426164 161774 426216 161780
rect 421380 161696 421432 161702
rect 421380 161638 421432 161644
rect 421392 160342 421420 161638
rect 426176 160410 426204 161774
rect 428660 161770 428688 162687
rect 428648 161764 428700 161770
rect 428648 161706 428700 161712
rect 425152 160404 425204 160410
rect 425152 160346 425204 160352
rect 426164 160404 426216 160410
rect 426164 160346 426216 160352
rect 421380 160336 421432 160342
rect 421380 160278 421432 160284
rect 414768 159854 415104 159882
rect 418172 159854 418752 159882
rect 421392 159882 421420 160278
rect 421392 159854 421728 159882
rect 425164 159746 425192 160346
rect 428004 160268 428056 160274
rect 428004 160210 428056 160216
rect 428016 159882 428044 160210
rect 428660 159882 428688 161706
rect 431880 161634 431908 329054
rect 432616 318209 432644 330006
rect 432708 325553 432736 344286
rect 435364 335368 435416 335374
rect 435364 335310 435416 335316
rect 432972 332648 433024 332654
rect 432972 332590 433024 332596
rect 432788 331288 432840 331294
rect 432788 331230 432840 331236
rect 432694 325544 432750 325553
rect 432694 325479 432750 325488
rect 432696 323604 432748 323610
rect 432696 323546 432748 323552
rect 432602 318200 432658 318209
rect 432602 318135 432658 318144
rect 432708 314537 432736 323546
rect 432800 321881 432828 331230
rect 432984 329225 433012 332590
rect 432970 329216 433026 329225
rect 432970 329151 433026 329160
rect 432786 321872 432842 321881
rect 432786 321807 432842 321816
rect 432694 314528 432750 314537
rect 432694 314463 432750 314472
rect 432604 311160 432656 311166
rect 432604 311102 432656 311108
rect 432616 310865 432644 311102
rect 432602 310856 432658 310865
rect 432602 310791 432658 310800
rect 432420 307760 432472 307766
rect 432420 307702 432472 307708
rect 432432 307193 432460 307702
rect 432418 307184 432474 307193
rect 432418 307119 432474 307128
rect 435376 249762 435404 335310
rect 435468 330070 435496 360198
rect 436848 343942 436876 377946
rect 439516 368490 439544 413986
rect 439504 368484 439556 368490
rect 439504 368426 439556 368432
rect 440896 368422 440924 418746
rect 442920 412634 442948 420135
rect 442828 412606 442948 412634
rect 442264 403028 442316 403034
rect 442264 402970 442316 402976
rect 440976 392012 441028 392018
rect 440976 391954 441028 391960
rect 440884 368416 440936 368422
rect 440884 368358 440936 368364
rect 440988 367062 441016 391954
rect 440976 367056 441028 367062
rect 440976 366998 441028 367004
rect 442276 366994 442304 402970
rect 442356 380928 442408 380934
rect 442356 380870 442408 380876
rect 442264 366988 442316 366994
rect 442264 366930 442316 366936
rect 442368 365634 442396 380870
rect 442356 365628 442408 365634
rect 442356 365570 442408 365576
rect 437020 363044 437072 363050
rect 437020 362986 437072 362992
rect 436928 358828 436980 358834
rect 436928 358770 436980 358776
rect 436836 343936 436888 343942
rect 436836 343878 436888 343884
rect 436836 338224 436888 338230
rect 436836 338166 436888 338172
rect 435548 335436 435600 335442
rect 435548 335378 435600 335384
rect 435456 330064 435508 330070
rect 435456 330006 435508 330012
rect 435560 325582 435588 335378
rect 436744 332716 436796 332722
rect 436744 332658 436796 332664
rect 436008 328500 436060 328506
rect 436008 328442 436060 328448
rect 435548 325576 435600 325582
rect 435548 325518 435600 325524
rect 435456 267028 435508 267034
rect 435456 266970 435508 266976
rect 435364 249756 435416 249762
rect 435364 249698 435416 249704
rect 435364 240780 435416 240786
rect 435364 240722 435416 240728
rect 435376 232558 435404 240722
rect 435364 232552 435416 232558
rect 435364 232494 435416 232500
rect 435468 221474 435496 266970
rect 435456 221468 435508 221474
rect 435456 221410 435508 221416
rect 431868 161628 431920 161634
rect 431868 161570 431920 161576
rect 431316 160200 431368 160206
rect 431316 160142 431368 160148
rect 428016 159854 428688 159882
rect 431328 159882 431356 160142
rect 431880 159882 431908 161570
rect 436020 160206 436048 328442
rect 436756 183530 436784 332658
rect 436848 282878 436876 338166
rect 436940 307766 436968 358770
rect 437032 332654 437060 362986
rect 442264 361684 442316 361690
rect 442264 361626 442316 361632
rect 439688 361616 439740 361622
rect 439688 361558 439740 361564
rect 439136 343936 439188 343942
rect 439136 343878 439188 343884
rect 439148 338094 439176 343878
rect 439136 338088 439188 338094
rect 439136 338030 439188 338036
rect 438124 336252 438176 336258
rect 438124 336194 438176 336200
rect 437020 332648 437072 332654
rect 437020 332590 437072 332596
rect 438136 320754 438164 336194
rect 439504 332852 439556 332858
rect 439504 332794 439556 332800
rect 438768 330540 438820 330546
rect 438768 330482 438820 330488
rect 438124 320748 438176 320754
rect 438124 320690 438176 320696
rect 436928 307760 436980 307766
rect 436928 307702 436980 307708
rect 436836 282872 436888 282878
rect 436836 282814 436888 282820
rect 436744 183524 436796 183530
rect 436744 183466 436796 183472
rect 438780 161566 438808 330482
rect 439516 205630 439544 332794
rect 439700 331294 439728 361558
rect 441068 358896 441120 358902
rect 441068 358838 441120 358844
rect 439872 336796 439924 336802
rect 439872 336738 439924 336744
rect 440976 336796 441028 336802
rect 440976 336738 441028 336744
rect 439780 335436 439832 335442
rect 439780 335378 439832 335384
rect 439688 331288 439740 331294
rect 439688 331230 439740 331236
rect 439792 316034 439820 335378
rect 439884 327010 439912 336738
rect 440884 331288 440936 331294
rect 440884 331230 440936 331236
rect 439872 327004 439924 327010
rect 439872 326946 439924 326952
rect 439608 316006 439820 316034
rect 439608 238746 439636 316006
rect 439688 289672 439740 289678
rect 439688 289614 439740 289620
rect 439700 264314 439728 289614
rect 439688 264308 439740 264314
rect 439688 264250 439740 264256
rect 439596 238740 439648 238746
rect 439596 238682 439648 238688
rect 439504 205624 439556 205630
rect 439504 205566 439556 205572
rect 440896 171834 440924 331230
rect 440988 260846 441016 336738
rect 441080 311166 441108 358838
rect 442276 344350 442304 361626
rect 442356 360324 442408 360330
rect 442356 360266 442408 360272
rect 442264 344344 442316 344350
rect 442264 344286 442316 344292
rect 441252 338088 441304 338094
rect 441252 338030 441304 338036
rect 441160 336048 441212 336054
rect 441160 335990 441212 335996
rect 441172 320822 441200 335990
rect 441264 322318 441292 338030
rect 441344 336184 441396 336190
rect 441344 336126 441396 336132
rect 441252 322312 441304 322318
rect 441252 322254 441304 322260
rect 441160 320816 441212 320822
rect 441160 320758 441212 320764
rect 441356 320550 441384 336126
rect 442264 334076 442316 334082
rect 442264 334018 442316 334024
rect 441344 320544 441396 320550
rect 441344 320486 441396 320492
rect 441068 311160 441120 311166
rect 441068 311102 441120 311108
rect 440976 260840 441028 260846
rect 440976 260782 441028 260788
rect 442276 227730 442304 334018
rect 442368 323610 442396 360266
rect 442356 323604 442408 323610
rect 442356 323546 442408 323552
rect 442828 318782 442856 412606
rect 443736 339584 443788 339590
rect 443736 339526 443788 339532
rect 443644 332648 443696 332654
rect 443644 332590 443696 332596
rect 442908 330608 442960 330614
rect 442908 330550 442960 330556
rect 442816 318776 442868 318782
rect 442816 318718 442868 318724
rect 442264 227724 442316 227730
rect 442264 227666 442316 227672
rect 440884 171828 440936 171834
rect 440884 171770 440936 171776
rect 438768 161560 438820 161566
rect 438768 161502 438820 161508
rect 438780 161474 438808 161502
rect 442920 161498 442948 330550
rect 443656 194546 443684 332590
rect 443748 304978 443776 339526
rect 443828 335096 443880 335102
rect 443828 335038 443880 335044
rect 443840 319802 443868 335038
rect 443920 335028 443972 335034
rect 443920 334970 443972 334976
rect 443932 322250 443960 334970
rect 444012 334892 444064 334898
rect 444012 334834 444064 334840
rect 443920 322244 443972 322250
rect 443920 322186 443972 322192
rect 444024 321842 444052 334834
rect 444116 331362 444144 444382
rect 444208 444378 444236 447170
rect 444196 444372 444248 444378
rect 444196 444314 444248 444320
rect 444194 422920 444250 422929
rect 444194 422855 444250 422864
rect 444104 331356 444156 331362
rect 444104 331298 444156 331304
rect 444012 321836 444064 321842
rect 444012 321778 444064 321784
rect 444208 320006 444236 422855
rect 444300 421977 444328 700402
rect 444380 444508 444432 444514
rect 444380 444450 444432 444456
rect 444286 421968 444342 421977
rect 444286 421903 444342 421912
rect 444288 331356 444340 331362
rect 444288 331298 444340 331304
rect 444196 320000 444248 320006
rect 444196 319942 444248 319948
rect 443828 319796 443880 319802
rect 443828 319738 443880 319744
rect 443736 304972 443788 304978
rect 443736 304914 443788 304920
rect 443644 194540 443696 194546
rect 443644 194482 443696 194488
rect 438596 161446 438808 161474
rect 441620 161492 441672 161498
rect 435272 160200 435324 160206
rect 435272 160142 435324 160148
rect 436008 160200 436060 160206
rect 436008 160142 436060 160148
rect 435284 159882 435312 160142
rect 438262 160132 438314 160138
rect 438262 160074 438314 160080
rect 431328 159854 431908 159882
rect 434824 159854 435312 159882
rect 438274 159882 438302 160074
rect 438596 159882 438624 161446
rect 441620 161434 441672 161440
rect 442908 161492 442960 161498
rect 442908 161434 442960 161440
rect 441632 160154 441660 161434
rect 444300 161430 444328 331298
rect 444392 330614 444420 444450
rect 444380 330608 444432 330614
rect 444380 330550 444432 330556
rect 445036 321502 445064 700674
rect 446404 700664 446456 700670
rect 446404 700606 446456 700612
rect 445116 700392 445168 700398
rect 445116 700334 445168 700340
rect 445024 321496 445076 321502
rect 445024 321438 445076 321444
rect 445128 320618 445156 700334
rect 445208 700324 445260 700330
rect 445208 700266 445260 700272
rect 445220 321745 445248 700266
rect 445390 683360 445446 683369
rect 445300 683324 445352 683330
rect 445390 683295 445446 683304
rect 445300 683266 445352 683272
rect 445206 321736 445262 321745
rect 445206 321671 445262 321680
rect 445116 320612 445168 320618
rect 445116 320554 445168 320560
rect 445312 319734 445340 683266
rect 445300 319728 445352 319734
rect 445300 319670 445352 319676
rect 445404 319326 445432 683295
rect 445484 683256 445536 683262
rect 445484 683198 445536 683204
rect 445496 321366 445524 683198
rect 446310 682816 446366 682825
rect 446310 682751 446366 682760
rect 445576 447160 445628 447166
rect 445576 447102 445628 447108
rect 445588 386578 445616 447102
rect 446220 444576 446272 444582
rect 446220 444518 446272 444524
rect 445666 387696 445722 387705
rect 445666 387631 445722 387640
rect 445576 386572 445628 386578
rect 445576 386514 445628 386520
rect 445588 354278 445616 386514
rect 445576 354272 445628 354278
rect 445576 354214 445628 354220
rect 445680 322046 445708 387631
rect 446232 344962 446260 444518
rect 446220 344956 446272 344962
rect 446220 344898 446272 344904
rect 446220 334960 446272 334966
rect 446220 334902 446272 334908
rect 445668 322040 445720 322046
rect 445668 321982 445720 321988
rect 446232 321978 446260 334902
rect 446220 321972 446272 321978
rect 446220 321914 446272 321920
rect 446324 321609 446352 682751
rect 446310 321600 446366 321609
rect 446310 321535 446366 321544
rect 445484 321360 445536 321366
rect 445484 321302 445536 321308
rect 446416 321094 446444 700606
rect 446496 686520 446548 686526
rect 446496 686462 446548 686468
rect 446404 321088 446456 321094
rect 446404 321030 446456 321036
rect 445392 319320 445444 319326
rect 445392 319262 445444 319268
rect 446508 319054 446536 686462
rect 446588 685228 446640 685234
rect 446588 685170 446640 685176
rect 446600 319705 446628 685170
rect 446772 685160 446824 685166
rect 446772 685102 446824 685108
rect 446680 683188 446732 683194
rect 446680 683130 446732 683136
rect 446586 319696 446642 319705
rect 446586 319631 446642 319640
rect 446692 319190 446720 683130
rect 446784 320113 446812 685102
rect 446956 684548 447008 684554
rect 446956 684490 447008 684496
rect 446862 683224 446918 683233
rect 446862 683159 446918 683168
rect 446770 320104 446826 320113
rect 446770 320039 446826 320048
rect 446680 319184 446732 319190
rect 446680 319126 446732 319132
rect 446876 319122 446904 683159
rect 446968 320686 446996 684490
rect 447048 682712 447100 682718
rect 447048 682654 447100 682660
rect 447060 320958 447088 682654
rect 447968 598256 448020 598262
rect 447968 598198 448020 598204
rect 447980 514457 448008 598198
rect 448060 522300 448112 522306
rect 448060 522242 448112 522248
rect 447966 514448 448022 514457
rect 447966 514383 448022 514392
rect 447414 512816 447470 512825
rect 447414 512751 447470 512760
rect 447428 499594 447456 512751
rect 447966 505200 448022 505209
rect 447966 505135 448022 505144
rect 447416 499588 447468 499594
rect 447416 499530 447468 499536
rect 447232 444372 447284 444378
rect 447232 444314 447284 444320
rect 447138 383616 447194 383625
rect 447138 383551 447140 383560
rect 447192 383551 447194 383560
rect 447140 383522 447192 383528
rect 447138 382256 447194 382265
rect 447138 382191 447194 382200
rect 447152 382158 447180 382191
rect 447140 382152 447192 382158
rect 447140 382094 447192 382100
rect 447138 380896 447194 380905
rect 447138 380831 447194 380840
rect 447152 380798 447180 380831
rect 447140 380792 447192 380798
rect 447140 380734 447192 380740
rect 447140 379432 447192 379438
rect 447140 379374 447192 379380
rect 447152 378865 447180 379374
rect 447138 378856 447194 378865
rect 447138 378791 447194 378800
rect 447140 378072 447192 378078
rect 447140 378014 447192 378020
rect 447152 377505 447180 378014
rect 447138 377496 447194 377505
rect 447138 377431 447194 377440
rect 447140 376712 447192 376718
rect 447140 376654 447192 376660
rect 447152 376145 447180 376654
rect 447138 376136 447194 376145
rect 447138 376071 447194 376080
rect 447140 375352 447192 375358
rect 447140 375294 447192 375300
rect 447152 374785 447180 375294
rect 447138 374776 447194 374785
rect 447138 374711 447194 374720
rect 447140 373992 447192 373998
rect 447140 373934 447192 373940
rect 447152 373425 447180 373934
rect 447138 373416 447194 373425
rect 447138 373351 447194 373360
rect 447140 372496 447192 372502
rect 447140 372438 447192 372444
rect 447152 372065 447180 372438
rect 447138 372056 447194 372065
rect 447138 371991 447194 372000
rect 447140 371136 447192 371142
rect 447140 371078 447192 371084
rect 447152 370705 447180 371078
rect 447138 370696 447194 370705
rect 447138 370631 447194 370640
rect 447140 369844 447192 369850
rect 447140 369786 447192 369792
rect 447152 369345 447180 369786
rect 447138 369336 447194 369345
rect 447138 369271 447194 369280
rect 447140 368416 447192 368422
rect 447140 368358 447192 368364
rect 447152 367985 447180 368358
rect 447138 367976 447194 367985
rect 447138 367911 447194 367920
rect 447140 367056 447192 367062
rect 447140 366998 447192 367004
rect 447152 365945 447180 366998
rect 447138 365936 447194 365945
rect 447138 365871 447194 365880
rect 447140 365696 447192 365702
rect 447140 365638 447192 365644
rect 447152 364585 447180 365638
rect 447138 364576 447194 364585
rect 447138 364511 447194 364520
rect 447138 363216 447194 363225
rect 447138 363151 447194 363160
rect 447152 363050 447180 363151
rect 447140 363044 447192 363050
rect 447140 362986 447192 362992
rect 447138 361856 447194 361865
rect 447138 361791 447194 361800
rect 447152 361622 447180 361791
rect 447140 361616 447192 361622
rect 447140 361558 447192 361564
rect 447138 361176 447194 361185
rect 447138 361111 447194 361120
rect 447152 360262 447180 361111
rect 447140 360256 447192 360262
rect 447140 360198 447192 360204
rect 447138 359136 447194 359145
rect 447138 359071 447194 359080
rect 447152 358834 447180 359071
rect 447140 358828 447192 358834
rect 447140 358770 447192 358776
rect 447138 350976 447194 350985
rect 447138 350911 447194 350920
rect 447152 350606 447180 350911
rect 447140 350600 447192 350606
rect 447140 350542 447192 350548
rect 447140 347744 447192 347750
rect 447140 347686 447192 347692
rect 447152 347585 447180 347686
rect 447138 347576 447194 347585
rect 447138 347511 447194 347520
rect 447244 342242 447272 444314
rect 447324 383648 447376 383654
rect 447324 383590 447376 383596
rect 447336 382945 447364 383590
rect 447322 382936 447378 382945
rect 447322 382871 447378 382880
rect 447324 382220 447376 382226
rect 447324 382162 447376 382168
rect 447336 381585 447364 382162
rect 447322 381576 447378 381585
rect 447322 381511 447378 381520
rect 447324 380724 447376 380730
rect 447324 380666 447376 380672
rect 447336 379545 447364 380666
rect 447322 379536 447378 379545
rect 447322 379471 447378 379480
rect 447324 378140 447376 378146
rect 447324 378082 447376 378088
rect 447336 376825 447364 378082
rect 447322 376816 447378 376825
rect 447322 376751 447378 376760
rect 447324 376644 447376 376650
rect 447324 376586 447376 376592
rect 447336 375465 447364 376586
rect 447322 375456 447378 375465
rect 447322 375391 447378 375400
rect 447324 375284 447376 375290
rect 447324 375226 447376 375232
rect 447336 374105 447364 375226
rect 447322 374096 447378 374105
rect 447322 374031 447378 374040
rect 447324 373924 447376 373930
rect 447324 373866 447376 373872
rect 447336 372745 447364 373866
rect 447322 372736 447378 372745
rect 447322 372671 447378 372680
rect 447324 372564 447376 372570
rect 447324 372506 447376 372512
rect 447336 371385 447364 372506
rect 447322 371376 447378 371385
rect 447322 371311 447378 371320
rect 447324 371204 447376 371210
rect 447324 371146 447376 371152
rect 447336 370025 447364 371146
rect 447322 370016 447378 370025
rect 447322 369951 447378 369960
rect 447324 369776 447376 369782
rect 447324 369718 447376 369724
rect 447336 368665 447364 369718
rect 447322 368656 447378 368665
rect 447322 368591 447378 368600
rect 447324 368484 447376 368490
rect 447324 368426 447376 368432
rect 447336 367305 447364 368426
rect 447322 367296 447378 367305
rect 447322 367231 447378 367240
rect 447324 366988 447376 366994
rect 447324 366930 447376 366936
rect 447336 366625 447364 366930
rect 447322 366616 447378 366625
rect 447322 366551 447378 366560
rect 447324 365628 447376 365634
rect 447324 365570 447376 365576
rect 447336 365265 447364 365570
rect 447322 365256 447378 365265
rect 447322 365191 447378 365200
rect 447322 363896 447378 363905
rect 447322 363831 447378 363840
rect 447336 362982 447364 363831
rect 447324 362976 447376 362982
rect 447324 362918 447376 362924
rect 447322 362536 447378 362545
rect 447322 362471 447378 362480
rect 447336 361690 447364 362471
rect 447324 361684 447376 361690
rect 447324 361626 447376 361632
rect 447322 360496 447378 360505
rect 447322 360431 447378 360440
rect 447336 360330 447364 360431
rect 447324 360324 447376 360330
rect 447324 360266 447376 360272
rect 447322 359816 447378 359825
rect 447322 359751 447378 359760
rect 447336 358902 447364 359751
rect 447324 358896 447376 358902
rect 447324 358838 447376 358844
rect 447324 354272 447376 354278
rect 447324 354214 447376 354220
rect 447336 344282 447364 354214
rect 447324 344276 447376 344282
rect 447324 344218 447376 344224
rect 447322 344176 447378 344185
rect 447322 344111 447378 344120
rect 447232 342236 447284 342242
rect 447232 342178 447284 342184
rect 447230 342136 447286 342145
rect 447230 342071 447286 342080
rect 447138 341456 447194 341465
rect 447138 341391 447194 341400
rect 447152 341018 447180 341391
rect 447140 341012 447192 341018
rect 447140 340954 447192 340960
rect 447244 340950 447272 342071
rect 447232 340944 447284 340950
rect 447232 340886 447284 340892
rect 447138 340776 447194 340785
rect 447138 340711 447194 340720
rect 447152 339522 447180 340711
rect 447230 340096 447286 340105
rect 447230 340031 447286 340040
rect 447244 339590 447272 340031
rect 447232 339584 447284 339590
rect 447232 339526 447284 339532
rect 447140 339516 447192 339522
rect 447140 339458 447192 339464
rect 447230 339416 447286 339425
rect 447230 339351 447286 339360
rect 447138 338736 447194 338745
rect 447138 338671 447194 338680
rect 447152 338230 447180 338671
rect 447140 338224 447192 338230
rect 447140 338166 447192 338172
rect 447244 338162 447272 339351
rect 447232 338156 447284 338162
rect 447232 338098 447284 338104
rect 447230 338056 447286 338065
rect 447230 337991 447286 338000
rect 447138 337376 447194 337385
rect 447138 337311 447194 337320
rect 447152 336802 447180 337311
rect 447244 336870 447272 337991
rect 447232 336864 447284 336870
rect 447232 336806 447284 336812
rect 447140 336796 447192 336802
rect 447140 336738 447192 336744
rect 447230 336696 447286 336705
rect 447230 336631 447286 336640
rect 447138 336016 447194 336025
rect 447138 335951 447194 335960
rect 447152 335442 447180 335951
rect 447140 335436 447192 335442
rect 447140 335378 447192 335384
rect 447244 335374 447272 336631
rect 447232 335368 447284 335374
rect 447232 335310 447284 335316
rect 447230 334656 447286 334665
rect 447230 334591 447286 334600
rect 447244 334014 447272 334591
rect 447232 334008 447284 334014
rect 447138 333976 447194 333985
rect 447232 333950 447284 333956
rect 447138 333911 447194 333920
rect 447152 332858 447180 333911
rect 447230 333296 447286 333305
rect 447230 333231 447286 333240
rect 447140 332852 447192 332858
rect 447140 332794 447192 332800
rect 447244 332654 447272 333231
rect 447232 332648 447284 332654
rect 447232 332590 447284 332596
rect 447138 331936 447194 331945
rect 447138 331871 447194 331880
rect 447152 331294 447180 331871
rect 447232 331356 447284 331362
rect 447232 331298 447284 331304
rect 447140 331288 447192 331294
rect 447244 331265 447272 331298
rect 447140 331230 447192 331236
rect 447230 331256 447286 331265
rect 447230 331191 447286 331200
rect 447140 330608 447192 330614
rect 447138 330576 447140 330585
rect 447192 330576 447194 330585
rect 447138 330511 447194 330520
rect 447138 329216 447194 329225
rect 447138 329151 447194 329160
rect 447152 328506 447180 329151
rect 447140 328500 447192 328506
rect 447140 328442 447192 328448
rect 447048 320952 447100 320958
rect 447048 320894 447100 320900
rect 446956 320680 447008 320686
rect 446956 320622 447008 320628
rect 446864 319116 446916 319122
rect 446864 319058 446916 319064
rect 446496 319048 446548 319054
rect 446496 318990 446548 318996
rect 446404 304496 446456 304502
rect 446404 304438 446456 304444
rect 446416 289678 446444 304438
rect 446404 289672 446456 289678
rect 446404 289614 446456 289620
rect 445024 288380 445076 288386
rect 445024 288322 445076 288328
rect 445036 262886 445064 288322
rect 445668 268592 445720 268598
rect 445668 268534 445720 268540
rect 445680 264246 445708 268534
rect 445668 264240 445720 264246
rect 445668 264182 445720 264188
rect 445024 262880 445076 262886
rect 445024 262822 445076 262828
rect 447336 171134 447364 344111
rect 447428 334150 447456 499530
rect 447980 499526 448008 505135
rect 448072 501945 448100 522242
rect 448336 518220 448388 518226
rect 448336 518162 448388 518168
rect 448150 516760 448206 516769
rect 448150 516695 448206 516704
rect 448164 507793 448192 516695
rect 448348 512825 448376 518162
rect 448428 516180 448480 516186
rect 448428 516122 448480 516128
rect 448334 512816 448390 512825
rect 448334 512751 448390 512760
rect 448440 510513 448468 516122
rect 448518 514448 448574 514457
rect 448518 514383 448574 514392
rect 448426 510504 448482 510513
rect 448256 510462 448426 510490
rect 448150 507784 448206 507793
rect 448150 507719 448206 507728
rect 448058 501936 448114 501945
rect 448058 501871 448114 501880
rect 448060 501832 448112 501838
rect 448060 501774 448112 501780
rect 447968 499520 448020 499526
rect 447968 499462 448020 499468
rect 447876 387184 447928 387190
rect 447876 387126 447928 387132
rect 447784 385416 447836 385422
rect 447784 385358 447836 385364
rect 447508 380860 447560 380866
rect 447508 380802 447560 380808
rect 447520 380225 447548 380802
rect 447506 380216 447562 380225
rect 447506 380151 447562 380160
rect 447508 379500 447560 379506
rect 447508 379442 447560 379448
rect 447520 378185 447548 379442
rect 447506 378176 447562 378185
rect 447506 378111 447562 378120
rect 447796 352345 447824 385358
rect 447888 353705 447916 387126
rect 447874 353696 447930 353705
rect 447874 353631 447930 353640
rect 447782 352336 447838 352345
rect 447782 352271 447838 352280
rect 447508 344276 447560 344282
rect 447508 344218 447560 344224
rect 447520 343505 447548 344218
rect 447506 343496 447562 343505
rect 447506 343431 447562 343440
rect 447520 342922 447548 343431
rect 447508 342916 447560 342922
rect 447508 342858 447560 342864
rect 447600 342236 447652 342242
rect 447600 342178 447652 342184
rect 447506 335336 447562 335345
rect 447506 335271 447562 335280
rect 447416 334144 447468 334150
rect 447416 334086 447468 334092
rect 447428 332874 447456 334086
rect 447520 334082 447548 335271
rect 447508 334076 447560 334082
rect 447508 334018 447560 334024
rect 447428 332846 447548 332874
rect 447416 332784 447468 332790
rect 447416 332726 447468 332732
rect 447428 332625 447456 332726
rect 447414 332616 447470 332625
rect 447414 332551 447470 332560
rect 447416 329112 447468 329118
rect 447416 329054 447468 329060
rect 447428 328545 447456 329054
rect 447414 328536 447470 328545
rect 447414 328471 447470 328480
rect 447520 327865 447548 332846
rect 447612 330546 447640 342178
rect 447600 330540 447652 330546
rect 447600 330482 447652 330488
rect 447612 329905 447640 330482
rect 447598 329896 447654 329905
rect 447598 329831 447654 329840
rect 447506 327856 447562 327865
rect 447506 327791 447562 327800
rect 447416 327072 447468 327078
rect 447416 327014 447468 327020
rect 447428 326505 447456 327014
rect 447980 327010 448008 499462
rect 448072 499458 448100 501774
rect 448060 499452 448112 499458
rect 448060 499394 448112 499400
rect 447968 327004 448020 327010
rect 447968 326946 448020 326952
rect 447414 326496 447470 326505
rect 447414 326431 447470 326440
rect 447980 325825 448008 326946
rect 447966 325816 448022 325825
rect 447966 325751 448022 325760
rect 447784 305584 447836 305590
rect 447784 305526 447836 305532
rect 447796 288386 447824 305526
rect 447784 288380 447836 288386
rect 447784 288322 447836 288328
rect 447784 268524 447836 268530
rect 447784 268466 447836 268472
rect 447796 240786 447824 268466
rect 447980 265674 448008 325751
rect 448072 325582 448100 499394
rect 448164 327078 448192 507719
rect 448256 328438 448284 510462
rect 448426 510439 448482 510448
rect 448532 509234 448560 514383
rect 448440 509206 448560 509234
rect 448334 503432 448390 503441
rect 448334 503367 448390 503376
rect 448348 501838 448376 503367
rect 448336 501832 448388 501838
rect 448336 501774 448388 501780
rect 448440 500290 448468 509206
rect 448440 500274 448560 500290
rect 448440 500268 448572 500274
rect 448440 500262 448520 500268
rect 448440 489914 448468 500262
rect 448520 500210 448572 500216
rect 448348 489886 448468 489914
rect 448348 328545 448376 489886
rect 448980 387116 449032 387122
rect 448980 387058 449032 387064
rect 448428 386028 448480 386034
rect 448428 385970 448480 385976
rect 448440 358465 448468 385970
rect 448426 358456 448482 358465
rect 448426 358391 448482 358400
rect 448992 357785 449020 387058
rect 449070 387016 449126 387025
rect 449070 386951 449126 386960
rect 448978 357776 449034 357785
rect 448978 357711 449034 357720
rect 449084 355745 449112 386951
rect 449070 355736 449126 355745
rect 449070 355671 449126 355680
rect 448428 344956 448480 344962
rect 448428 344898 448480 344904
rect 448440 344865 448468 344898
rect 448426 344856 448482 344865
rect 448426 344791 448482 344800
rect 449072 334824 449124 334830
rect 449072 334766 449124 334772
rect 448426 332616 448482 332625
rect 448426 332551 448482 332560
rect 448334 328536 448390 328545
rect 448334 328471 448390 328480
rect 448244 328432 448296 328438
rect 448244 328374 448296 328380
rect 448256 327185 448284 328374
rect 448242 327176 448298 327185
rect 448242 327111 448298 327120
rect 448152 327072 448204 327078
rect 448152 327014 448204 327020
rect 448060 325576 448112 325582
rect 448060 325518 448112 325524
rect 448072 325122 448100 325518
rect 448242 325136 448298 325145
rect 448072 325094 448242 325122
rect 448242 325071 448298 325080
rect 448256 318102 448284 325071
rect 448336 324964 448388 324970
rect 448336 324906 448388 324912
rect 448244 318096 448296 318102
rect 448244 318038 448296 318044
rect 447968 265668 448020 265674
rect 447968 265610 448020 265616
rect 447784 240780 447836 240786
rect 447784 240722 447836 240728
rect 448348 207670 448376 324906
rect 448336 207664 448388 207670
rect 448336 207606 448388 207612
rect 447336 171106 447824 171134
rect 445208 163124 445260 163130
rect 445208 163066 445260 163072
rect 444288 161424 444340 161430
rect 444288 161366 444340 161372
rect 444300 160750 444328 161366
rect 444288 160744 444340 160750
rect 444288 160686 444340 160692
rect 438274 159868 438624 159882
rect 441586 160126 441660 160154
rect 445220 160138 445248 163066
rect 444886 160132 444938 160138
rect 441586 159868 441614 160126
rect 444886 160074 444938 160080
rect 445208 160132 445260 160138
rect 445208 160074 445260 160080
rect 444898 159868 444926 160074
rect 447796 159882 447824 171106
rect 448440 163538 448468 332551
rect 449084 321910 449112 334766
rect 449072 321904 449124 321910
rect 449072 321846 449124 321852
rect 449176 321706 449204 700742
rect 450544 700596 450596 700602
rect 450544 700538 450596 700544
rect 449256 700528 449308 700534
rect 449256 700470 449308 700476
rect 449268 322182 449296 700470
rect 449348 687948 449400 687954
rect 449348 687890 449400 687896
rect 449256 322176 449308 322182
rect 449256 322118 449308 322124
rect 449164 321700 449216 321706
rect 449164 321642 449216 321648
rect 449360 320074 449388 687890
rect 449808 595468 449860 595474
rect 449808 595410 449860 595416
rect 449820 503441 449848 595410
rect 449992 520396 450044 520402
rect 449992 520338 450044 520344
rect 449806 503432 449862 503441
rect 449806 503367 449862 503376
rect 449716 499588 449768 499594
rect 449716 499530 449768 499536
rect 449728 498846 449756 499530
rect 449716 498840 449768 498846
rect 449716 498782 449768 498788
rect 449900 496120 449952 496126
rect 449898 496088 449900 496097
rect 449952 496088 449954 496097
rect 449898 496023 449954 496032
rect 449900 494760 449952 494766
rect 449900 494702 449952 494708
rect 449808 457496 449860 457502
rect 449808 457438 449860 457444
rect 449716 454776 449768 454782
rect 449716 454718 449768 454724
rect 449624 454708 449676 454714
rect 449624 454650 449676 454656
rect 449438 387152 449494 387161
rect 449438 387087 449494 387096
rect 449452 354385 449480 387087
rect 449530 385656 449586 385665
rect 449530 385591 449586 385600
rect 449438 354376 449494 354385
rect 449438 354311 449494 354320
rect 449440 336116 449492 336122
rect 449440 336058 449492 336064
rect 449348 320068 449400 320074
rect 449348 320010 449400 320016
rect 449452 319870 449480 336058
rect 449544 324970 449572 385591
rect 449636 356425 449664 454650
rect 449622 356416 449678 356425
rect 449622 356351 449678 356360
rect 449728 355065 449756 454718
rect 449820 357105 449848 457438
rect 449912 389298 449940 494702
rect 449900 389292 449952 389298
rect 449900 389234 449952 389240
rect 449806 357096 449862 357105
rect 449806 357031 449862 357040
rect 449714 355056 449770 355065
rect 449714 354991 449770 355000
rect 449898 351112 449954 351121
rect 449898 351047 449954 351056
rect 449714 350296 449770 350305
rect 449714 350231 449770 350240
rect 449622 345536 449678 345545
rect 449622 345471 449678 345480
rect 449532 324964 449584 324970
rect 449532 324906 449584 324912
rect 449544 324465 449572 324906
rect 449530 324456 449586 324465
rect 449530 324391 449586 324400
rect 449440 319864 449492 319870
rect 449440 319806 449492 319812
rect 449636 307154 449664 345471
rect 449624 307148 449676 307154
rect 449624 307090 449676 307096
rect 449728 263566 449756 350231
rect 449806 343496 449862 343505
rect 449806 343431 449862 343440
rect 449716 263560 449768 263566
rect 449716 263502 449768 263508
rect 449820 249762 449848 343431
rect 449808 249756 449860 249762
rect 449808 249698 449860 249704
rect 448428 163532 448480 163538
rect 448428 163474 448480 163480
rect 438288 159854 438624 159868
rect 447796 159854 448224 159882
rect 425040 159718 425192 159746
rect 434824 159390 434852 159854
rect 434812 159384 434864 159390
rect 434812 159326 434864 159332
rect 410708 139392 410760 139398
rect 410708 139334 410760 139340
rect 410616 95192 410668 95198
rect 410616 95134 410668 95140
rect 410524 73160 410576 73166
rect 410524 73102 410576 73108
rect 449912 62830 449940 351047
rect 450004 350033 450032 520338
rect 450084 464364 450136 464370
rect 450084 464306 450136 464312
rect 449990 350024 450046 350033
rect 449990 349959 450046 349968
rect 450096 346361 450124 464306
rect 450176 460964 450228 460970
rect 450176 460906 450228 460912
rect 450188 347313 450216 460906
rect 450268 454844 450320 454850
rect 450268 454786 450320 454792
rect 450280 353297 450308 454786
rect 450360 385144 450412 385150
rect 450360 385086 450412 385092
rect 450266 353288 450322 353297
rect 450266 353223 450322 353232
rect 450372 348673 450400 385086
rect 450358 348664 450414 348673
rect 450358 348599 450414 348608
rect 450174 347304 450230 347313
rect 450174 347239 450230 347248
rect 450082 346352 450138 346361
rect 450082 346287 450138 346296
rect 450452 334756 450504 334762
rect 450452 334698 450504 334704
rect 450464 322386 450492 334698
rect 450452 322380 450504 322386
rect 450452 322322 450504 322328
rect 450556 321434 450584 700538
rect 462332 669905 462360 703520
rect 478524 700505 478552 703520
rect 478510 700496 478566 700505
rect 478510 700431 478566 700440
rect 494808 700369 494836 703520
rect 494794 700360 494850 700369
rect 494794 700295 494850 700304
rect 527192 699825 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 462318 669896 462374 669905
rect 462318 669831 462374 669840
rect 457810 667992 457866 668001
rect 457810 667927 457866 667936
rect 457718 653304 457774 653313
rect 457718 653239 457774 653248
rect 457626 650856 457682 650865
rect 457626 650791 457682 650800
rect 457534 645960 457590 645969
rect 457534 645895 457590 645904
rect 457442 621480 457498 621489
rect 457442 621415 457498 621424
rect 457350 616584 457406 616593
rect 457350 616519 457406 616528
rect 457258 609240 457314 609249
rect 457258 609175 457314 609184
rect 457272 599690 457300 609175
rect 457260 599684 457312 599690
rect 457260 599626 457312 599632
rect 457364 543046 457392 616519
rect 457456 595542 457484 621415
rect 457548 600234 457576 645895
rect 457536 600228 457588 600234
rect 457536 600170 457588 600176
rect 457640 598330 457668 650791
rect 457628 598324 457680 598330
rect 457628 598266 457680 598272
rect 457732 596630 457760 653239
rect 457824 600302 457852 667927
rect 458086 660648 458142 660657
rect 458086 660583 458142 660592
rect 457994 658200 458050 658209
rect 457994 658135 458050 658144
rect 457902 641064 457958 641073
rect 457902 640999 457958 641008
rect 457812 600296 457864 600302
rect 457812 600238 457864 600244
rect 457916 599622 457944 640999
rect 457904 599616 457956 599622
rect 457904 599558 457956 599564
rect 457720 596624 457772 596630
rect 457720 596566 457772 596572
rect 457444 595536 457496 595542
rect 457444 595478 457496 595484
rect 457352 543040 457404 543046
rect 457352 542982 457404 542988
rect 458008 523734 458036 658135
rect 457996 523728 458048 523734
rect 457996 523670 458048 523676
rect 458100 522374 458128 660583
rect 459190 655752 459246 655761
rect 459190 655687 459246 655696
rect 459098 648408 459154 648417
rect 459098 648343 459154 648352
rect 459006 643512 459062 643521
rect 459006 643447 459062 643456
rect 458914 638616 458970 638625
rect 458914 638551 458970 638560
rect 458822 619032 458878 619041
rect 458822 618967 458878 618976
rect 458638 611688 458694 611697
rect 458638 611623 458694 611632
rect 458652 599758 458680 611623
rect 458732 602812 458784 602818
rect 458732 602754 458784 602760
rect 458640 599752 458692 599758
rect 458640 599694 458692 599700
rect 458744 596873 458772 602754
rect 458836 598398 458864 618967
rect 458824 598392 458876 598398
rect 458824 598334 458876 598340
rect 458928 598233 458956 638551
rect 458914 598224 458970 598233
rect 458914 598159 458970 598168
rect 459020 597009 459048 643447
rect 459112 602818 459140 648343
rect 459100 602812 459152 602818
rect 459100 602754 459152 602760
rect 459204 602698 459232 655687
rect 459466 631272 459522 631281
rect 459466 631207 459522 631216
rect 459282 628824 459338 628833
rect 459282 628759 459338 628768
rect 459112 602670 459232 602698
rect 459112 599593 459140 602670
rect 459190 601896 459246 601905
rect 459190 601831 459246 601840
rect 459204 600030 459232 601831
rect 459192 600024 459244 600030
rect 459192 599966 459244 599972
rect 459098 599584 459154 599593
rect 459098 599519 459154 599528
rect 459006 597000 459062 597009
rect 459006 596935 459062 596944
rect 458730 596864 458786 596873
rect 458730 596799 458786 596808
rect 458088 522368 458140 522374
rect 458088 522310 458140 522316
rect 459296 520946 459324 628759
rect 459374 626376 459430 626385
rect 459374 626311 459430 626320
rect 459284 520940 459336 520946
rect 459284 520882 459336 520888
rect 450636 519580 450688 519586
rect 450636 519522 450688 519528
rect 450648 516361 450676 519522
rect 459388 518294 459416 626311
rect 459480 522345 459508 631207
rect 459558 623860 459614 623869
rect 459558 623795 459614 623804
rect 459572 536110 459600 623795
rect 459650 614136 459706 614145
rect 459650 614071 459706 614080
rect 459664 594114 459692 614071
rect 459742 606724 459798 606733
rect 459742 606659 459798 606668
rect 459756 596902 459784 606659
rect 459834 604276 459890 604285
rect 459834 604211 459890 604220
rect 459848 598466 459876 604211
rect 461676 600296 461728 600302
rect 461676 600238 461728 600244
rect 461584 600228 461636 600234
rect 461584 600170 461636 600176
rect 459836 598460 459888 598466
rect 459836 598402 459888 598408
rect 459744 596896 459796 596902
rect 459744 596838 459796 596844
rect 459652 594108 459704 594114
rect 459652 594050 459704 594056
rect 459560 536104 459612 536110
rect 459560 536046 459612 536052
rect 459466 522336 459522 522345
rect 459466 522271 459522 522280
rect 459376 518288 459428 518294
rect 459376 518230 459428 518236
rect 450634 516352 450690 516361
rect 450634 516287 450690 516296
rect 450648 500126 450754 500154
rect 451292 500126 452226 500154
rect 450648 494766 450676 500126
rect 450636 494760 450688 494766
rect 450636 494702 450688 494708
rect 450636 455524 450688 455530
rect 450636 455466 450688 455472
rect 450648 349081 450676 455466
rect 450728 389292 450780 389298
rect 450728 389234 450780 389240
rect 450740 385914 450768 389234
rect 451292 385914 451320 500126
rect 453304 497548 453356 497554
rect 453304 497490 453356 497496
rect 451924 497480 451976 497486
rect 451924 497422 451976 497428
rect 451372 496868 451424 496874
rect 451372 496810 451424 496816
rect 451384 402974 451412 496810
rect 451384 402946 451872 402974
rect 451844 385914 451872 402946
rect 451936 386034 451964 497422
rect 452844 496936 452896 496942
rect 452844 496878 452896 496884
rect 451924 386028 451976 386034
rect 451924 385970 451976 385976
rect 452856 385914 452884 496878
rect 450740 385886 450846 385914
rect 451292 385886 451582 385914
rect 451844 385886 452318 385914
rect 452856 385886 453054 385914
rect 453316 385422 453344 497490
rect 453684 496874 453712 500140
rect 454132 497072 454184 497078
rect 454132 497014 454184 497020
rect 454040 497004 454092 497010
rect 454040 496946 454092 496952
rect 453672 496868 453724 496874
rect 453672 496810 453724 496816
rect 453764 389156 453816 389162
rect 453764 389098 453816 389104
rect 453776 385900 453804 389098
rect 454052 385914 454080 496946
rect 454144 402974 454172 497014
rect 455156 496942 455184 500140
rect 455144 496936 455196 496942
rect 455144 496878 455196 496884
rect 455420 496936 455472 496942
rect 455420 496878 455472 496884
rect 454684 496868 454736 496874
rect 454684 496810 454736 496816
rect 454144 402946 454632 402974
rect 454604 386050 454632 402946
rect 454696 389162 454724 496810
rect 455432 402974 455460 496878
rect 456628 496874 456656 500140
rect 457444 497616 457496 497622
rect 457444 497558 457496 497564
rect 456616 496868 456668 496874
rect 456616 496810 456668 496816
rect 456892 429888 456944 429894
rect 456892 429830 456944 429836
rect 456904 402974 456932 429830
rect 455432 402946 455552 402974
rect 456904 402946 457024 402974
rect 454684 389156 454736 389162
rect 454684 389098 454736 389104
rect 454604 386022 454816 386050
rect 454788 385914 454816 386022
rect 455524 385914 455552 402946
rect 456708 388884 456760 388890
rect 456708 388826 456760 388832
rect 454052 385886 454526 385914
rect 454788 385886 455262 385914
rect 455524 385886 455998 385914
rect 456720 385900 456748 388826
rect 456996 385914 457024 402946
rect 457456 387190 457484 497558
rect 458100 497010 458128 500140
rect 459572 497078 459600 500140
rect 459560 497072 459612 497078
rect 459560 497014 459612 497020
rect 458088 497004 458140 497010
rect 458088 496946 458140 496952
rect 461044 496942 461072 500140
rect 461032 496936 461084 496942
rect 461032 496878 461084 496884
rect 457536 428460 457588 428466
rect 457536 428402 457588 428408
rect 457548 388890 457576 428402
rect 459928 398132 459980 398138
rect 459928 398074 459980 398080
rect 458456 396772 458508 396778
rect 458456 396714 458508 396720
rect 458180 395344 458232 395350
rect 458180 395286 458232 395292
rect 457536 388884 457588 388890
rect 457536 388826 457588 388832
rect 457444 387184 457496 387190
rect 457444 387126 457496 387132
rect 456996 385886 457470 385914
rect 458192 385900 458220 395286
rect 458468 385914 458496 396714
rect 459652 391332 459704 391338
rect 459652 391274 459704 391280
rect 458468 385886 458942 385914
rect 459664 385900 459692 391274
rect 459940 385914 459968 398074
rect 461124 389836 461176 389842
rect 461124 389778 461176 389784
rect 459940 385886 460414 385914
rect 461136 385900 461164 389778
rect 461596 388618 461624 600170
rect 461688 389162 461716 600238
rect 462424 600086 463542 600114
rect 469232 600086 470534 600114
rect 461768 596624 461820 596630
rect 461768 596566 461820 596572
rect 461676 389156 461728 389162
rect 461676 389098 461728 389104
rect 461584 388612 461636 388618
rect 461584 388554 461636 388560
rect 461780 388550 461808 596566
rect 462424 522306 462452 600086
rect 462504 600024 462556 600030
rect 462504 599966 462556 599972
rect 462412 522300 462464 522306
rect 462412 522242 462464 522248
rect 462516 402974 462544 599966
rect 465080 599752 465132 599758
rect 465080 599694 465132 599700
rect 463700 598460 463752 598466
rect 463700 598402 463752 598408
rect 462962 517576 463018 517585
rect 462962 517511 463018 517520
rect 462516 402946 462912 402974
rect 462596 389156 462648 389162
rect 462596 389098 462648 389104
rect 461860 389088 461912 389094
rect 461860 389030 461912 389036
rect 461768 388544 461820 388550
rect 461768 388486 461820 388492
rect 461872 385900 461900 389030
rect 462608 385900 462636 389098
rect 462884 385914 462912 402946
rect 462976 388482 463004 517511
rect 462964 388476 463016 388482
rect 462964 388418 463016 388424
rect 463712 385914 463740 598402
rect 463792 596896 463844 596902
rect 463792 596838 463844 596844
rect 463804 402974 463832 596838
rect 464344 595536 464396 595542
rect 464344 595478 464396 595484
rect 463804 402946 464292 402974
rect 464264 386050 464292 402946
rect 464356 389162 464384 595478
rect 465092 389298 465120 599694
rect 465172 599684 465224 599690
rect 465172 599626 465224 599632
rect 465080 389292 465132 389298
rect 465080 389234 465132 389240
rect 464344 389156 464396 389162
rect 464344 389098 464396 389104
rect 464264 386022 464384 386050
rect 464356 385914 464384 386022
rect 465184 385914 465212 599626
rect 468484 599616 468536 599622
rect 468484 599558 468536 599564
rect 467932 598392 467984 598398
rect 467932 598334 467984 598340
rect 466460 594108 466512 594114
rect 466460 594050 466512 594056
rect 465540 393984 465592 393990
rect 465540 393926 465592 393932
rect 465552 389094 465580 393926
rect 465908 389292 465960 389298
rect 465908 389234 465960 389240
rect 465540 389088 465592 389094
rect 465540 389030 465592 389036
rect 465920 385914 465948 389234
rect 466472 385914 466500 594050
rect 466552 543040 466604 543046
rect 466552 542982 466604 542988
rect 466564 402974 466592 542982
rect 467104 523728 467156 523734
rect 467104 523670 467156 523676
rect 466564 402946 467052 402974
rect 467024 386730 467052 402946
rect 467116 388754 467144 523670
rect 467194 519480 467250 519489
rect 467194 519415 467250 519424
rect 467104 388748 467156 388754
rect 467104 388690 467156 388696
rect 467208 388686 467236 519415
rect 467944 402974 467972 598334
rect 467944 402946 468064 402974
rect 467196 388680 467248 388686
rect 467196 388622 467248 388628
rect 467024 386702 467328 386730
rect 467300 385914 467328 386702
rect 468036 385914 468064 402946
rect 468496 388958 468524 599558
rect 468576 598324 468628 598330
rect 468576 598266 468628 598272
rect 468484 388952 468536 388958
rect 468484 388894 468536 388900
rect 468588 388822 468616 598266
rect 469232 595474 469260 600086
rect 477512 598330 477540 600100
rect 484504 598398 484532 600100
rect 484492 598392 484544 598398
rect 484492 598334 484544 598340
rect 477500 598324 477552 598330
rect 477500 598266 477552 598272
rect 491496 597854 491524 600100
rect 498212 600086 498502 600114
rect 494152 598392 494204 598398
rect 494152 598334 494204 598340
rect 494060 598324 494112 598330
rect 494060 598266 494112 598272
rect 491484 597848 491536 597854
rect 491484 597790 491536 597796
rect 469220 595468 469272 595474
rect 469220 595410 469272 595416
rect 469404 536104 469456 536110
rect 469404 536046 469456 536052
rect 468668 522368 468720 522374
rect 468668 522310 468720 522316
rect 468680 388890 468708 522310
rect 469416 402974 469444 536046
rect 470876 520940 470928 520946
rect 470876 520882 470928 520888
rect 482928 520940 482980 520946
rect 482928 520882 482980 520888
rect 470692 518288 470744 518294
rect 470692 518230 470744 518236
rect 469416 402946 469536 402974
rect 469220 389156 469272 389162
rect 469220 389098 469272 389104
rect 468668 388884 468720 388890
rect 468668 388826 468720 388832
rect 468576 388816 468628 388822
rect 468576 388758 468628 388764
rect 462884 385886 463358 385914
rect 463712 385886 464094 385914
rect 464356 385886 464830 385914
rect 465184 385886 465566 385914
rect 465920 385886 466302 385914
rect 466472 385886 467038 385914
rect 467300 385886 467774 385914
rect 468036 385886 468510 385914
rect 469232 385900 469260 389098
rect 469508 385914 469536 402946
rect 469508 385886 469982 385914
rect 470704 385900 470732 518230
rect 470888 402974 470916 520882
rect 482940 517562 482968 520882
rect 488632 520396 488684 520402
rect 488632 520338 488684 520344
rect 488644 517970 488672 520338
rect 488644 517942 488980 517970
rect 482664 517546 483000 517562
rect 480168 517540 480220 517546
rect 480168 517482 480220 517488
rect 482652 517540 483000 517546
rect 482704 517534 483000 517540
rect 482652 517482 482704 517488
rect 480180 461650 480208 517482
rect 491850 516216 491906 516225
rect 491850 516151 491852 516160
rect 491904 516151 491906 516160
rect 491852 516122 491904 516128
rect 494072 508881 494100 598266
rect 494164 516769 494192 598334
rect 494244 597848 494296 597854
rect 494244 597790 494296 597796
rect 494150 516760 494206 516769
rect 494150 516695 494206 516704
rect 494150 515944 494206 515953
rect 494256 515930 494284 597790
rect 498212 518226 498240 600086
rect 505480 598262 505508 600100
rect 512012 600086 512486 600114
rect 518912 600086 519478 600114
rect 525812 600086 526470 600114
rect 505468 598256 505520 598262
rect 505468 598198 505520 598204
rect 511264 590708 511316 590714
rect 511264 590650 511316 590656
rect 498200 518220 498252 518226
rect 498200 518162 498252 518168
rect 494334 516760 494390 516769
rect 494334 516695 494390 516704
rect 494206 515902 494284 515930
rect 494150 515879 494206 515888
rect 494164 515438 494192 515879
rect 494152 515432 494204 515438
rect 494152 515374 494204 515380
rect 494348 512650 494376 516695
rect 494152 512644 494204 512650
rect 494152 512586 494204 512592
rect 494336 512644 494388 512650
rect 494336 512586 494388 512592
rect 494164 512553 494192 512586
rect 494150 512544 494206 512553
rect 494150 512479 494206 512488
rect 494058 508872 494114 508881
rect 494058 508807 494114 508816
rect 494072 507890 494100 508807
rect 494060 507884 494112 507890
rect 494060 507826 494112 507832
rect 480272 500126 480608 500154
rect 481744 500126 481804 500154
rect 482664 500126 483000 500154
rect 483860 500126 484196 500154
rect 484412 500126 485392 500154
rect 486436 500126 486588 500154
rect 487172 500126 487784 500154
rect 488552 500126 488980 500154
rect 490176 500126 491156 500154
rect 480272 497554 480300 500126
rect 480260 497548 480312 497554
rect 480260 497490 480312 497496
rect 480168 461644 480220 461650
rect 480168 461586 480220 461592
rect 480180 456822 480208 461586
rect 473728 456816 473780 456822
rect 473728 456758 473780 456764
rect 480168 456816 480220 456822
rect 480168 456758 480220 456764
rect 473740 455462 473768 456758
rect 480996 455524 481048 455530
rect 480996 455466 481048 455472
rect 473728 455456 473780 455462
rect 473728 455398 473780 455404
rect 473740 453900 473768 455398
rect 481008 453900 481036 455466
rect 481744 454850 481772 500126
rect 482664 497622 482692 500126
rect 482652 497616 482704 497622
rect 482652 497558 482704 497564
rect 483860 496913 483888 500126
rect 483846 496904 483902 496913
rect 483846 496839 483902 496848
rect 481732 454844 481784 454850
rect 481732 454786 481784 454792
rect 484412 454782 484440 500126
rect 486436 496913 486464 500126
rect 486422 496904 486478 496913
rect 486422 496839 486478 496848
rect 484400 454776 484452 454782
rect 484400 454718 484452 454724
rect 487172 454714 487200 500126
rect 488552 457502 488580 500126
rect 488540 457496 488592 457502
rect 488540 457438 488592 457444
rect 488264 456068 488316 456074
rect 488264 456010 488316 456016
rect 487160 454708 487212 454714
rect 487160 454650 487212 454656
rect 487986 453928 488042 453937
rect 488276 453914 488304 456010
rect 488042 453900 488304 453914
rect 488042 453886 488290 453900
rect 487986 453863 488042 453872
rect 471624 428466 471652 432140
rect 474292 429894 474320 432140
rect 476132 432126 476974 432154
rect 478892 432126 479642 432154
rect 474280 429888 474332 429894
rect 474280 429830 474332 429836
rect 471612 428460 471664 428466
rect 471612 428402 471664 428408
rect 470888 402946 471008 402974
rect 470980 385914 471008 402946
rect 476132 395350 476160 432126
rect 478892 396778 478920 432126
rect 482296 429214 482324 432140
rect 484964 429214 484992 432140
rect 487632 429214 487660 432140
rect 490024 432126 490314 432154
rect 480904 429208 480956 429214
rect 480904 429150 480956 429156
rect 482284 429208 482336 429214
rect 482284 429150 482336 429156
rect 483664 429208 483716 429214
rect 483664 429150 483716 429156
rect 484952 429208 485004 429214
rect 484952 429150 485004 429156
rect 486424 429208 486476 429214
rect 486424 429150 486476 429156
rect 487620 429208 487672 429214
rect 487620 429150 487672 429156
rect 478880 396772 478932 396778
rect 478880 396714 478932 396720
rect 476120 395344 476172 395350
rect 476120 395286 476172 395292
rect 473358 393952 473414 393961
rect 473358 393887 473414 393896
rect 472898 392592 472954 392601
rect 472898 392527 472954 392536
rect 472162 389056 472218 389065
rect 472162 388991 472218 389000
rect 470980 385886 471454 385914
rect 472176 385900 472204 388991
rect 472912 385900 472940 392527
rect 473372 385914 473400 393887
rect 480916 391338 480944 429150
rect 483020 421592 483072 421598
rect 483020 421534 483072 421540
rect 480904 391332 480956 391338
rect 480904 391274 480956 391280
rect 474370 389056 474426 389065
rect 474370 388991 474426 389000
rect 475842 389056 475898 389065
rect 475842 388991 475898 389000
rect 477314 389056 477370 389065
rect 477314 388991 477370 389000
rect 479522 389056 479578 389065
rect 479522 388991 479578 389000
rect 473372 385886 473662 385914
rect 474384 385900 474412 388991
rect 475108 388952 475160 388958
rect 475108 388894 475160 388900
rect 475120 385900 475148 388894
rect 475856 385900 475884 388991
rect 476580 388612 476632 388618
rect 476580 388554 476632 388560
rect 476592 385900 476620 388554
rect 477328 385900 477356 388991
rect 478052 388816 478104 388822
rect 478052 388758 478104 388764
rect 478064 385900 478092 388758
rect 478788 388544 478840 388550
rect 478788 388486 478840 388492
rect 478800 385900 478828 388486
rect 479536 385900 479564 388991
rect 480996 388884 481048 388890
rect 480996 388826 481048 388832
rect 480260 388748 480312 388754
rect 480260 388690 480312 388696
rect 480272 385900 480300 388690
rect 481008 385900 481036 388826
rect 481732 388680 481784 388686
rect 481732 388622 481784 388628
rect 481744 385900 481772 388622
rect 482468 388476 482520 388482
rect 482468 388418 482520 388424
rect 482480 385900 482508 388418
rect 483032 385914 483060 421534
rect 483676 398138 483704 429150
rect 485780 423360 485832 423366
rect 485780 423302 485832 423308
rect 483664 398132 483716 398138
rect 483664 398074 483716 398080
rect 483940 389020 483992 389026
rect 483940 388962 483992 388968
rect 483032 385886 483230 385914
rect 483952 385900 483980 388962
rect 484676 388748 484728 388754
rect 484676 388690 484728 388696
rect 484688 385900 484716 388690
rect 485412 388680 485464 388686
rect 485412 388622 485464 388628
rect 485424 385900 485452 388622
rect 485792 385914 485820 423302
rect 486436 389842 486464 429150
rect 487160 423292 487212 423298
rect 487160 423234 487212 423240
rect 486424 389836 486476 389842
rect 486424 389778 486476 389784
rect 486884 388612 486936 388618
rect 486884 388554 486936 388560
rect 485792 385886 486174 385914
rect 486896 385900 486924 388554
rect 487172 385914 487200 423234
rect 488540 423224 488592 423230
rect 488540 423166 488592 423172
rect 488552 402974 488580 423166
rect 488552 402946 488672 402974
rect 488356 388544 488408 388550
rect 488356 388486 488408 388492
rect 487172 385886 487646 385914
rect 488368 385900 488396 388486
rect 488644 385914 488672 402946
rect 490024 393990 490052 432126
rect 490012 393984 490064 393990
rect 490012 393926 490064 393932
rect 490564 389836 490616 389842
rect 490564 389778 490616 389784
rect 489828 388476 489880 388482
rect 489828 388418 489880 388424
rect 488644 385886 489118 385914
rect 489840 385900 489868 388418
rect 490576 385900 490604 389778
rect 491128 387122 491156 500126
rect 491312 500126 491372 500154
rect 491312 497486 491340 500126
rect 494072 499526 494100 507826
rect 494242 505200 494298 505209
rect 494242 505135 494244 505144
rect 494296 505135 494298 505144
rect 494244 505106 494296 505112
rect 494060 499520 494112 499526
rect 494060 499462 494112 499468
rect 494256 499458 494284 505106
rect 494702 501256 494758 501265
rect 494702 501191 494758 501200
rect 494244 499452 494296 499458
rect 494244 499394 494296 499400
rect 491300 497480 491352 497486
rect 491300 497422 491352 497428
rect 494716 462534 494744 501191
rect 494704 462528 494756 462534
rect 494704 462470 494756 462476
rect 494716 456074 494744 462470
rect 494704 456068 494756 456074
rect 494704 456010 494756 456016
rect 502524 424380 502576 424386
rect 502524 424322 502576 424328
rect 496820 423156 496872 423162
rect 496820 423098 496872 423104
rect 494060 420232 494112 420238
rect 494060 420174 494112 420180
rect 492680 398132 492732 398138
rect 492680 398074 492732 398080
rect 491576 395344 491628 395350
rect 491576 395286 491628 395292
rect 491300 393984 491352 393990
rect 491300 393926 491352 393932
rect 491116 387116 491168 387122
rect 491116 387058 491168 387064
rect 491312 385900 491340 393926
rect 491588 385914 491616 395286
rect 492692 389298 492720 398074
rect 492772 396772 492824 396778
rect 492772 396714 492824 396720
rect 492680 389292 492732 389298
rect 492680 389234 492732 389240
rect 491588 385886 492062 385914
rect 492784 385900 492812 396714
rect 494072 389298 494100 420174
rect 494152 399492 494204 399498
rect 494152 399434 494204 399440
rect 493140 389292 493192 389298
rect 493140 389234 493192 389240
rect 494060 389292 494112 389298
rect 494060 389234 494112 389240
rect 493152 385914 493180 389234
rect 494164 385914 494192 399434
rect 496452 392692 496504 392698
rect 496452 392634 496504 392640
rect 495716 391332 495768 391338
rect 495716 391274 495768 391280
rect 494612 389292 494664 389298
rect 494612 389234 494664 389240
rect 494624 385914 494652 389234
rect 493152 385886 493534 385914
rect 494164 385886 494270 385914
rect 494624 385886 495006 385914
rect 495728 385900 495756 391274
rect 496464 385900 496492 392634
rect 496832 385914 496860 423098
rect 498200 423088 498252 423094
rect 498200 423030 498252 423036
rect 497464 400920 497516 400926
rect 497464 400862 497516 400868
rect 497476 385914 497504 400862
rect 498212 385914 498240 423030
rect 499580 423020 499632 423026
rect 499580 422962 499632 422968
rect 499592 402974 499620 422962
rect 501052 422952 501104 422958
rect 501052 422894 501104 422900
rect 501064 402974 501092 422894
rect 502536 402974 502564 424322
rect 502984 423428 503036 423434
rect 502984 423370 503036 423376
rect 499592 402946 499712 402974
rect 501064 402946 501184 402974
rect 502536 402946 502656 402974
rect 499396 388952 499448 388958
rect 499396 388894 499448 388900
rect 496832 385886 497214 385914
rect 497476 385886 497950 385914
rect 498212 385886 498686 385914
rect 499408 385900 499436 388894
rect 499684 385914 499712 402946
rect 500868 388884 500920 388890
rect 500868 388826 500920 388832
rect 499684 385886 500158 385914
rect 500880 385900 500908 388826
rect 501156 385914 501184 402946
rect 502340 388816 502392 388822
rect 502340 388758 502392 388764
rect 501156 385886 501630 385914
rect 502352 385900 502380 388758
rect 502628 385914 502656 402946
rect 502996 389026 503024 423370
rect 503720 417784 503772 417790
rect 503720 417726 503772 417732
rect 502984 389020 503036 389026
rect 502984 388962 503036 388968
rect 503732 385914 503760 417726
rect 507860 417716 507912 417722
rect 507860 417658 507912 417664
rect 506480 417648 506532 417654
rect 506480 417590 506532 417596
rect 503996 417512 504048 417518
rect 503996 417454 504048 417460
rect 504008 402974 504036 417454
rect 504008 402946 504128 402974
rect 504100 385914 504128 402946
rect 506020 392624 506072 392630
rect 506020 392566 506072 392572
rect 505284 391264 505336 391270
rect 505284 391206 505336 391212
rect 502628 385886 503102 385914
rect 503732 385886 503838 385914
rect 504100 385886 504574 385914
rect 505296 385900 505324 391206
rect 506032 385900 506060 392566
rect 506492 385914 506520 417590
rect 506572 417580 506624 417586
rect 506572 417522 506624 417528
rect 506584 402974 506612 417522
rect 506584 402946 507072 402974
rect 507044 385914 507072 402946
rect 507872 385914 507900 417658
rect 507952 417444 508004 417450
rect 507952 417386 508004 417392
rect 507964 402974 507992 417386
rect 507964 402946 508544 402974
rect 508516 385914 508544 402946
rect 506492 385886 506782 385914
rect 507044 385886 507518 385914
rect 507872 385886 508254 385914
rect 508516 385886 508990 385914
rect 453304 385416 453356 385422
rect 453304 385358 453356 385364
rect 509514 375592 509570 375601
rect 509514 375527 509570 375536
rect 509330 370152 509386 370161
rect 509330 370087 509386 370096
rect 450634 349072 450690 349081
rect 450634 349007 450690 349016
rect 450728 334688 450780 334694
rect 450728 334630 450780 334636
rect 450636 334620 450688 334626
rect 450636 334562 450688 334568
rect 450544 321428 450596 321434
rect 450544 321370 450596 321376
rect 450648 321026 450676 334562
rect 450740 322114 450768 334630
rect 507492 322720 507544 322726
rect 507492 322662 507544 322668
rect 507400 322584 507452 322590
rect 507400 322526 507452 322532
rect 507308 322516 507360 322522
rect 507308 322458 507360 322464
rect 463516 322448 463568 322454
rect 507124 322448 507176 322454
rect 463568 322396 463634 322402
rect 463516 322390 463634 322396
rect 507124 322390 507176 322396
rect 463528 322374 463634 322390
rect 464896 322380 464948 322386
rect 464896 322322 464948 322328
rect 459652 322312 459704 322318
rect 459494 322260 459652 322266
rect 463516 322312 463568 322318
rect 459494 322254 459704 322260
rect 459494 322238 459692 322254
rect 463252 322250 463358 322266
rect 463516 322254 463568 322260
rect 463240 322244 463358 322250
rect 463292 322238 463358 322244
rect 463240 322186 463292 322192
rect 450728 322108 450780 322114
rect 450728 322050 450780 322056
rect 455708 322102 455906 322130
rect 456076 322102 456182 322130
rect 456352 322102 456458 322130
rect 456628 322102 456734 322130
rect 450636 321020 450688 321026
rect 450636 320962 450688 320968
rect 455512 319252 455564 319258
rect 455512 319194 455564 319200
rect 455420 318912 455472 318918
rect 455420 318854 455472 318860
rect 452108 318232 452160 318238
rect 452108 318174 452160 318180
rect 450728 316872 450780 316878
rect 450728 316814 450780 316820
rect 450636 316804 450688 316810
rect 450636 316746 450688 316752
rect 450544 316736 450596 316742
rect 450544 316678 450596 316684
rect 449992 249756 450044 249762
rect 449992 249698 450044 249704
rect 450004 248470 450032 249698
rect 449992 248464 450044 248470
rect 449992 248406 450044 248412
rect 450004 163130 450032 248406
rect 449992 163124 450044 163130
rect 449992 163066 450044 163072
rect 449900 62824 449952 62830
rect 449900 62766 449952 62772
rect 409234 44840 409290 44849
rect 409234 44775 409290 44784
rect 405004 3528 405056 3534
rect 405004 3470 405056 3476
rect 361120 3392 361172 3398
rect 361120 3334 361172 3340
rect 361028 3256 361080 3262
rect 361028 3198 361080 3204
rect 450556 2174 450584 316678
rect 450648 3466 450676 316746
rect 450740 3505 450768 316814
rect 452016 315376 452068 315382
rect 452016 315318 452068 315324
rect 451096 314288 451148 314294
rect 451096 314230 451148 314236
rect 451004 314220 451056 314226
rect 451004 314162 451056 314168
rect 450820 314016 450872 314022
rect 450820 313958 450872 313964
rect 450832 39370 450860 313958
rect 450912 313948 450964 313954
rect 450912 313890 450964 313896
rect 450924 46442 450952 313890
rect 450912 46436 450964 46442
rect 450912 46378 450964 46384
rect 451016 46238 451044 314162
rect 451108 46306 451136 314230
rect 451924 311228 451976 311234
rect 451924 311170 451976 311176
rect 451188 160200 451240 160206
rect 451188 160142 451240 160148
rect 451200 142866 451228 160142
rect 451740 158432 451792 158438
rect 451740 158374 451792 158380
rect 451752 158273 451780 158374
rect 451738 158264 451794 158273
rect 451738 158199 451794 158208
rect 451188 142860 451240 142866
rect 451188 142802 451240 142808
rect 451936 125633 451964 311170
rect 452028 148753 452056 315318
rect 452120 155553 452148 318174
rect 455236 318096 455288 318102
rect 455236 318038 455288 318044
rect 453580 317280 453632 317286
rect 453580 317222 453632 317228
rect 454958 317248 455014 317257
rect 453396 317144 453448 317150
rect 453396 317086 453448 317092
rect 453302 316976 453358 316985
rect 453302 316911 453358 316920
rect 452200 314084 452252 314090
rect 452200 314026 452252 314032
rect 452106 155544 452162 155553
rect 452106 155479 452162 155488
rect 452212 154193 452240 314026
rect 452476 283620 452528 283626
rect 452476 283562 452528 283568
rect 452292 275324 452344 275330
rect 452292 275266 452344 275272
rect 452198 154184 452254 154193
rect 452198 154119 452254 154128
rect 452108 152992 452160 152998
rect 452108 152934 452160 152940
rect 452120 152833 452148 152934
rect 452106 152824 452162 152833
rect 452106 152759 452162 152768
rect 452014 148744 452070 148753
rect 452014 148679 452070 148688
rect 452108 140684 452160 140690
rect 452108 140626 452160 140632
rect 452120 140593 452148 140626
rect 452106 140584 452162 140593
rect 452106 140519 452162 140528
rect 452108 132456 452160 132462
rect 452106 132424 452108 132433
rect 452160 132424 452162 132433
rect 452106 132359 452162 132368
rect 452304 128353 452332 275266
rect 452384 268456 452436 268462
rect 452384 268398 452436 268404
rect 452396 129713 452424 268398
rect 452488 150113 452516 283562
rect 453212 271176 453264 271182
rect 453212 271118 453264 271124
rect 452568 156936 452620 156942
rect 452566 156904 452568 156913
rect 452620 156904 452622 156913
rect 452566 156839 452622 156848
rect 452568 151496 452620 151502
rect 452566 151464 452568 151473
rect 452620 151464 452622 151473
rect 452566 151399 452622 151408
rect 452474 150104 452530 150113
rect 452474 150039 452530 150048
rect 452568 147416 452620 147422
rect 452566 147384 452568 147393
rect 452620 147384 452622 147393
rect 452566 147319 452622 147328
rect 452568 146192 452620 146198
rect 452568 146134 452620 146140
rect 452580 146033 452608 146134
rect 452566 146024 452622 146033
rect 452566 145959 452622 145968
rect 452568 144696 452620 144702
rect 452566 144664 452568 144673
rect 452620 144664 452622 144673
rect 452566 144599 452622 144608
rect 452568 143336 452620 143342
rect 452566 143304 452568 143313
rect 452620 143304 452622 143313
rect 452566 143239 452622 143248
rect 452568 141976 452620 141982
rect 452566 141944 452568 141953
rect 452620 141944 452622 141953
rect 452566 141879 452622 141888
rect 452568 139392 452620 139398
rect 452568 139334 452620 139340
rect 452580 139233 452608 139334
rect 452566 139224 452622 139233
rect 452566 139159 452622 139168
rect 452568 137896 452620 137902
rect 452566 137864 452568 137873
rect 452620 137864 452622 137873
rect 452566 137799 452622 137808
rect 452568 136536 452620 136542
rect 452566 136504 452568 136513
rect 452620 136504 452622 136513
rect 452566 136439 452622 136448
rect 452568 135176 452620 135182
rect 452566 135144 452568 135153
rect 452620 135144 452622 135153
rect 452566 135079 452622 135088
rect 452476 133816 452528 133822
rect 452474 133784 452476 133793
rect 452528 133784 452530 133793
rect 452474 133719 452530 133728
rect 452568 131096 452620 131102
rect 452566 131064 452568 131073
rect 452620 131064 452622 131073
rect 452566 130999 452622 131008
rect 452382 129704 452438 129713
rect 452382 129639 452438 129648
rect 452290 128344 452346 128353
rect 452290 128279 452346 128288
rect 452198 126984 452254 126993
rect 453224 126954 453252 271118
rect 452198 126919 452200 126928
rect 452252 126919 452254 126928
rect 453212 126948 453264 126954
rect 452200 126890 452252 126896
rect 453212 126890 453264 126896
rect 451922 125624 451978 125633
rect 451922 125559 451978 125568
rect 451740 124772 451792 124778
rect 451740 124714 451792 124720
rect 451752 124273 451780 124714
rect 451738 124264 451794 124273
rect 451738 124199 451794 124208
rect 451740 123140 451792 123146
rect 451740 123082 451792 123088
rect 451752 122913 451780 123082
rect 451738 122904 451794 122913
rect 451738 122839 451794 122848
rect 451740 121644 451792 121650
rect 451740 121586 451792 121592
rect 451752 121553 451780 121586
rect 451738 121544 451794 121553
rect 451738 121479 451794 121488
rect 451096 46300 451148 46306
rect 451096 46242 451148 46248
rect 451004 46232 451056 46238
rect 451004 46174 451056 46180
rect 450820 39364 450872 39370
rect 450820 39306 450872 39312
rect 450726 3496 450782 3505
rect 450636 3460 450688 3466
rect 450726 3431 450782 3440
rect 450636 3402 450688 3408
rect 450544 2168 450596 2174
rect 450544 2110 450596 2116
rect 453316 2106 453344 316911
rect 453408 45558 453436 317086
rect 453488 316600 453540 316606
rect 453488 316542 453540 316548
rect 453500 46510 453528 316542
rect 453592 46578 453620 317222
rect 454776 317212 454828 317218
rect 454958 317183 455014 317192
rect 454776 317154 454828 317160
rect 454682 316704 454738 316713
rect 454682 316639 454738 316648
rect 453672 309800 453724 309806
rect 453672 309742 453724 309748
rect 453684 132462 453712 309742
rect 453764 308508 453816 308514
rect 453764 308450 453816 308456
rect 453776 133822 453804 308450
rect 453856 285048 453908 285054
rect 453856 284990 453908 284996
rect 453764 133816 453816 133822
rect 453764 133758 453816 133764
rect 453672 132456 453724 132462
rect 453672 132398 453724 132404
rect 453868 124778 453896 284990
rect 453948 279472 454000 279478
rect 453948 279414 454000 279420
rect 453960 131102 453988 279414
rect 454040 207664 454092 207670
rect 454040 207606 454092 207612
rect 454052 164898 454080 207606
rect 454040 164892 454092 164898
rect 454040 164834 454092 164840
rect 453948 131096 454000 131102
rect 453948 131038 454000 131044
rect 453856 124772 453908 124778
rect 453856 124714 453908 124720
rect 453580 46572 453632 46578
rect 453580 46514 453632 46520
rect 453488 46504 453540 46510
rect 453488 46446 453540 46452
rect 453396 45552 453448 45558
rect 453396 45494 453448 45500
rect 454696 3369 454724 316639
rect 454788 136542 454816 317154
rect 454868 316940 454920 316946
rect 454868 316882 454920 316888
rect 454880 306202 454908 316882
rect 454972 306338 455000 317183
rect 455052 317076 455104 317082
rect 455052 317018 455104 317024
rect 454960 306332 455012 306338
rect 454960 306274 455012 306280
rect 455064 306270 455092 317018
rect 455052 306264 455104 306270
rect 455052 306206 455104 306212
rect 454868 306196 454920 306202
rect 454868 306138 454920 306144
rect 455052 282260 455104 282266
rect 455052 282202 455104 282208
rect 454868 276684 454920 276690
rect 454868 276626 454920 276632
rect 454776 136536 454828 136542
rect 454776 136478 454828 136484
rect 454880 123146 454908 276626
rect 454960 271244 455012 271250
rect 454960 271186 455012 271192
rect 454868 123140 454920 123146
rect 454868 123082 454920 123088
rect 454972 121650 455000 271186
rect 455064 144702 455092 282202
rect 455144 274032 455196 274038
rect 455144 273974 455196 273980
rect 455052 144696 455104 144702
rect 455052 144638 455104 144644
rect 455156 140690 455184 273974
rect 455248 222154 455276 318038
rect 455432 301510 455460 318854
rect 455524 303006 455552 319194
rect 455604 318980 455656 318986
rect 455604 318922 455656 318928
rect 455616 304434 455644 318922
rect 455708 315314 455736 322102
rect 456076 318986 456104 322102
rect 456156 319456 456208 319462
rect 456156 319398 456208 319404
rect 456064 318980 456116 318986
rect 456064 318922 456116 318928
rect 456064 318096 456116 318102
rect 456064 318038 456116 318044
rect 455696 315308 455748 315314
rect 455696 315250 455748 315256
rect 455604 304428 455656 304434
rect 455604 304370 455656 304376
rect 455512 303000 455564 303006
rect 455512 302942 455564 302948
rect 455420 301504 455472 301510
rect 455420 301446 455472 301452
rect 455236 222148 455288 222154
rect 455236 222090 455288 222096
rect 455144 140684 455196 140690
rect 455144 140626 455196 140632
rect 454960 121644 455012 121650
rect 454960 121586 455012 121592
rect 456076 3738 456104 318038
rect 456168 46617 456196 319398
rect 456352 319258 456380 322102
rect 456340 319252 456392 319258
rect 456340 319194 456392 319200
rect 456628 318918 456656 322102
rect 456892 318980 456944 318986
rect 456892 318922 456944 318928
rect 456616 318912 456668 318918
rect 456616 318854 456668 318860
rect 456340 317416 456392 317422
rect 456340 317358 456392 317364
rect 456248 317008 456300 317014
rect 456248 316950 456300 316956
rect 456154 46608 456210 46617
rect 456154 46543 456210 46552
rect 456260 44878 456288 316950
rect 456352 46714 456380 317358
rect 456524 317348 456576 317354
rect 456524 317290 456576 317296
rect 456432 316668 456484 316674
rect 456432 316610 456484 316616
rect 456340 46708 456392 46714
rect 456340 46650 456392 46656
rect 456444 46646 456472 316610
rect 456536 47054 456564 317290
rect 456904 296002 456932 318922
rect 456996 300762 457024 322116
rect 457180 322102 457286 322130
rect 457456 322102 457562 322130
rect 456984 300756 457036 300762
rect 456984 300698 457036 300704
rect 457180 298110 457208 322102
rect 457456 318986 457484 322102
rect 457444 318980 457496 318986
rect 457444 318922 457496 318928
rect 457824 318374 457852 322116
rect 458100 321230 458128 322116
rect 458088 321224 458140 321230
rect 458088 321166 458140 321172
rect 458376 321162 458404 322116
rect 458364 321156 458416 321162
rect 458364 321098 458416 321104
rect 458652 320142 458680 322116
rect 458928 321570 458956 322116
rect 459204 321774 459232 322116
rect 459192 321768 459244 321774
rect 459192 321710 459244 321716
rect 459756 321638 459784 322116
rect 459744 321632 459796 321638
rect 459744 321574 459796 321580
rect 458916 321564 458968 321570
rect 458916 321506 458968 321512
rect 460032 321473 460060 322116
rect 460202 322008 460258 322017
rect 460202 321943 460258 321952
rect 460018 321464 460074 321473
rect 460018 321399 460074 321408
rect 458640 320136 458692 320142
rect 458640 320078 458692 320084
rect 458916 319660 458968 319666
rect 458916 319602 458968 319608
rect 457812 318368 457864 318374
rect 457812 318310 457864 318316
rect 458824 318164 458876 318170
rect 458824 318106 458876 318112
rect 457444 314152 457496 314158
rect 457444 314094 457496 314100
rect 457168 298104 457220 298110
rect 457168 298046 457220 298052
rect 456892 295996 456944 296002
rect 456892 295938 456944 295944
rect 456616 273964 456668 273970
rect 456616 273906 456668 273912
rect 456628 156942 456656 273906
rect 456708 269952 456760 269958
rect 456708 269894 456760 269900
rect 456720 158438 456748 269894
rect 456800 263560 456852 263566
rect 456800 263502 456852 263508
rect 456812 262721 456840 263502
rect 456798 262712 456854 262721
rect 456798 262647 456854 262656
rect 456798 248840 456854 248849
rect 456798 248775 456854 248784
rect 456812 248470 456840 248775
rect 456800 248464 456852 248470
rect 456800 248406 456852 248412
rect 456800 222148 456852 222154
rect 456800 222090 456852 222096
rect 456812 221105 456840 222090
rect 456798 221096 456854 221105
rect 456798 221031 456854 221040
rect 456812 198014 456840 221031
rect 456892 207664 456944 207670
rect 456892 207606 456944 207612
rect 456904 207233 456932 207606
rect 456890 207224 456946 207233
rect 456890 207159 456946 207168
rect 456800 198008 456852 198014
rect 456800 197950 456852 197956
rect 456812 162178 456840 197950
rect 456800 162172 456852 162178
rect 456800 162114 456852 162120
rect 456708 158432 456760 158438
rect 456708 158374 456760 158380
rect 456616 156936 456668 156942
rect 456616 156878 456668 156884
rect 456524 47048 456576 47054
rect 456524 46990 456576 46996
rect 456432 46640 456484 46646
rect 456432 46582 456484 46588
rect 457456 46374 457484 314094
rect 457536 306196 457588 306202
rect 457536 306138 457588 306144
rect 457548 146198 457576 306138
rect 457628 280832 457680 280838
rect 457628 280774 457680 280780
rect 457536 146192 457588 146198
rect 457536 146134 457588 146140
rect 457640 141982 457668 280774
rect 457720 272604 457772 272610
rect 457720 272546 457772 272552
rect 457628 141976 457680 141982
rect 457628 141918 457680 141924
rect 457732 137902 457760 272546
rect 457812 272536 457864 272542
rect 457812 272478 457864 272484
rect 457824 151502 457852 272478
rect 457904 265668 457956 265674
rect 457904 265610 457956 265616
rect 457916 248414 457944 265610
rect 457916 248386 458128 248414
rect 458100 234977 458128 248386
rect 458086 234968 458142 234977
rect 458086 234903 458142 234912
rect 458100 162246 458128 234903
rect 458730 207224 458786 207233
rect 458730 207159 458786 207168
rect 458744 200802 458772 207159
rect 458732 200796 458784 200802
rect 458732 200738 458784 200744
rect 458088 162240 458140 162246
rect 458088 162182 458140 162188
rect 457812 151496 457864 151502
rect 457812 151438 457864 151444
rect 457720 137896 457772 137902
rect 457720 137838 457772 137844
rect 457444 46368 457496 46374
rect 457444 46310 457496 46316
rect 456248 44872 456300 44878
rect 456248 44814 456300 44820
rect 458836 4010 458864 318106
rect 458928 46889 458956 319602
rect 459100 319592 459152 319598
rect 459100 319534 459152 319540
rect 459008 316532 459060 316538
rect 459008 316474 459060 316480
rect 458914 46880 458970 46889
rect 458914 46815 458970 46824
rect 459020 46782 459048 316474
rect 459008 46776 459060 46782
rect 459112 46753 459140 319534
rect 459192 318300 459244 318306
rect 459192 318242 459244 318248
rect 459204 135182 459232 318242
rect 459284 279540 459336 279546
rect 459284 279482 459336 279488
rect 459296 139398 459324 279482
rect 459468 275392 459520 275398
rect 459468 275334 459520 275340
rect 459376 271312 459428 271318
rect 459376 271254 459428 271260
rect 459388 143342 459416 271254
rect 459480 147422 459508 275334
rect 459468 147416 459520 147422
rect 459468 147358 459520 147364
rect 459376 143336 459428 143342
rect 459376 143278 459428 143284
rect 459284 139392 459336 139398
rect 459284 139334 459336 139340
rect 459192 135176 459244 135182
rect 459192 135118 459244 135124
rect 459008 46718 459060 46724
rect 459098 46744 459154 46753
rect 459098 46679 459154 46688
rect 460216 39778 460244 321943
rect 460308 320006 460336 322116
rect 460584 321706 460612 322116
rect 460572 321700 460624 321706
rect 460572 321642 460624 321648
rect 460860 321502 460888 322116
rect 460848 321496 460900 321502
rect 460848 321438 460900 321444
rect 461136 320074 461164 322116
rect 461412 321434 461440 322116
rect 461400 321428 461452 321434
rect 461400 321370 461452 321376
rect 461688 321201 461716 322116
rect 461674 321192 461730 321201
rect 461674 321127 461730 321136
rect 461860 320884 461912 320890
rect 461860 320826 461912 320832
rect 461872 320142 461900 320826
rect 461964 320618 461992 322116
rect 462240 321881 462268 322116
rect 462226 321872 462282 321881
rect 462226 321807 462282 321816
rect 462516 321366 462544 322116
rect 462504 321360 462556 321366
rect 462504 321302 462556 321308
rect 461952 320612 462004 320618
rect 461952 320554 462004 320560
rect 461860 320136 461912 320142
rect 461860 320078 461912 320084
rect 461124 320068 461176 320074
rect 461124 320010 461176 320016
rect 460296 320000 460348 320006
rect 460296 319942 460348 319948
rect 462792 319734 462820 322116
rect 463068 319802 463096 322116
rect 463528 321638 463556 322254
rect 463896 321842 463924 322116
rect 464080 322102 464186 322130
rect 464356 322102 464462 322130
rect 463884 321836 463936 321842
rect 463884 321778 463936 321784
rect 463516 321632 463568 321638
rect 463516 321574 463568 321580
rect 463056 319796 463108 319802
rect 463056 319738 463108 319744
rect 462780 319728 462832 319734
rect 462780 319670 462832 319676
rect 460388 319524 460440 319530
rect 460388 319466 460440 319472
rect 460296 319388 460348 319394
rect 460296 319330 460348 319336
rect 460308 46918 460336 319330
rect 460296 46912 460348 46918
rect 460296 46854 460348 46860
rect 460400 46850 460428 319466
rect 464080 319138 464108 322102
rect 463804 319110 464108 319138
rect 461584 318368 461636 318374
rect 461584 318310 461636 318316
rect 461596 299470 461624 318310
rect 463804 310962 463832 319110
rect 464356 316034 464384 322102
rect 464080 316006 464384 316034
rect 461676 310956 461728 310962
rect 461676 310898 461728 310904
rect 463792 310956 463844 310962
rect 463792 310898 463844 310904
rect 461688 304502 461716 310898
rect 464080 305590 464108 316006
rect 464724 314294 464752 322116
rect 464908 320142 464936 322322
rect 502156 322244 502208 322250
rect 502156 322186 502208 322192
rect 471796 322176 471848 322182
rect 464896 320136 464948 320142
rect 464896 320078 464948 320084
rect 465000 316606 465028 322116
rect 464988 316600 465040 316606
rect 464988 316542 465040 316548
rect 465276 316538 465304 322116
rect 465552 319666 465580 322116
rect 465540 319660 465592 319666
rect 465540 319602 465592 319608
rect 465828 319394 465856 322116
rect 466012 322102 466118 322130
rect 466288 322102 466394 322130
rect 465816 319388 465868 319394
rect 465816 319330 465868 319336
rect 466012 319138 466040 322102
rect 465460 319110 466040 319138
rect 465264 316532 465316 316538
rect 465264 316474 465316 316480
rect 464712 314288 464764 314294
rect 464712 314230 464764 314236
rect 465460 306134 465488 319110
rect 466288 316034 466316 322102
rect 466552 319252 466604 319258
rect 466552 319194 466604 319200
rect 465736 316006 466316 316034
rect 465736 307086 465764 316006
rect 465724 307080 465776 307086
rect 465724 307022 465776 307028
rect 465448 306128 465500 306134
rect 465448 306070 465500 306076
rect 464068 305584 464120 305590
rect 464068 305526 464120 305532
rect 461676 304496 461728 304502
rect 461676 304438 461728 304444
rect 461584 299464 461636 299470
rect 461584 299406 461636 299412
rect 465724 288448 465776 288454
rect 465724 288390 465776 288396
rect 460480 278044 460532 278050
rect 460480 277986 460532 277992
rect 460492 152998 460520 277986
rect 465736 274106 465764 288390
rect 460572 274100 460624 274106
rect 460572 274042 460624 274048
rect 465724 274100 465776 274106
rect 465724 274042 465776 274048
rect 460584 267034 460612 274042
rect 466564 268394 466592 319194
rect 466656 312594 466684 322116
rect 466828 318980 466880 318986
rect 466828 318922 466880 318928
rect 466644 312588 466696 312594
rect 466644 312530 466696 312536
rect 466840 282198 466868 318922
rect 466932 291718 466960 322116
rect 467116 322102 467222 322130
rect 467392 322102 467498 322130
rect 467668 322102 467774 322130
rect 467944 322102 468050 322130
rect 468220 322102 468326 322130
rect 471848 322124 471914 322130
rect 471796 322118 471914 322124
rect 467116 318986 467144 322102
rect 467392 319258 467420 322102
rect 467380 319252 467432 319258
rect 467380 319194 467432 319200
rect 467104 318980 467156 318986
rect 467104 318922 467156 318928
rect 467668 316034 467696 322102
rect 467116 316006 467696 316034
rect 467116 293282 467144 316006
rect 467104 293276 467156 293282
rect 467104 293218 467156 293224
rect 466920 291712 466972 291718
rect 466920 291654 466972 291660
rect 466828 282192 466880 282198
rect 466828 282134 466880 282140
rect 467944 269890 467972 322102
rect 468220 313274 468248 322102
rect 468588 321366 468616 322116
rect 468576 321360 468628 321366
rect 468576 321302 468628 321308
rect 468864 319258 468892 322116
rect 469140 321842 469168 322116
rect 469128 321836 469180 321842
rect 469128 321778 469180 321784
rect 469416 319666 469444 322116
rect 469692 320074 469720 322116
rect 469968 321434 469996 322116
rect 470244 321502 470272 322116
rect 470232 321496 470284 321502
rect 470232 321438 470284 321444
rect 469956 321428 470008 321434
rect 469956 321370 470008 321376
rect 469680 320068 469732 320074
rect 469680 320010 469732 320016
rect 470520 319938 470548 322116
rect 470508 319932 470560 319938
rect 470508 319874 470560 319880
rect 469404 319660 469456 319666
rect 469404 319602 469456 319608
rect 468852 319252 468904 319258
rect 468852 319194 468904 319200
rect 470796 318782 470824 322116
rect 471072 319870 471100 322116
rect 471348 321094 471376 322116
rect 471336 321088 471388 321094
rect 471336 321030 471388 321036
rect 471060 319864 471112 319870
rect 471624 319841 471652 322116
rect 471808 322102 471914 322118
rect 471060 319806 471112 319812
rect 471610 319832 471666 319841
rect 471610 319767 471666 319776
rect 472176 319569 472204 322116
rect 472452 320754 472480 322116
rect 472440 320748 472492 320754
rect 472440 320690 472492 320696
rect 472728 319705 472756 322116
rect 472714 319696 472770 319705
rect 472714 319631 472770 319640
rect 472162 319560 472218 319569
rect 472162 319495 472218 319504
rect 473004 319190 473032 322116
rect 473280 319326 473308 322116
rect 473556 320958 473584 322116
rect 473544 320952 473596 320958
rect 473544 320894 473596 320900
rect 473832 320686 473860 322116
rect 474108 321910 474136 322116
rect 474096 321904 474148 321910
rect 474096 321846 474148 321852
rect 473820 320680 473872 320686
rect 473820 320622 473872 320628
rect 474384 320142 474412 322116
rect 474568 322102 474674 322130
rect 474372 320136 474424 320142
rect 474372 320078 474424 320084
rect 473268 319320 473320 319326
rect 473268 319262 473320 319268
rect 472992 319184 473044 319190
rect 472992 319126 473044 319132
rect 470784 318776 470836 318782
rect 470784 318718 470836 318724
rect 474568 316034 474596 322102
rect 474832 319184 474884 319190
rect 474832 319126 474884 319132
rect 473740 316006 474596 316034
rect 468208 313268 468260 313274
rect 468208 313210 468260 313216
rect 473740 307766 473768 316006
rect 474844 313954 474872 319126
rect 474936 316034 474964 322116
rect 475120 322102 475226 322130
rect 475120 319190 475148 322102
rect 475108 319184 475160 319190
rect 475108 319126 475160 319132
rect 475488 316674 475516 322116
rect 475764 317422 475792 322116
rect 476040 319598 476068 322116
rect 476028 319592 476080 319598
rect 476028 319534 476080 319540
rect 476316 319530 476344 322116
rect 476592 321554 476620 322116
rect 476776 322102 476882 322130
rect 477052 322102 477158 322130
rect 477328 322102 477434 322130
rect 476592 321526 476712 321554
rect 476304 319524 476356 319530
rect 476304 319466 476356 319472
rect 476212 319184 476264 319190
rect 476212 319126 476264 319132
rect 475752 317416 475804 317422
rect 475752 317358 475804 317364
rect 475476 316668 475528 316674
rect 475476 316610 475528 316616
rect 474936 316006 475056 316034
rect 475028 314226 475056 316006
rect 475016 314220 475068 314226
rect 475016 314162 475068 314168
rect 474832 313948 474884 313954
rect 474832 313890 474884 313896
rect 471244 307760 471296 307766
rect 471244 307702 471296 307708
rect 473728 307760 473780 307766
rect 473728 307702 473780 307708
rect 471256 288454 471284 307702
rect 476224 294574 476252 319126
rect 476488 318980 476540 318986
rect 476488 318922 476540 318928
rect 476500 306134 476528 318922
rect 476684 316034 476712 321526
rect 476776 318986 476804 322102
rect 476764 318980 476816 318986
rect 476764 318922 476816 318928
rect 477052 316034 477080 322102
rect 477328 319190 477356 322102
rect 477316 319184 477368 319190
rect 477316 319126 477368 319132
rect 477592 319184 477644 319190
rect 477592 319126 477644 319132
rect 476592 316006 476712 316034
rect 476776 316006 477080 316034
rect 476488 306128 476540 306134
rect 476488 306070 476540 306076
rect 476212 294568 476264 294574
rect 476212 294510 476264 294516
rect 471244 288448 471296 288454
rect 471244 288390 471296 288396
rect 476592 284986 476620 316006
rect 476776 313954 476804 316006
rect 476764 313948 476816 313954
rect 476764 313890 476816 313896
rect 477604 289678 477632 319126
rect 477696 311166 477724 322116
rect 477880 322102 477986 322130
rect 478156 322102 478262 322130
rect 477684 311160 477736 311166
rect 477684 311102 477736 311108
rect 477880 290494 477908 322102
rect 478156 319190 478184 322102
rect 478144 319184 478196 319190
rect 478144 319126 478196 319132
rect 478524 318782 478552 322116
rect 478800 320006 478828 322116
rect 479076 321094 479104 322116
rect 479064 321088 479116 321094
rect 479064 321030 479116 321036
rect 479352 320142 479380 322116
rect 479628 321910 479656 322116
rect 479616 321904 479668 321910
rect 479616 321846 479668 321852
rect 479340 320136 479392 320142
rect 479340 320078 479392 320084
rect 478788 320000 478840 320006
rect 478788 319942 478840 319948
rect 479904 319734 479932 322116
rect 479892 319728 479944 319734
rect 479892 319670 479944 319676
rect 480180 319598 480208 322116
rect 480456 319802 480484 322116
rect 480732 321298 480760 322116
rect 480720 321292 480772 321298
rect 480720 321234 480772 321240
rect 481008 319870 481036 322116
rect 481192 322102 481298 322130
rect 481192 322046 481220 322102
rect 481180 322040 481232 322046
rect 481180 321982 481232 321988
rect 481560 320822 481588 322116
rect 481548 320816 481600 320822
rect 481548 320758 481600 320764
rect 481836 320550 481864 322116
rect 481824 320544 481876 320550
rect 481824 320486 481876 320492
rect 480996 319864 481048 319870
rect 480996 319806 481048 319812
rect 480444 319796 480496 319802
rect 480444 319738 480496 319744
rect 480168 319592 480220 319598
rect 480168 319534 480220 319540
rect 482112 319054 482140 322116
rect 482388 321337 482416 322116
rect 482374 321328 482430 321337
rect 482374 321263 482430 321272
rect 482664 319977 482692 322116
rect 482940 321745 482968 322116
rect 482926 321736 482982 321745
rect 482926 321671 482982 321680
rect 483216 320113 483244 322116
rect 483202 320104 483258 320113
rect 483202 320039 483258 320048
rect 482650 319968 482706 319977
rect 482650 319903 482706 319912
rect 483492 319122 483520 322116
rect 483768 321609 483796 322116
rect 483952 322102 484058 322130
rect 484228 322114 484334 322130
rect 484216 322108 484334 322114
rect 483952 321978 483980 322102
rect 484268 322102 484334 322108
rect 484216 322050 484268 322056
rect 483940 321972 483992 321978
rect 483940 321914 483992 321920
rect 483754 321600 483810 321609
rect 483754 321535 483810 321544
rect 484596 321026 484624 322116
rect 484780 322102 484886 322130
rect 485056 322102 485162 322130
rect 485332 322102 485438 322130
rect 484584 321020 484636 321026
rect 484584 320962 484636 320968
rect 484780 319138 484808 322102
rect 483480 319116 483532 319122
rect 483480 319058 483532 319064
rect 484504 319110 484808 319138
rect 482100 319048 482152 319054
rect 482100 318990 482152 318996
rect 478512 318776 478564 318782
rect 478512 318718 478564 318724
rect 479524 318776 479576 318782
rect 479524 318718 479576 318724
rect 477868 290488 477920 290494
rect 477868 290430 477920 290436
rect 477592 289672 477644 289678
rect 477592 289614 477644 289620
rect 476764 288448 476816 288454
rect 476764 288390 476816 288396
rect 476580 284980 476632 284986
rect 476580 284922 476632 284928
rect 467932 269884 467984 269890
rect 467932 269826 467984 269832
rect 476776 268598 476804 288390
rect 479536 273222 479564 318718
rect 484504 313342 484532 319110
rect 485056 316034 485084 322102
rect 484780 316006 485084 316034
rect 482284 313336 482336 313342
rect 482284 313278 482336 313284
rect 484492 313336 484544 313342
rect 484492 313278 484544 313284
rect 482296 288454 482324 313278
rect 482284 288448 482336 288454
rect 482284 288390 482336 288396
rect 479524 273216 479576 273222
rect 479524 273158 479576 273164
rect 484780 269346 484808 316006
rect 485332 314158 485360 322102
rect 485700 317286 485728 322116
rect 485872 319116 485924 319122
rect 485872 319058 485924 319064
rect 485688 317280 485740 317286
rect 485688 317222 485740 317228
rect 485320 314152 485372 314158
rect 485320 314094 485372 314100
rect 485884 302802 485912 319058
rect 485976 317150 486004 322116
rect 486252 317354 486280 322116
rect 486528 319462 486556 322116
rect 486712 322102 486818 322130
rect 486988 322102 487094 322130
rect 486516 319456 486568 319462
rect 486516 319398 486568 319404
rect 486240 317348 486292 317354
rect 486240 317290 486292 317296
rect 485964 317144 486016 317150
rect 485964 317086 486016 317092
rect 486712 316034 486740 322102
rect 486988 319122 487016 322102
rect 487252 319320 487304 319326
rect 487252 319262 487304 319268
rect 486976 319116 487028 319122
rect 486976 319058 487028 319064
rect 486160 316006 486740 316034
rect 485872 302796 485924 302802
rect 485872 302738 485924 302744
rect 486160 291650 486188 316006
rect 486148 291644 486200 291650
rect 486148 291586 486200 291592
rect 487264 287706 487292 319262
rect 487356 317150 487384 322116
rect 487540 322102 487646 322130
rect 487816 322102 487922 322130
rect 488092 322102 488198 322130
rect 488368 322102 488474 322130
rect 488644 322102 488750 322130
rect 487344 317144 487396 317150
rect 487344 317086 487396 317092
rect 487540 307222 487568 322102
rect 487816 319326 487844 322102
rect 487804 319320 487856 319326
rect 487804 319262 487856 319268
rect 488092 319138 488120 322102
rect 487816 319110 488120 319138
rect 487816 308446 487844 319110
rect 488368 316034 488396 322102
rect 488092 316006 488396 316034
rect 487804 308440 487856 308446
rect 487804 308382 487856 308388
rect 487528 307216 487580 307222
rect 487528 307158 487580 307164
rect 487252 287700 487304 287706
rect 487252 287642 487304 287648
rect 488092 269958 488120 316006
rect 488644 271250 488672 322102
rect 488908 319116 488960 319122
rect 488908 319058 488960 319064
rect 488632 271244 488684 271250
rect 488632 271186 488684 271192
rect 488920 271182 488948 319058
rect 489012 276690 489040 322116
rect 489196 322102 489302 322130
rect 489472 322102 489578 322130
rect 489748 322102 489854 322130
rect 490024 322102 490130 322130
rect 490300 322102 490406 322130
rect 490576 322102 490682 322130
rect 490852 322102 490958 322130
rect 491128 322102 491234 322130
rect 489196 285054 489224 322102
rect 489472 311234 489500 322102
rect 489748 319122 489776 322102
rect 489736 319116 489788 319122
rect 489736 319058 489788 319064
rect 489460 311228 489512 311234
rect 489460 311170 489512 311176
rect 489184 285048 489236 285054
rect 489184 284990 489236 284996
rect 489000 276684 489052 276690
rect 489000 276626 489052 276632
rect 490024 275330 490052 322102
rect 490012 275324 490064 275330
rect 490012 275266 490064 275272
rect 488908 271176 488960 271182
rect 488908 271118 488960 271124
rect 488080 269952 488132 269958
rect 488080 269894 488132 269900
rect 481088 269340 481140 269346
rect 481088 269282 481140 269288
rect 484768 269340 484820 269346
rect 484768 269282 484820 269288
rect 476764 268592 476816 268598
rect 476764 268534 476816 268540
rect 481100 268530 481128 269282
rect 481088 268524 481140 268530
rect 481088 268466 481140 268472
rect 490300 268462 490328 322102
rect 490576 279478 490604 322102
rect 490852 309806 490880 322102
rect 490840 309800 490892 309806
rect 490840 309742 490892 309748
rect 491128 308514 491156 322102
rect 491496 318306 491524 322116
rect 491680 322102 491786 322130
rect 491956 322102 492062 322130
rect 492232 322102 492338 322130
rect 492508 322102 492614 322130
rect 491680 319274 491708 322102
rect 491588 319246 491708 319274
rect 491484 318300 491536 318306
rect 491484 318242 491536 318248
rect 491588 317218 491616 319246
rect 491956 319104 491984 322102
rect 491680 319076 491984 319104
rect 491576 317212 491628 317218
rect 491576 317154 491628 317160
rect 491116 308508 491168 308514
rect 491116 308450 491168 308456
rect 490564 279472 490616 279478
rect 490564 279414 490616 279420
rect 491680 272610 491708 319076
rect 491944 318980 491996 318986
rect 491944 318922 491996 318928
rect 491956 274038 491984 318922
rect 492232 279546 492260 322102
rect 492508 318986 492536 322102
rect 492772 319048 492824 319054
rect 492772 318990 492824 318996
rect 492496 318980 492548 318986
rect 492496 318922 492548 318928
rect 492220 279540 492272 279546
rect 492220 279482 492272 279488
rect 492784 275398 492812 318990
rect 492876 280838 492904 322116
rect 493048 319116 493100 319122
rect 493048 319058 493100 319064
rect 493060 306202 493088 319058
rect 493048 306196 493100 306202
rect 493048 306138 493100 306144
rect 492864 280832 492916 280838
rect 492864 280774 492916 280780
rect 492772 275392 492824 275398
rect 492772 275334 492824 275340
rect 491944 274032 491996 274038
rect 491944 273974 491996 273980
rect 491668 272604 491720 272610
rect 491668 272546 491720 272552
rect 493152 271318 493180 322116
rect 493336 322102 493442 322130
rect 493612 322102 493718 322130
rect 493888 322102 493994 322130
rect 494164 322102 494270 322130
rect 493336 282266 493364 322102
rect 493612 319122 493640 322102
rect 493600 319116 493652 319122
rect 493600 319058 493652 319064
rect 493888 319054 493916 322102
rect 493876 319048 493928 319054
rect 493876 318990 493928 318996
rect 494164 315382 494192 322102
rect 494428 319320 494480 319326
rect 494428 319262 494480 319268
rect 494152 315376 494204 315382
rect 494152 315318 494204 315324
rect 493324 282260 493376 282266
rect 493324 282202 493376 282208
rect 494440 272542 494468 319262
rect 494532 283626 494560 322116
rect 494716 322102 494822 322130
rect 494992 322102 495098 322130
rect 495268 322102 495374 322130
rect 494716 319326 494744 322102
rect 494704 319320 494756 319326
rect 494704 319262 494756 319268
rect 494992 319104 495020 322102
rect 494716 319076 495020 319104
rect 494520 283620 494572 283626
rect 494520 283562 494572 283568
rect 494716 278050 494744 319076
rect 495268 316034 495296 322102
rect 495532 319048 495584 319054
rect 495532 318990 495584 318996
rect 494992 316006 495296 316034
rect 494992 314090 495020 316006
rect 494980 314084 495032 314090
rect 494980 314026 495032 314032
rect 495544 309874 495572 318990
rect 495636 318238 495664 322116
rect 495808 319116 495860 319122
rect 495808 319058 495860 319064
rect 495624 318232 495676 318238
rect 495624 318174 495676 318180
rect 495820 315353 495848 319058
rect 495806 315344 495862 315353
rect 495806 315279 495862 315288
rect 495532 309868 495584 309874
rect 495532 309810 495584 309816
rect 494704 278044 494756 278050
rect 494704 277986 494756 277992
rect 495912 273970 495940 322116
rect 496188 318238 496216 322116
rect 496372 322102 496478 322130
rect 496648 322102 496754 322130
rect 496372 319122 496400 322102
rect 496360 319116 496412 319122
rect 496360 319058 496412 319064
rect 496648 319054 496676 322102
rect 497016 321554 497044 322116
rect 497200 322102 497306 322130
rect 497476 322102 497582 322130
rect 497752 322102 497858 322130
rect 497016 321526 497136 321554
rect 496820 320952 496872 320958
rect 496820 320894 496872 320900
rect 496832 320142 496860 320894
rect 496820 320136 496872 320142
rect 496820 320078 496872 320084
rect 496912 319116 496964 319122
rect 496912 319058 496964 319064
rect 496636 319048 496688 319054
rect 496636 318990 496688 318996
rect 496176 318232 496228 318238
rect 496176 318174 496228 318180
rect 495900 273964 495952 273970
rect 495900 273906 495952 273912
rect 494428 272536 494480 272542
rect 494428 272478 494480 272484
rect 493140 271312 493192 271318
rect 493140 271254 493192 271260
rect 496924 268462 496952 319058
rect 497108 316034 497136 321526
rect 497200 319122 497228 322102
rect 497188 319116 497240 319122
rect 497188 319058 497240 319064
rect 497188 318980 497240 318986
rect 497188 318922 497240 318928
rect 497016 316006 497136 316034
rect 497016 309806 497044 316006
rect 497004 309800 497056 309806
rect 497004 309742 497056 309748
rect 497200 269958 497228 318922
rect 497476 273970 497504 322102
rect 497752 318986 497780 322102
rect 498120 319530 498148 322116
rect 498108 319524 498160 319530
rect 498108 319466 498160 319472
rect 498292 319048 498344 319054
rect 498292 318990 498344 318996
rect 497740 318980 497792 318986
rect 497740 318922 497792 318928
rect 497464 273964 497516 273970
rect 497464 273906 497516 273912
rect 498304 271250 498332 318990
rect 498396 284986 498424 322116
rect 498672 319394 498700 322116
rect 498856 322102 498962 322130
rect 499132 322102 499238 322130
rect 499408 322102 499514 322130
rect 498660 319388 498712 319394
rect 498660 319330 498712 319336
rect 498568 319116 498620 319122
rect 498568 319058 498620 319064
rect 498384 284980 498436 284986
rect 498384 284922 498436 284928
rect 498580 274038 498608 319058
rect 498856 275330 498884 322102
rect 499132 319054 499160 322102
rect 499408 319122 499436 322102
rect 499396 319116 499448 319122
rect 499396 319058 499448 319064
rect 499672 319116 499724 319122
rect 499672 319058 499724 319064
rect 499120 319048 499172 319054
rect 499120 318990 499172 318996
rect 498844 275324 498896 275330
rect 498844 275266 498896 275272
rect 498568 274032 498620 274038
rect 498568 273974 498620 273980
rect 498292 271244 498344 271250
rect 498292 271186 498344 271192
rect 499684 271182 499712 319058
rect 499776 276690 499804 322116
rect 499960 322102 500066 322130
rect 499960 278050 499988 322102
rect 500328 317286 500356 322116
rect 500512 322102 500618 322130
rect 500788 322102 500894 322130
rect 500316 317280 500368 317286
rect 500316 317222 500368 317228
rect 500512 316034 500540 322102
rect 500788 319122 500816 322102
rect 500776 319116 500828 319122
rect 500776 319058 500828 319064
rect 501052 319116 501104 319122
rect 501052 319058 501104 319064
rect 500236 316006 500540 316034
rect 500236 279478 500264 316006
rect 500224 279472 500276 279478
rect 500224 279414 500276 279420
rect 499948 278044 500000 278050
rect 499948 277986 500000 277992
rect 499764 276684 499816 276690
rect 499764 276626 499816 276632
rect 501064 272542 501092 319058
rect 501156 315382 501184 322116
rect 501340 322102 501446 322130
rect 501340 319122 501368 322102
rect 501328 319116 501380 319122
rect 501328 319058 501380 319064
rect 501708 318306 501736 322116
rect 501892 322102 501998 322130
rect 501696 318300 501748 318306
rect 501696 318242 501748 318248
rect 501892 316034 501920 322102
rect 502168 319666 502196 322186
rect 502156 319660 502208 319666
rect 502156 319602 502208 319608
rect 502260 319433 502288 322116
rect 502246 319424 502302 319433
rect 502246 319359 502302 319368
rect 502432 319116 502484 319122
rect 502432 319058 502484 319064
rect 501340 316006 501920 316034
rect 501144 315376 501196 315382
rect 501144 315318 501196 315324
rect 501340 314090 501368 316006
rect 501328 314084 501380 314090
rect 501328 314026 501380 314032
rect 502444 280838 502472 319058
rect 502536 317218 502564 322116
rect 502812 319462 502840 322116
rect 502996 322102 503102 322130
rect 503272 322102 503378 322130
rect 503548 322102 503654 322130
rect 503824 322102 503930 322130
rect 502800 319456 502852 319462
rect 502800 319398 502852 319404
rect 502996 319138 503024 322102
rect 502720 319110 503024 319138
rect 502524 317212 502576 317218
rect 502524 317154 502576 317160
rect 502720 311234 502748 319110
rect 503272 316034 503300 322102
rect 503548 319122 503576 322102
rect 503536 319116 503588 319122
rect 503536 319058 503588 319064
rect 502996 316006 503300 316034
rect 502996 314158 503024 316006
rect 502984 314152 503036 314158
rect 502984 314094 503036 314100
rect 502708 311228 502760 311234
rect 502708 311170 502760 311176
rect 502432 280832 502484 280838
rect 502432 280774 502484 280780
rect 501052 272536 501104 272542
rect 501052 272478 501104 272484
rect 499672 271176 499724 271182
rect 499672 271118 499724 271124
rect 503824 270026 503852 322102
rect 507136 289542 507164 322390
rect 507214 322280 507270 322289
rect 507214 322215 507270 322224
rect 507124 289536 507176 289542
rect 507124 289478 507176 289484
rect 507228 289406 507256 322215
rect 507320 289474 507348 322458
rect 507412 295322 507440 322526
rect 507400 295316 507452 295322
rect 507400 295258 507452 295264
rect 507504 295254 507532 322662
rect 507584 322652 507636 322658
rect 507584 322594 507636 322600
rect 507596 297294 507624 322594
rect 509344 303482 509372 370087
rect 509422 357640 509478 357649
rect 509422 357575 509478 357584
rect 509332 303476 509384 303482
rect 509332 303418 509384 303424
rect 509436 302870 509464 357575
rect 509528 322153 509556 375527
rect 510710 365664 510766 365673
rect 510710 365599 510766 365608
rect 509606 357640 509662 357649
rect 509606 357575 509662 357584
rect 509620 322658 509648 357575
rect 510724 354674 510752 365599
rect 510802 355872 510858 355881
rect 510802 355807 510858 355816
rect 510632 354646 510752 354674
rect 509790 348392 509846 348401
rect 509790 348327 509846 348336
rect 509698 344040 509754 344049
rect 509698 343975 509754 343984
rect 509712 323474 509740 343975
rect 509700 323468 509752 323474
rect 509700 323410 509752 323416
rect 509698 323368 509754 323377
rect 509698 323303 509754 323312
rect 509608 322652 509660 322658
rect 509608 322594 509660 322600
rect 509514 322144 509570 322153
rect 509514 322079 509570 322088
rect 509712 316878 509740 323303
rect 509804 322969 509832 348327
rect 509882 342408 509938 342417
rect 509882 342343 509938 342352
rect 509790 322960 509846 322969
rect 509790 322895 509846 322904
rect 509896 317082 509924 342343
rect 509974 334248 510030 334257
rect 509974 334183 510030 334192
rect 509988 322522 510016 334183
rect 510066 331936 510122 331945
rect 510066 331871 510122 331880
rect 510080 322726 510108 331871
rect 510158 330304 510214 330313
rect 510158 330239 510214 330248
rect 510068 322720 510120 322726
rect 510068 322662 510120 322668
rect 510172 322590 510200 330239
rect 510252 323468 510304 323474
rect 510252 323410 510304 323416
rect 510160 322584 510212 322590
rect 510160 322526 510212 322532
rect 509976 322516 510028 322522
rect 509976 322458 510028 322464
rect 509884 317076 509936 317082
rect 509884 317018 509936 317024
rect 510264 316946 510292 323410
rect 510252 316940 510304 316946
rect 510252 316882 510304 316888
rect 509700 316872 509752 316878
rect 509700 316814 509752 316820
rect 510632 303618 510660 354646
rect 510816 305930 510844 355807
rect 510894 354240 510950 354249
rect 510894 354175 510950 354184
rect 510908 305998 510936 354175
rect 510986 347712 511042 347721
rect 510986 347647 511042 347656
rect 511000 306066 511028 347647
rect 511078 346080 511134 346089
rect 511078 346015 511134 346024
rect 511092 317014 511120 346015
rect 511170 335744 511226 335753
rect 511170 335679 511226 335688
rect 511184 322454 511212 335679
rect 511172 322448 511224 322454
rect 511172 322390 511224 322396
rect 511276 319598 511304 590650
rect 512012 519586 512040 600086
rect 515404 599616 515456 599622
rect 515404 599558 515456 599564
rect 514024 536852 514076 536858
rect 514024 536794 514076 536800
rect 512000 519580 512052 519586
rect 512000 519522 512052 519528
rect 511448 423564 511500 423570
rect 511448 423506 511500 423512
rect 511356 404388 511408 404394
rect 511356 404330 511408 404336
rect 511368 321162 511396 404330
rect 511460 388754 511488 423506
rect 511448 388748 511500 388754
rect 511448 388690 511500 388696
rect 512184 386504 512236 386510
rect 512184 386446 512236 386452
rect 512000 386436 512052 386442
rect 512000 386378 512052 386384
rect 512012 380458 512040 386378
rect 512092 385076 512144 385082
rect 512092 385018 512144 385024
rect 512000 380452 512052 380458
rect 512000 380394 512052 380400
rect 511998 380352 512054 380361
rect 511998 380287 512000 380296
rect 512052 380287 512054 380296
rect 512000 380258 512052 380264
rect 512104 378978 512132 385018
rect 512012 378950 512132 378978
rect 512012 376553 512040 378950
rect 512196 378842 512224 386446
rect 512734 384704 512790 384713
rect 512734 384639 512790 384648
rect 512748 383790 512776 384639
rect 513286 384160 513342 384169
rect 513286 384095 513342 384104
rect 512736 383784 512788 383790
rect 512736 383726 512788 383732
rect 513300 383722 513328 384095
rect 513288 383716 513340 383722
rect 513288 383658 513340 383664
rect 513010 383616 513066 383625
rect 513010 383551 513066 383560
rect 512458 383072 512514 383081
rect 512458 383007 512460 383016
rect 512512 383007 512514 383016
rect 512460 382978 512512 382984
rect 512274 382528 512330 382537
rect 513024 382498 513052 383551
rect 512274 382463 512330 382472
rect 513012 382492 513064 382498
rect 512288 382362 512316 382463
rect 513012 382434 513064 382440
rect 512276 382356 512328 382362
rect 512276 382298 512328 382304
rect 512458 381984 512514 381993
rect 512458 381919 512514 381928
rect 512368 380452 512420 380458
rect 512368 380394 512420 380400
rect 512104 378814 512224 378842
rect 512104 377641 512132 378814
rect 512182 378720 512238 378729
rect 512182 378655 512238 378664
rect 512196 378350 512224 378655
rect 512184 378344 512236 378350
rect 512184 378286 512236 378292
rect 512274 378176 512330 378185
rect 512274 378111 512330 378120
rect 512090 377632 512146 377641
rect 512090 377567 512146 377576
rect 511998 376544 512054 376553
rect 511998 376479 512054 376488
rect 512090 372736 512146 372745
rect 512090 372671 512092 372680
rect 512144 372671 512146 372680
rect 512092 372642 512144 372648
rect 512090 371648 512146 371657
rect 512090 371583 512146 371592
rect 511998 367296 512054 367305
rect 511998 367231 512000 367240
rect 512052 367231 512054 367240
rect 512000 367202 512052 367208
rect 511998 364576 512054 364585
rect 511998 364511 512000 364520
rect 512052 364511 512054 364520
rect 512000 364482 512052 364488
rect 512104 364334 512132 371583
rect 512182 368384 512238 368393
rect 512182 368319 512238 368328
rect 512012 364306 512132 364334
rect 511538 354784 511594 354793
rect 511538 354719 511594 354728
rect 511448 352164 511500 352170
rect 511448 352106 511500 352112
rect 511460 321230 511488 352106
rect 511448 321224 511500 321230
rect 511448 321166 511500 321172
rect 511356 321156 511408 321162
rect 511356 321098 511408 321104
rect 511264 319592 511316 319598
rect 511264 319534 511316 319540
rect 511080 317008 511132 317014
rect 511080 316950 511132 316956
rect 510988 306060 511040 306066
rect 510988 306002 511040 306008
rect 510896 305992 510948 305998
rect 510896 305934 510948 305940
rect 510804 305924 510856 305930
rect 510804 305866 510856 305872
rect 510620 303612 510672 303618
rect 510620 303554 510672 303560
rect 509424 302864 509476 302870
rect 509424 302806 509476 302812
rect 511552 297362 511580 354719
rect 511906 325816 511962 325825
rect 511906 325751 511962 325760
rect 511920 322289 511948 325751
rect 511906 322280 511962 322289
rect 511906 322215 511962 322224
rect 512012 300150 512040 364306
rect 512090 364032 512146 364041
rect 512090 363967 512146 363976
rect 512104 363594 512132 363967
rect 512092 363588 512144 363594
rect 512092 363530 512144 363536
rect 512090 363488 512146 363497
rect 512090 363423 512146 363432
rect 512000 300144 512052 300150
rect 512000 300086 512052 300092
rect 512104 297430 512132 363423
rect 512196 304298 512224 368319
rect 512288 318170 512316 378111
rect 512380 374921 512408 380394
rect 512472 376038 512500 381919
rect 513286 381440 513342 381449
rect 513286 381375 513342 381384
rect 513300 380934 513328 381375
rect 513288 380928 513340 380934
rect 512826 380896 512882 380905
rect 513288 380870 513340 380876
rect 512826 380831 512882 380840
rect 512840 377466 512868 380831
rect 513286 379808 513342 379817
rect 513286 379743 513342 379752
rect 513300 379574 513328 379743
rect 513288 379568 513340 379574
rect 513288 379510 513340 379516
rect 513286 379264 513342 379273
rect 513286 379199 513342 379208
rect 513300 378282 513328 379199
rect 513288 378276 513340 378282
rect 513288 378218 513340 378224
rect 512828 377460 512880 377466
rect 512828 377402 512880 377408
rect 513194 377088 513250 377097
rect 513194 377023 513250 377032
rect 513208 376786 513236 377023
rect 513196 376780 513248 376786
rect 513196 376722 513248 376728
rect 512460 376032 512512 376038
rect 512460 375974 512512 375980
rect 513286 376000 513342 376009
rect 513286 375935 513342 375944
rect 513300 375698 513328 375935
rect 513288 375692 513340 375698
rect 513288 375634 513340 375640
rect 512366 374912 512422 374921
rect 512366 374847 512422 374856
rect 512458 374368 512514 374377
rect 512458 374303 512514 374312
rect 512472 374202 512500 374303
rect 512460 374196 512512 374202
rect 512460 374138 512512 374144
rect 512642 373824 512698 373833
rect 512642 373759 512644 373768
rect 512696 373759 512698 373768
rect 512644 373730 512696 373736
rect 513286 373280 513342 373289
rect 513286 373215 513342 373224
rect 513300 372774 513328 373215
rect 513288 372768 513340 372774
rect 513288 372710 513340 372716
rect 512458 372192 512514 372201
rect 512458 372127 512514 372136
rect 512472 371822 512500 372127
rect 512460 371816 512512 371822
rect 512460 371758 512512 371764
rect 513286 371104 513342 371113
rect 513286 371039 513342 371048
rect 513300 370122 513328 371039
rect 513288 370116 513340 370122
rect 513288 370058 513340 370064
rect 512734 370016 512790 370025
rect 512734 369951 512736 369960
rect 512788 369951 512790 369960
rect 512736 369922 512788 369928
rect 513286 369472 513342 369481
rect 513286 369407 513342 369416
rect 513300 368558 513328 369407
rect 513470 368928 513526 368937
rect 513470 368863 513526 368872
rect 513288 368552 513340 368558
rect 513288 368494 513340 368500
rect 512642 367840 512698 367849
rect 512642 367775 512698 367784
rect 512656 367402 512684 367775
rect 512644 367396 512696 367402
rect 512644 367338 512696 367344
rect 513194 366752 513250 366761
rect 513194 366687 513250 366696
rect 513208 365770 513236 366687
rect 513286 366208 513342 366217
rect 513286 366143 513342 366152
rect 513300 365906 513328 366143
rect 513288 365900 513340 365906
rect 513288 365842 513340 365848
rect 513196 365764 513248 365770
rect 513196 365706 513248 365712
rect 513286 365120 513342 365129
rect 513286 365055 513342 365064
rect 513300 364410 513328 365055
rect 513288 364404 513340 364410
rect 513288 364346 513340 364352
rect 513194 362944 513250 362953
rect 513194 362879 513250 362888
rect 512366 362400 512422 362409
rect 512366 362335 512368 362344
rect 512420 362335 512422 362344
rect 512368 362306 512420 362312
rect 513208 361826 513236 362879
rect 513286 361856 513342 361865
rect 513196 361820 513248 361826
rect 513286 361791 513342 361800
rect 513196 361762 513248 361768
rect 513300 361622 513328 361791
rect 513288 361616 513340 361622
rect 513288 361558 513340 361564
rect 512826 361312 512882 361321
rect 512826 361247 512882 361256
rect 512366 360768 512422 360777
rect 512366 360703 512422 360712
rect 512380 360330 512408 360703
rect 512840 360466 512868 361247
rect 512828 360460 512880 360466
rect 512828 360402 512880 360408
rect 513288 360392 513340 360398
rect 513288 360334 513340 360340
rect 512368 360324 512420 360330
rect 512368 360266 512420 360272
rect 513300 360233 513328 360334
rect 513286 360224 513342 360233
rect 513286 360159 513342 360168
rect 512918 359680 512974 359689
rect 512918 359615 512974 359624
rect 512366 359136 512422 359145
rect 512366 359071 512422 359080
rect 512380 358970 512408 359071
rect 512368 358964 512420 358970
rect 512368 358906 512420 358912
rect 512932 358902 512960 359615
rect 512920 358896 512972 358902
rect 512920 358838 512972 358844
rect 512458 358592 512514 358601
rect 512458 358527 512514 358536
rect 512366 353696 512422 353705
rect 512366 353631 512368 353640
rect 512420 353631 512422 353640
rect 512368 353602 512420 353608
rect 512366 352608 512422 352617
rect 512366 352543 512422 352552
rect 512380 352442 512408 352543
rect 512368 352436 512420 352442
rect 512368 352378 512420 352384
rect 512366 350976 512422 350985
rect 512366 350911 512368 350920
rect 512420 350911 512422 350920
rect 512368 350882 512420 350888
rect 512366 349344 512422 349353
rect 512366 349279 512368 349288
rect 512420 349279 512422 349288
rect 512368 349250 512420 349256
rect 512366 345536 512422 345545
rect 512366 345471 512422 345480
rect 512276 318164 512328 318170
rect 512276 318106 512328 318112
rect 512380 316810 512408 345471
rect 512472 318102 512500 358527
rect 512918 356416 512974 356425
rect 512918 356351 512974 356360
rect 512932 356250 512960 356351
rect 512920 356244 512972 356250
rect 512920 356186 512972 356192
rect 513286 355328 513342 355337
rect 513286 355263 513342 355272
rect 513300 355162 513328 355263
rect 513288 355156 513340 355162
rect 513288 355098 513340 355104
rect 512826 353152 512882 353161
rect 512826 353087 512828 353096
rect 512880 353087 512882 353096
rect 512828 353058 512880 353064
rect 513286 352064 513342 352073
rect 513286 351999 513288 352008
rect 513340 351999 513342 352008
rect 513288 351970 513340 351976
rect 513010 351520 513066 351529
rect 513010 351455 513066 351464
rect 513024 350674 513052 351455
rect 513012 350668 513064 350674
rect 513012 350610 513064 350616
rect 513194 350432 513250 350441
rect 513194 350367 513250 350376
rect 513010 349888 513066 349897
rect 513010 349823 513066 349832
rect 513024 349246 513052 349823
rect 513208 349586 513236 350367
rect 513196 349580 513248 349586
rect 513196 349522 513248 349528
rect 513012 349240 513064 349246
rect 513012 349182 513064 349188
rect 513010 348256 513066 348265
rect 513010 348191 513066 348200
rect 513024 348090 513052 348191
rect 513012 348084 513064 348090
rect 513012 348026 513064 348032
rect 513286 347168 513342 347177
rect 513286 347103 513342 347112
rect 513300 346730 513328 347103
rect 513288 346724 513340 346730
rect 513288 346666 513340 346672
rect 513102 346624 513158 346633
rect 513102 346559 513104 346568
rect 513156 346559 513158 346568
rect 513104 346530 513156 346536
rect 512550 344992 512606 345001
rect 512550 344927 512606 344936
rect 512460 318096 512512 318102
rect 512460 318038 512512 318044
rect 512368 316804 512420 316810
rect 512368 316746 512420 316752
rect 512564 305658 512592 344927
rect 512642 343904 512698 343913
rect 512642 343839 512698 343848
rect 512656 343738 512684 343839
rect 512644 343732 512696 343738
rect 512644 343674 512696 343680
rect 513010 343360 513066 343369
rect 513010 343295 513066 343304
rect 513024 343194 513052 343295
rect 513012 343188 513064 343194
rect 513012 343130 513064 343136
rect 513288 342304 513340 342310
rect 513286 342272 513288 342281
rect 513340 342272 513342 342281
rect 513286 342207 513342 342216
rect 513010 341728 513066 341737
rect 513010 341663 513066 341672
rect 513024 341154 513052 341663
rect 513286 341184 513342 341193
rect 513012 341148 513064 341154
rect 513286 341119 513342 341128
rect 513012 341090 513064 341096
rect 513300 341018 513328 341119
rect 513288 341012 513340 341018
rect 513288 340954 513340 340960
rect 513194 340640 513250 340649
rect 513194 340575 513250 340584
rect 513104 339584 513156 339590
rect 513102 339552 513104 339561
rect 513156 339552 513158 339561
rect 513208 339522 513236 340575
rect 513286 340096 513342 340105
rect 513286 340031 513342 340040
rect 513300 339658 513328 340031
rect 513288 339652 513340 339658
rect 513288 339594 513340 339600
rect 513102 339487 513158 339496
rect 513196 339516 513248 339522
rect 513196 339458 513248 339464
rect 512826 339008 512882 339017
rect 512826 338943 512882 338952
rect 512642 338464 512698 338473
rect 512642 338399 512698 338408
rect 512656 338298 512684 338399
rect 512644 338292 512696 338298
rect 512644 338234 512696 338240
rect 512840 338162 512868 338943
rect 512828 338156 512880 338162
rect 512828 338098 512880 338104
rect 513286 337920 513342 337929
rect 513286 337855 513342 337864
rect 512642 337376 512698 337385
rect 512642 337311 512698 337320
rect 512552 305652 512604 305658
rect 512552 305594 512604 305600
rect 512184 304292 512236 304298
rect 512184 304234 512236 304240
rect 512656 302938 512684 337311
rect 513300 337074 513328 337855
rect 513288 337068 513340 337074
rect 513288 337010 513340 337016
rect 513288 336932 513340 336938
rect 513288 336874 513340 336880
rect 513300 336841 513328 336874
rect 513286 336832 513342 336841
rect 513286 336767 513342 336776
rect 513286 336288 513342 336297
rect 513342 336246 513420 336274
rect 513286 336223 513342 336232
rect 512734 334656 512790 334665
rect 512734 334591 512790 334600
rect 512748 334354 512776 334591
rect 512736 334348 512788 334354
rect 512736 334290 512788 334296
rect 512918 332480 512974 332489
rect 512918 332415 512974 332424
rect 512932 331498 512960 332415
rect 512920 331492 512972 331498
rect 512920 331434 512972 331440
rect 512734 329216 512790 329225
rect 512734 329151 512790 329160
rect 512644 302932 512696 302938
rect 512644 302874 512696 302880
rect 512092 297424 512144 297430
rect 512092 297366 512144 297372
rect 511540 297356 511592 297362
rect 511540 297298 511592 297304
rect 507584 297288 507636 297294
rect 507584 297230 507636 297236
rect 507492 295248 507544 295254
rect 507492 295190 507544 295196
rect 507308 289468 507360 289474
rect 507308 289410 507360 289416
rect 507216 289400 507268 289406
rect 507216 289342 507268 289348
rect 503812 270020 503864 270026
rect 503812 269962 503864 269968
rect 497188 269952 497240 269958
rect 497188 269894 497240 269900
rect 512748 269822 512776 329151
rect 512826 325408 512882 325417
rect 512826 325343 512882 325352
rect 512840 304366 512868 325343
rect 513392 314022 513420 336246
rect 513380 314016 513432 314022
rect 513380 313958 513432 313964
rect 512828 304360 512880 304366
rect 512828 304302 512880 304308
rect 513484 303142 513512 368863
rect 513656 363588 513708 363594
rect 513656 363530 513708 363536
rect 513562 356960 513618 356969
rect 513562 356895 513618 356904
rect 513472 303136 513524 303142
rect 513472 303078 513524 303084
rect 513576 292534 513604 356895
rect 513668 303414 513696 363530
rect 513748 362364 513800 362370
rect 513748 362306 513800 362312
rect 513656 303408 513708 303414
rect 513656 303350 513708 303356
rect 513760 303346 513788 362306
rect 513840 358964 513892 358970
rect 513840 358906 513892 358912
rect 513852 303550 513880 358906
rect 513932 349308 513984 349314
rect 513932 349250 513984 349256
rect 513944 305862 513972 349250
rect 514036 319734 514064 536794
rect 514116 464432 514168 464438
rect 514116 464374 514168 464380
rect 514128 319938 514156 464374
rect 514208 380316 514260 380322
rect 514208 380258 514260 380264
rect 514220 358834 514248 380258
rect 514852 372700 514904 372706
rect 514852 372642 514904 372648
rect 514300 364540 514352 364546
rect 514300 364482 514352 364488
rect 514208 358828 514260 358834
rect 514208 358770 514260 358776
rect 514116 319932 514168 319938
rect 514116 319874 514168 319880
rect 514024 319728 514076 319734
rect 514024 319670 514076 319676
rect 513932 305856 513984 305862
rect 513932 305798 513984 305804
rect 513840 303544 513892 303550
rect 513840 303486 513892 303492
rect 513748 303340 513800 303346
rect 513748 303282 513800 303288
rect 514312 297974 514340 364482
rect 514760 334348 514812 334354
rect 514760 334290 514812 334296
rect 514772 316742 514800 334290
rect 514760 316736 514812 316742
rect 514760 316678 514812 316684
rect 514300 297968 514352 297974
rect 514300 297910 514352 297916
rect 514864 295186 514892 372642
rect 514944 367260 514996 367266
rect 514944 367202 514996 367208
rect 514956 303210 514984 367202
rect 515128 360324 515180 360330
rect 515128 360266 515180 360272
rect 515036 353660 515088 353666
rect 515036 353602 515088 353608
rect 514944 303204 514996 303210
rect 514944 303146 514996 303152
rect 514852 295180 514904 295186
rect 514852 295122 514904 295128
rect 513564 292528 513616 292534
rect 513564 292470 513616 292476
rect 515048 291786 515076 353602
rect 515140 303278 515168 360266
rect 515220 352436 515272 352442
rect 515220 352378 515272 352384
rect 515232 305794 515260 352378
rect 515312 350940 515364 350946
rect 515312 350882 515364 350888
rect 515220 305788 515272 305794
rect 515220 305730 515272 305736
rect 515324 305726 515352 350882
rect 515416 319802 515444 599558
rect 515496 563100 515548 563106
rect 515496 563042 515548 563048
rect 515508 321774 515536 563042
rect 518912 520946 518940 600086
rect 518900 520940 518952 520946
rect 518900 520882 518952 520888
rect 518164 484424 518216 484430
rect 518164 484366 518216 484372
rect 515588 382356 515640 382362
rect 515588 382298 515640 382304
rect 515600 358494 515628 382298
rect 516784 378208 516836 378214
rect 516784 378150 516836 378156
rect 515680 374196 515732 374202
rect 515680 374138 515732 374144
rect 515588 358488 515640 358494
rect 515588 358430 515640 358436
rect 515496 321768 515548 321774
rect 515496 321710 515548 321716
rect 515404 319796 515456 319802
rect 515404 319738 515456 319744
rect 515312 305720 515364 305726
rect 515312 305662 515364 305668
rect 515128 303272 515180 303278
rect 515128 303214 515180 303220
rect 515692 295118 515720 374138
rect 516232 373788 516284 373794
rect 516232 373730 516284 373736
rect 516140 369980 516192 369986
rect 516140 369922 516192 369928
rect 515680 295112 515732 295118
rect 515680 295054 515732 295060
rect 516152 292126 516180 369922
rect 516244 300694 516272 373730
rect 516324 371816 516376 371822
rect 516324 371758 516376 371764
rect 516336 303074 516364 371758
rect 516508 356244 516560 356250
rect 516508 356186 516560 356192
rect 516416 331492 516468 331498
rect 516416 331434 516468 331440
rect 516324 303068 516376 303074
rect 516324 303010 516376 303016
rect 516232 300688 516284 300694
rect 516232 300630 516284 300636
rect 516140 292120 516192 292126
rect 516140 292062 516192 292068
rect 515036 291780 515088 291786
rect 515036 291722 515088 291728
rect 516428 289610 516456 331434
rect 516520 297906 516548 356186
rect 516600 349240 516652 349246
rect 516600 349182 516652 349188
rect 516612 300422 516640 349182
rect 516692 341148 516744 341154
rect 516692 341090 516744 341096
rect 516600 300416 516652 300422
rect 516600 300358 516652 300364
rect 516508 297900 516560 297906
rect 516508 297842 516560 297848
rect 516704 294846 516732 341090
rect 516796 321094 516824 378150
rect 516968 376780 517020 376786
rect 516968 376722 517020 376728
rect 516876 346588 516928 346594
rect 516876 346530 516928 346536
rect 516784 321088 516836 321094
rect 516784 321030 516836 321036
rect 516888 300354 516916 346530
rect 516980 316849 517008 376722
rect 517520 355156 517572 355162
rect 517520 355098 517572 355104
rect 516966 316840 517022 316849
rect 516966 316775 517022 316784
rect 516876 300348 516928 300354
rect 516876 300290 516928 300296
rect 516692 294840 516744 294846
rect 516692 294782 516744 294788
rect 517532 292398 517560 355098
rect 517612 353116 517664 353122
rect 517612 353058 517664 353064
rect 517624 297838 517652 353058
rect 517704 350668 517756 350674
rect 517704 350610 517756 350616
rect 517716 298042 517744 350610
rect 517796 348084 517848 348090
rect 517796 348026 517848 348032
rect 517808 300286 517836 348026
rect 517888 343188 517940 343194
rect 517888 343130 517940 343136
rect 517796 300280 517848 300286
rect 517796 300222 517848 300228
rect 517900 300218 517928 343130
rect 517980 341012 518032 341018
rect 517980 340954 518032 340960
rect 517992 300626 518020 340954
rect 518072 339584 518124 339590
rect 518072 339526 518124 339532
rect 517980 300620 518032 300626
rect 517980 300562 518032 300568
rect 518084 300490 518112 339526
rect 518176 321910 518204 484366
rect 518256 470620 518308 470626
rect 518256 470562 518308 470568
rect 518164 321904 518216 321910
rect 518164 321846 518216 321852
rect 518268 321842 518296 470562
rect 519542 465760 519598 465769
rect 519542 465695 519598 465704
rect 518348 383036 518400 383042
rect 518348 382978 518400 382984
rect 518360 358630 518388 382978
rect 518992 367396 519044 367402
rect 518992 367338 519044 367344
rect 518900 365764 518952 365770
rect 518900 365706 518952 365712
rect 518348 358624 518400 358630
rect 518348 358566 518400 358572
rect 518348 337068 518400 337074
rect 518348 337010 518400 337016
rect 518256 321836 518308 321842
rect 518256 321778 518308 321784
rect 518360 300558 518388 337010
rect 518348 300552 518400 300558
rect 518348 300494 518400 300500
rect 518072 300484 518124 300490
rect 518072 300426 518124 300432
rect 517888 300212 517940 300218
rect 517888 300154 517940 300160
rect 517704 298036 517756 298042
rect 517704 297978 517756 297984
rect 517612 297832 517664 297838
rect 517612 297774 517664 297780
rect 517520 292392 517572 292398
rect 517520 292334 517572 292340
rect 518912 292058 518940 365706
rect 519004 297566 519032 367338
rect 519084 361820 519136 361826
rect 519084 361762 519136 361768
rect 519096 297634 519124 361762
rect 519176 360460 519228 360466
rect 519176 360402 519228 360408
rect 519188 297702 519216 360402
rect 519268 358896 519320 358902
rect 519268 358838 519320 358844
rect 519280 297770 519308 358838
rect 519360 352028 519412 352034
rect 519360 351970 519412 351976
rect 519268 297764 519320 297770
rect 519268 297706 519320 297712
rect 519176 297696 519228 297702
rect 519176 297638 519228 297644
rect 519084 297628 519136 297634
rect 519084 297570 519136 297576
rect 518992 297560 519044 297566
rect 518992 297502 519044 297508
rect 519372 292262 519400 351970
rect 519452 346724 519504 346730
rect 519452 346666 519504 346672
rect 519464 292466 519492 346666
rect 519556 319870 519584 465695
rect 525812 464370 525840 600086
rect 538220 515432 538272 515438
rect 538220 515374 538272 515380
rect 535460 512644 535512 512650
rect 535460 512586 535512 512592
rect 532700 507884 532752 507890
rect 532700 507826 532752 507832
rect 529940 505164 529992 505170
rect 529940 505106 529992 505112
rect 529952 480254 529980 505106
rect 532712 480254 532740 507826
rect 535472 480254 535500 512586
rect 538232 480254 538260 515374
rect 529952 480226 530256 480254
rect 532712 480226 533200 480254
rect 535472 480226 536144 480254
rect 538232 480226 539088 480254
rect 525800 464364 525852 464370
rect 525800 464306 525852 464312
rect 527640 462528 527692 462534
rect 527640 462470 527692 462476
rect 521752 461644 521804 461650
rect 521752 461586 521804 461592
rect 521764 460972 521792 461586
rect 524432 460970 524722 460986
rect 527652 460972 527680 462470
rect 530228 460986 530256 480226
rect 533172 460986 533200 480226
rect 536116 460986 536144 480226
rect 539060 460986 539088 480226
rect 542372 464438 542400 702406
rect 559668 699825 559696 703520
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 573364 696992 573416 696998
rect 573364 696934 573416 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 567844 670744 567896 670750
rect 567844 670686 567896 670692
rect 545120 500268 545172 500274
rect 545120 500210 545172 500216
rect 542452 498840 542504 498846
rect 542452 498782 542504 498788
rect 542360 464432 542412 464438
rect 542360 464374 542412 464380
rect 542464 460986 542492 498782
rect 524420 460964 524722 460970
rect 524472 460958 524722 460964
rect 530228 460958 530610 460986
rect 533172 460958 533554 460986
rect 536116 460958 536498 460986
rect 539060 460958 539442 460986
rect 542386 460958 542492 460986
rect 545132 460986 545160 500210
rect 547880 496120 547932 496126
rect 547880 496062 547932 496068
rect 547892 460986 547920 496062
rect 554136 462460 554188 462466
rect 554136 462402 554188 462408
rect 551192 462392 551244 462398
rect 551192 462334 551244 462340
rect 545132 460958 545330 460986
rect 547892 460958 548274 460986
rect 551204 460972 551232 462334
rect 554148 460972 554176 462402
rect 524420 460906 524472 460912
rect 557538 442912 557594 442921
rect 557538 442847 557594 442856
rect 521212 421598 521240 425068
rect 522304 423496 522356 423502
rect 522304 423438 522356 423444
rect 521200 421592 521252 421598
rect 521200 421534 521252 421540
rect 522316 388958 522344 423438
rect 522500 423434 522528 425068
rect 523788 423570 523816 425068
rect 524708 425054 525090 425082
rect 523776 423564 523828 423570
rect 523776 423506 523828 423512
rect 522488 423428 522540 423434
rect 522488 423370 522540 423376
rect 523684 423428 523736 423434
rect 523684 423370 523736 423376
rect 522304 388952 522356 388958
rect 522304 388894 522356 388900
rect 523696 388890 523724 423370
rect 524708 412634 524736 425054
rect 526364 423366 526392 425068
rect 527284 425054 527666 425082
rect 526352 423360 526404 423366
rect 526352 423302 526404 423308
rect 526444 423360 526496 423366
rect 526444 423302 526496 423308
rect 524432 412606 524736 412634
rect 523684 388884 523736 388890
rect 523684 388826 523736 388832
rect 524432 388686 524460 412606
rect 526456 388822 526484 423302
rect 527284 412634 527312 425054
rect 528940 423298 528968 425068
rect 530228 423638 530256 425068
rect 529204 423632 529256 423638
rect 529204 423574 529256 423580
rect 530216 423632 530268 423638
rect 530216 423574 530268 423580
rect 530584 423632 530636 423638
rect 530584 423574 530636 423580
rect 528928 423292 528980 423298
rect 528928 423234 528980 423240
rect 527192 412606 527312 412634
rect 526444 388816 526496 388822
rect 526444 388758 526496 388764
rect 524420 388680 524472 388686
rect 524420 388622 524472 388628
rect 527192 388618 527220 412606
rect 527180 388612 527232 388618
rect 527180 388554 527232 388560
rect 529216 388550 529244 423574
rect 529204 388544 529256 388550
rect 529204 388486 529256 388492
rect 530596 388482 530624 423574
rect 531516 423230 531544 425068
rect 532804 423638 532832 425068
rect 532792 423632 532844 423638
rect 532792 423574 532844 423580
rect 531504 423224 531556 423230
rect 531504 423166 531556 423172
rect 534092 389842 534120 425068
rect 535012 425054 535394 425082
rect 536300 425054 536682 425082
rect 537588 425054 537970 425082
rect 538876 425054 539258 425082
rect 540164 425054 540546 425082
rect 535012 412634 535040 425054
rect 536300 412634 536328 425054
rect 537588 412634 537616 425054
rect 538876 412634 538904 425054
rect 540164 412634 540192 425054
rect 541820 420238 541848 425068
rect 542740 425054 543122 425082
rect 544028 425054 544410 425082
rect 541808 420232 541860 420238
rect 541808 420174 541860 420180
rect 542740 412634 542768 425054
rect 544028 412634 544056 425054
rect 545684 423162 545712 425068
rect 546604 425054 546986 425082
rect 545672 423156 545724 423162
rect 545672 423098 545724 423104
rect 546604 412634 546632 425054
rect 548260 423094 548288 425068
rect 549548 423502 549576 425068
rect 549536 423496 549588 423502
rect 549536 423438 549588 423444
rect 548248 423088 548300 423094
rect 548248 423030 548300 423036
rect 550836 423026 550864 425068
rect 552124 423434 552152 425068
rect 552112 423428 552164 423434
rect 552112 423370 552164 423376
rect 550824 423020 550876 423026
rect 550824 422962 550876 422968
rect 553412 422958 553440 425068
rect 554700 423366 554728 425068
rect 557552 424386 557580 442847
rect 557540 424380 557592 424386
rect 557540 424322 557592 424328
rect 554688 423360 554740 423366
rect 554688 423302 554740 423308
rect 553400 422952 553452 422958
rect 553400 422894 553452 422900
rect 534184 412606 535040 412634
rect 535472 412606 536328 412634
rect 536852 412606 537616 412634
rect 538232 412606 538904 412634
rect 539612 412606 540192 412634
rect 542372 412606 542768 412634
rect 543752 412606 544056 412634
rect 546512 412606 546632 412634
rect 534184 393990 534212 412606
rect 535472 395350 535500 412606
rect 536852 396778 536880 412606
rect 538232 398138 538260 412606
rect 539612 399498 539640 412606
rect 539600 399492 539652 399498
rect 539600 399434 539652 399440
rect 538220 398132 538272 398138
rect 538220 398074 538272 398080
rect 536840 396772 536892 396778
rect 536840 396714 536892 396720
rect 535460 395344 535512 395350
rect 535460 395286 535512 395292
rect 534172 393984 534224 393990
rect 534172 393926 534224 393932
rect 542372 391338 542400 412606
rect 543752 392698 543780 412606
rect 546512 400926 546540 412606
rect 546500 400920 546552 400926
rect 546500 400862 546552 400868
rect 543740 392692 543792 392698
rect 543740 392634 543792 392640
rect 542360 391332 542412 391338
rect 542360 391274 542412 391280
rect 534080 389836 534132 389842
rect 534080 389778 534132 389784
rect 530584 388476 530636 388482
rect 530584 388418 530636 388424
rect 553952 386572 554004 386578
rect 553952 386514 554004 386520
rect 534724 383784 534776 383790
rect 534724 383726 534776 383732
rect 519636 382492 519688 382498
rect 519636 382434 519688 382440
rect 519648 358698 519676 382434
rect 522304 378344 522356 378350
rect 522304 378286 522356 378292
rect 520280 375692 520332 375698
rect 520280 375634 520332 375640
rect 519636 358692 519688 358698
rect 519636 358634 519688 358640
rect 519636 339652 519688 339658
rect 519636 339594 519688 339600
rect 519544 319864 519596 319870
rect 519544 319806 519596 319812
rect 519648 294710 519676 339594
rect 519728 336932 519780 336938
rect 519728 336874 519780 336880
rect 519740 294914 519768 336874
rect 519728 294908 519780 294914
rect 519728 294850 519780 294856
rect 520292 294778 520320 375634
rect 521660 372768 521712 372774
rect 521660 372710 521712 372716
rect 520372 370116 520424 370122
rect 520372 370058 520424 370064
rect 520384 294982 520412 370058
rect 520464 368552 520516 368558
rect 520464 368494 520516 368500
rect 520476 295050 520504 368494
rect 520556 365900 520608 365906
rect 520556 365842 520608 365848
rect 520568 297498 520596 365842
rect 520648 349580 520700 349586
rect 520648 349522 520700 349528
rect 520556 297492 520608 297498
rect 520556 297434 520608 297440
rect 520464 295044 520516 295050
rect 520464 294986 520516 294992
rect 520372 294976 520424 294982
rect 520372 294918 520424 294924
rect 520280 294772 520332 294778
rect 520280 294714 520332 294720
rect 519636 294704 519688 294710
rect 519636 294646 519688 294652
rect 519452 292460 519504 292466
rect 519452 292402 519504 292408
rect 519360 292256 519412 292262
rect 519360 292198 519412 292204
rect 520660 292194 520688 349522
rect 520740 343732 520792 343738
rect 520740 343674 520792 343680
rect 520752 292330 520780 343674
rect 520832 338292 520884 338298
rect 520832 338234 520884 338240
rect 520844 294642 520872 338234
rect 520832 294636 520884 294642
rect 520832 294578 520884 294584
rect 520740 292324 520792 292330
rect 520740 292266 520792 292272
rect 520648 292188 520700 292194
rect 520648 292130 520700 292136
rect 518900 292052 518952 292058
rect 518900 291994 518952 292000
rect 516416 289604 516468 289610
rect 516416 289546 516468 289552
rect 521672 289338 521700 372710
rect 521752 361616 521804 361622
rect 521752 361558 521804 361564
rect 521764 291990 521792 361558
rect 522316 360874 522344 378286
rect 523040 364404 523092 364410
rect 523040 364346 523092 364352
rect 522304 360868 522356 360874
rect 522304 360810 522356 360816
rect 521844 342304 521896 342310
rect 521844 342246 521896 342252
rect 521752 291984 521804 291990
rect 521752 291926 521804 291932
rect 521660 289332 521712 289338
rect 521660 289274 521712 289280
rect 521856 289270 521884 342246
rect 521936 339516 521988 339522
rect 521936 339458 521988 339464
rect 521844 289264 521896 289270
rect 521844 289206 521896 289212
rect 521948 289134 521976 339458
rect 522028 338156 522080 338162
rect 522028 338098 522080 338104
rect 522040 289202 522068 338098
rect 523052 291922 523080 364346
rect 523132 360392 523184 360398
rect 523132 360334 523184 360340
rect 523040 291916 523092 291922
rect 523040 291858 523092 291864
rect 523144 291854 523172 360334
rect 534736 358902 534764 383726
rect 547144 383716 547196 383722
rect 547144 383658 547196 383664
rect 544384 379568 544436 379574
rect 544384 379510 544436 379516
rect 544396 359038 544424 379510
rect 544384 359032 544436 359038
rect 544384 358974 544436 358980
rect 547156 358970 547184 383658
rect 548524 380928 548576 380934
rect 548524 380870 548576 380876
rect 547236 376032 547288 376038
rect 547236 375974 547288 375980
rect 547144 358964 547196 358970
rect 547144 358906 547196 358912
rect 534724 358896 534776 358902
rect 534724 358838 534776 358844
rect 547248 358562 547276 375974
rect 548536 359106 548564 380870
rect 548616 378276 548668 378282
rect 548616 378218 548668 378224
rect 548628 360194 548656 378218
rect 553964 377890 553992 386514
rect 563428 385144 563480 385150
rect 563428 385086 563480 385092
rect 553964 377862 554438 377890
rect 563440 377876 563468 385086
rect 549904 377460 549956 377466
rect 549904 377402 549956 377408
rect 548616 360188 548668 360194
rect 548616 360130 548668 360136
rect 548524 359100 548576 359106
rect 548524 359042 548576 359048
rect 549916 358766 549944 377402
rect 550640 360868 550692 360874
rect 550640 360810 550692 360816
rect 550652 360754 550680 360810
rect 550652 360726 550850 360754
rect 552032 360194 552322 360210
rect 552020 360188 552322 360194
rect 552072 360182 552322 360188
rect 552020 360130 552072 360136
rect 553780 359038 553808 360060
rect 553768 359032 553820 359038
rect 553768 358974 553820 358980
rect 555252 358834 555280 360060
rect 555240 358828 555292 358834
rect 555240 358770 555292 358776
rect 556724 358766 556752 360060
rect 558196 359106 558224 360060
rect 558184 359100 558236 359106
rect 558184 359042 558236 359048
rect 549904 358760 549956 358766
rect 549904 358702 549956 358708
rect 556712 358760 556764 358766
rect 556712 358702 556764 358708
rect 559668 358562 559696 360060
rect 547236 358556 547288 358562
rect 547236 358498 547288 358504
rect 559656 358556 559708 358562
rect 559656 358498 559708 358504
rect 561140 358494 561168 360060
rect 562612 358630 562640 360060
rect 564084 358698 564112 360060
rect 565556 358970 565584 360060
rect 565544 358964 565596 358970
rect 565544 358906 565596 358912
rect 567028 358902 567056 360060
rect 567016 358896 567068 358902
rect 567016 358838 567068 358844
rect 564072 358692 564124 358698
rect 564072 358634 564124 358640
rect 562600 358624 562652 358630
rect 562600 358566 562652 358572
rect 561128 358488 561180 358494
rect 561128 358430 561180 358436
rect 567856 321706 567884 670686
rect 569224 364404 569276 364410
rect 569224 364346 569276 364352
rect 567844 321700 567896 321706
rect 567844 321642 567896 321648
rect 569236 321366 569264 364346
rect 569224 321360 569276 321366
rect 569224 321302 569276 321308
rect 573376 321298 573404 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 576124 683188 576176 683194
rect 576124 683130 576176 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 574744 630692 574796 630698
rect 574744 630634 574796 630640
rect 574756 321434 574784 630634
rect 576136 321502 576164 683130
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580262 617536 580318 617545
rect 580262 617471 580318 617480
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 579894 564360 579950 564369
rect 579894 564295 579950 564304
rect 579908 563106 579936 564295
rect 579896 563100 579948 563106
rect 579896 563042 579948 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 352164 580224 352170
rect 580172 352106 580224 352112
rect 580184 351937 580212 352106
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 576124 321496 576176 321502
rect 576124 321438 576176 321444
rect 574744 321428 574796 321434
rect 574744 321370 574796 321376
rect 573364 321292 573416 321298
rect 573364 321234 573416 321240
rect 580184 320006 580212 325207
rect 580276 321638 580304 617471
rect 580368 599622 580396 643991
rect 580356 599616 580408 599622
rect 580356 599558 580408 599564
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580264 321632 580316 321638
rect 580264 321574 580316 321580
rect 580368 320074 580396 577623
rect 580446 524512 580502 524521
rect 580446 524447 580502 524456
rect 580460 322250 580488 524447
rect 580538 511320 580594 511329
rect 580538 511255 580594 511264
rect 580448 322244 580500 322250
rect 580448 322186 580500 322192
rect 580552 321570 580580 511255
rect 580630 458144 580686 458153
rect 580630 458079 580686 458088
rect 580540 321564 580592 321570
rect 580540 321506 580592 321512
rect 580644 320890 580672 458079
rect 580722 431624 580778 431633
rect 580722 431559 580778 431568
rect 580736 320958 580764 431559
rect 580814 418296 580870 418305
rect 580814 418231 580870 418240
rect 580724 320952 580776 320958
rect 580724 320894 580776 320900
rect 580632 320884 580684 320890
rect 580632 320826 580684 320832
rect 580356 320068 580408 320074
rect 580356 320010 580408 320016
rect 580172 320000 580224 320006
rect 580172 319942 580224 319948
rect 530676 319524 530728 319530
rect 530676 319466 530728 319472
rect 530584 319388 530636 319394
rect 530584 319330 530636 319336
rect 529940 317144 529992 317150
rect 529940 317086 529992 317092
rect 529204 308440 529256 308446
rect 529204 308382 529256 308388
rect 523132 291848 523184 291854
rect 523132 291790 523184 291796
rect 522028 289196 522080 289202
rect 522028 289138 522080 289144
rect 521936 289128 521988 289134
rect 521936 289070 521988 289076
rect 529216 287054 529244 308382
rect 529216 287026 529336 287054
rect 512736 269816 512788 269822
rect 512736 269758 512788 269764
rect 490288 268456 490340 268462
rect 490288 268398 490340 268404
rect 496912 268456 496964 268462
rect 496912 268398 496964 268404
rect 466552 268388 466604 268394
rect 466552 268330 466604 268336
rect 460572 267028 460624 267034
rect 460572 266970 460624 266976
rect 529308 261633 529336 287026
rect 529294 261624 529350 261633
rect 529294 261559 529350 261568
rect 529952 209273 529980 317086
rect 530032 307216 530084 307222
rect 530032 307158 530084 307164
rect 530044 226250 530072 307158
rect 530122 226264 530178 226273
rect 530044 226222 530122 226250
rect 530122 226199 530178 226208
rect 529938 209264 529994 209273
rect 529938 209199 529994 209208
rect 481640 200796 481692 200802
rect 481640 200738 481692 200744
rect 460480 152992 460532 152998
rect 460480 152934 460532 152940
rect 481652 151814 481680 200738
rect 485780 198008 485832 198014
rect 485780 197950 485832 197956
rect 483664 160132 483716 160138
rect 483664 160074 483716 160080
rect 481652 151786 481864 151814
rect 481836 139890 481864 151786
rect 483676 142934 483704 160074
rect 483664 142928 483716 142934
rect 483664 142870 483716 142876
rect 485792 139890 485820 197950
rect 524420 171828 524472 171834
rect 524420 171770 524472 171776
rect 489920 162172 489972 162178
rect 489920 162114 489972 162120
rect 489932 139890 489960 162114
rect 496820 161832 496872 161838
rect 496820 161774 496872 161780
rect 494060 161696 494112 161702
rect 494060 161638 494112 161644
rect 494072 139890 494100 161638
rect 496832 151814 496860 161774
rect 500960 161764 501012 161770
rect 500960 161706 501012 161712
rect 500972 151814 501000 161706
rect 505100 161628 505152 161634
rect 505100 161570 505152 161576
rect 505112 151814 505140 161570
rect 513380 161560 513432 161566
rect 513380 161502 513432 161508
rect 513392 151814 513420 161502
rect 517520 161492 517572 161498
rect 517520 161434 517572 161440
rect 496832 151786 497688 151814
rect 500972 151786 501644 151814
rect 505112 151786 505600 151814
rect 513392 151786 513512 151814
rect 497660 139890 497688 151786
rect 501616 139890 501644 151786
rect 505572 139890 505600 151786
rect 509608 142860 509660 142866
rect 509608 142802 509660 142808
rect 509620 139890 509648 142802
rect 513484 139890 513512 151786
rect 517532 139890 517560 161434
rect 521660 160744 521712 160750
rect 521660 160686 521712 160692
rect 521672 139890 521700 160686
rect 524432 151814 524460 171770
rect 528560 163532 528612 163538
rect 528560 163474 528612 163480
rect 528572 151814 528600 163474
rect 524432 151786 525380 151814
rect 528572 151786 529336 151814
rect 525352 139890 525380 151786
rect 529308 139890 529336 151786
rect 530596 140078 530624 319330
rect 530688 140146 530716 319466
rect 538864 319456 538916 319462
rect 538864 319398 538916 319404
rect 536840 307148 536892 307154
rect 536840 307090 536892 307096
rect 531320 287700 531372 287706
rect 531320 287642 531372 287648
rect 531332 243681 531360 287642
rect 531318 243672 531374 243681
rect 531318 243607 531374 243616
rect 536852 151814 536880 307090
rect 537484 300756 537536 300762
rect 537484 300698 537536 300704
rect 537496 167006 537524 300698
rect 537484 167000 537536 167006
rect 537484 166942 537536 166948
rect 536852 151786 537248 151814
rect 533988 142928 534040 142934
rect 533988 142870 534040 142876
rect 534000 142186 534028 142870
rect 533988 142180 534040 142186
rect 533988 142122 534040 142128
rect 530676 140140 530728 140146
rect 530676 140082 530728 140088
rect 530584 140072 530636 140078
rect 530584 140014 530636 140020
rect 534000 139890 534028 142122
rect 481836 139862 482264 139890
rect 485792 139862 486220 139890
rect 489932 139862 490176 139890
rect 494072 139862 494132 139890
rect 497660 139862 498088 139890
rect 501616 139862 502044 139890
rect 505572 139862 506000 139890
rect 509620 139862 509956 139890
rect 513484 139862 513912 139890
rect 517532 139862 517868 139890
rect 521672 139862 521824 139890
rect 525352 139862 525780 139890
rect 529308 139862 529736 139890
rect 533692 139862 534028 139890
rect 537220 139890 537248 151786
rect 537220 139862 537648 139890
rect 538876 139262 538904 319398
rect 580828 319258 580856 418231
rect 580816 319252 580868 319258
rect 580816 319194 580868 319200
rect 540336 318300 540388 318306
rect 540336 318242 540388 318248
rect 539692 317280 539744 317286
rect 539692 317222 539744 317228
rect 538956 314152 539008 314158
rect 538956 314094 539008 314100
rect 538864 139256 538916 139262
rect 538864 139198 538916 139204
rect 538968 136610 538996 314094
rect 539600 309868 539652 309874
rect 539600 309810 539652 309816
rect 539048 280832 539100 280838
rect 539048 280774 539100 280780
rect 539060 151814 539088 280774
rect 539060 151786 539364 151814
rect 539336 137737 539364 151786
rect 539322 137728 539378 137737
rect 539322 137663 539378 137672
rect 538956 136604 539008 136610
rect 538956 136546 539008 136552
rect 539508 136604 539560 136610
rect 539508 136546 539560 136552
rect 539520 135969 539548 136546
rect 539506 135960 539562 135969
rect 539506 135895 539562 135904
rect 539612 86873 539640 309810
rect 539704 113257 539732 317222
rect 539876 284980 539928 284986
rect 539876 284922 539928 284928
rect 539784 142180 539836 142186
rect 539784 142122 539836 142128
rect 539690 113248 539746 113257
rect 539690 113183 539746 113192
rect 539598 86864 539654 86873
rect 539598 86799 539654 86808
rect 537484 62824 537536 62830
rect 537484 62766 537536 62772
rect 460388 46844 460440 46850
rect 460388 46786 460440 46792
rect 537496 41041 537524 62766
rect 537482 41032 537538 41041
rect 537482 40967 537538 40976
rect 460204 39772 460256 39778
rect 460204 39714 460256 39720
rect 539796 33697 539824 142122
rect 539888 99249 539916 284922
rect 540152 279472 540204 279478
rect 540152 279414 540204 279420
rect 539968 276684 540020 276690
rect 539968 276626 540020 276632
rect 539980 108769 540008 276626
rect 540060 271244 540112 271250
rect 540060 271186 540112 271192
rect 539966 108760 540022 108769
rect 539966 108695 540022 108704
rect 540072 104689 540100 271186
rect 540164 115025 540192 279414
rect 540244 272536 540296 272542
rect 540244 272478 540296 272484
rect 540256 121145 540284 272478
rect 540348 123185 540376 318242
rect 540980 318232 541032 318238
rect 540980 318174 541032 318180
rect 540334 123176 540390 123185
rect 540334 123111 540390 123120
rect 540242 121136 540298 121145
rect 540242 121071 540298 121080
rect 540150 115016 540206 115025
rect 540150 114951 540206 114960
rect 540058 104680 540114 104689
rect 540058 104615 540114 104624
rect 539874 99240 539930 99249
rect 539874 99175 539930 99184
rect 540992 82385 541020 318174
rect 543096 317212 543148 317218
rect 543096 317154 543148 317160
rect 541072 315376 541124 315382
rect 541072 315318 541124 315324
rect 541084 119105 541112 315318
rect 543004 314084 543056 314090
rect 543004 314026 543056 314032
rect 542728 311228 542780 311234
rect 542728 311170 542780 311176
rect 541440 278044 541492 278050
rect 541440 277986 541492 277992
rect 541256 275324 541308 275330
rect 541256 275266 541308 275272
rect 541164 273964 541216 273970
rect 541164 273906 541216 273912
rect 541070 119096 541126 119105
rect 541070 119031 541126 119040
rect 541176 92585 541204 273906
rect 541268 102785 541296 275266
rect 541348 274032 541400 274038
rect 541348 273974 541400 273980
rect 541360 106865 541388 273974
rect 541452 110945 541480 277986
rect 541532 271176 541584 271182
rect 541532 271118 541584 271124
rect 541544 117065 541572 271118
rect 542636 268456 542688 268462
rect 542636 268398 542688 268404
rect 542544 140140 542596 140146
rect 542544 140082 542596 140088
rect 542452 140072 542504 140078
rect 542452 140014 542504 140020
rect 541530 117056 541586 117065
rect 541530 116991 541586 117000
rect 541438 110936 541494 110945
rect 541438 110871 541494 110880
rect 541346 106856 541402 106865
rect 541346 106791 541402 106800
rect 541254 102776 541310 102785
rect 541254 102711 541310 102720
rect 542464 100745 542492 140014
rect 542450 100736 542506 100745
rect 542450 100671 542506 100680
rect 542556 96665 542584 140082
rect 542542 96656 542598 96665
rect 542542 96591 542598 96600
rect 541162 92576 541218 92585
rect 541162 92511 541218 92520
rect 542648 90545 542676 268398
rect 542740 133385 542768 311170
rect 542912 309800 542964 309806
rect 542912 309742 542964 309748
rect 542820 269952 542872 269958
rect 542820 269894 542872 269900
rect 542726 133376 542782 133385
rect 542726 133311 542782 133320
rect 542832 94625 542860 269894
rect 542818 94616 542874 94625
rect 542818 94551 542874 94560
rect 542634 90536 542690 90545
rect 542634 90471 542690 90480
rect 542924 88505 542952 309742
rect 543016 125225 543044 314026
rect 543108 129305 543136 317154
rect 562324 315308 562376 315314
rect 562324 315250 562376 315256
rect 548524 313948 548576 313954
rect 548524 313890 548576 313896
rect 544384 312588 544436 312594
rect 544384 312530 544436 312536
rect 543740 270020 543792 270026
rect 543740 269962 543792 269968
rect 543188 139256 543240 139262
rect 543188 139198 543240 139204
rect 543200 131345 543228 139198
rect 543278 137864 543334 137873
rect 543278 137799 543334 137808
rect 543186 131336 543242 131345
rect 543186 131271 543242 131280
rect 543094 129296 543150 129305
rect 543094 129231 543150 129240
rect 543292 127265 543320 137799
rect 543278 127256 543334 127265
rect 543278 127191 543334 127200
rect 543002 125216 543058 125225
rect 543002 125151 543058 125160
rect 542910 88496 542966 88505
rect 542910 88431 542966 88440
rect 540978 82376 541034 82385
rect 540978 82311 541034 82320
rect 543752 51134 543780 269962
rect 544396 60722 544424 312530
rect 547144 311160 547196 311166
rect 547144 311102 547196 311108
rect 547156 153202 547184 311102
rect 547144 153196 547196 153202
rect 547144 153138 547196 153144
rect 548536 73166 548564 313890
rect 559564 293276 559616 293282
rect 559564 293218 559616 293224
rect 551284 290488 551336 290494
rect 551284 290430 551336 290436
rect 551296 193186 551324 290430
rect 554044 282192 554096 282198
rect 554044 282134 554096 282140
rect 551284 193180 551336 193186
rect 551284 193122 551336 193128
rect 554056 139398 554084 282134
rect 555424 268388 555476 268394
rect 555424 268330 555476 268336
rect 555436 179382 555464 268330
rect 559576 219434 559604 293218
rect 559564 219428 559616 219434
rect 559564 219370 559616 219376
rect 555424 179376 555476 179382
rect 555424 179318 555476 179324
rect 554044 139392 554096 139398
rect 554044 139334 554096 139340
rect 548524 73160 548576 73166
rect 548524 73102 548576 73108
rect 544384 60716 544436 60722
rect 544384 60658 544436 60664
rect 540612 51128 540664 51134
rect 540612 51070 540664 51076
rect 543740 51128 543792 51134
rect 543740 51070 543792 51076
rect 540624 48929 540652 51070
rect 540610 48920 540666 48929
rect 540610 48855 540666 48864
rect 539782 33688 539838 33697
rect 539782 33623 539838 33632
rect 562336 6866 562364 315250
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 566464 307080 566516 307086
rect 566464 307022 566516 307028
rect 565084 306128 565136 306134
rect 565084 306070 565136 306076
rect 563704 304428 563756 304434
rect 563704 304370 563756 304376
rect 563716 46918 563744 304370
rect 563704 46912 563756 46918
rect 563704 46854 563756 46860
rect 565096 33114 565124 306070
rect 565084 33108 565136 33114
rect 565084 33050 565136 33056
rect 566476 20670 566504 307022
rect 574744 303000 574796 303006
rect 574744 302942 574796 302948
rect 571984 295996 572036 296002
rect 571984 295938 572036 295944
rect 569224 291712 569276 291718
rect 569224 291654 569276 291660
rect 569236 100706 569264 291654
rect 570604 289672 570656 289678
rect 570604 289614 570656 289620
rect 570616 233238 570644 289614
rect 571996 245614 572024 295938
rect 573364 294568 573416 294574
rect 573364 294510 573416 294516
rect 571984 245608 572036 245614
rect 571984 245550 572036 245556
rect 570604 233232 570656 233238
rect 570604 233174 570656 233180
rect 573376 113150 573404 294510
rect 573364 113144 573416 113150
rect 573364 113086 573416 113092
rect 569224 100700 569276 100706
rect 569224 100642 569276 100648
rect 574756 86970 574784 302942
rect 576124 301504 576176 301510
rect 576124 301446 576176 301452
rect 576136 126954 576164 301446
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 578884 298104 578936 298110
rect 578884 298046 578936 298052
rect 578896 205737 578924 298046
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580264 269884 580316 269890
rect 580264 269826 580316 269832
rect 580276 258913 580304 269826
rect 580262 258904 580318 258913
rect 580262 258839 580318 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 578882 205728 578938 205737
rect 578882 205663 578938 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 576124 126948 576176 126954
rect 576124 126890 576176 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 574744 86964 574796 86970
rect 574744 86906 574796 86912
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 566464 20664 566516 20670
rect 566464 20606 566516 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 562324 6860 562376 6866
rect 562324 6802 562376 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 458824 4004 458876 4010
rect 458824 3946 458876 3952
rect 456064 3732 456116 3738
rect 456064 3674 456116 3680
rect 454682 3360 454738 3369
rect 454682 3295 454738 3304
rect 453304 2100 453356 2106
rect 453304 2042 453356 2048
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 40498 700304 40554 700360
rect 202786 700440 202842 700496
rect 153198 692008 153254 692064
rect 136638 689288 136694 689344
rect 282918 690648 282974 690704
rect 3422 684256 3478 684312
rect 3238 579944 3294 580000
rect 3330 566888 3386 566944
rect 3514 671200 3570 671256
rect 3514 669840 3570 669896
rect 3422 462576 3478 462632
rect 3698 632032 3754 632088
rect 3606 475632 3662 475688
rect 3514 449520 3570 449576
rect 4066 553832 4122 553888
rect 3974 527856 4030 527912
rect 3882 514800 3938 514856
rect 361762 678988 361764 679008
rect 361764 678988 361816 679008
rect 361816 678988 361818 679008
rect 361762 678952 361818 678988
rect 361762 667956 361818 667992
rect 361762 667936 361764 667956
rect 361764 667936 361816 667956
rect 361816 667936 361818 667956
rect 361762 656940 361818 656976
rect 361762 656920 361764 656940
rect 361764 656920 361816 656940
rect 361816 656920 361818 656940
rect 361762 645924 361818 645960
rect 361762 645904 361764 645924
rect 361764 645904 361816 645924
rect 361816 645904 361818 645924
rect 361578 634888 361634 634944
rect 361578 623872 361634 623928
rect 361578 612856 361634 612912
rect 361578 601840 361634 601896
rect 361762 590824 361818 590880
rect 361762 579808 361818 579864
rect 361578 568812 361634 568848
rect 361578 568792 361580 568812
rect 361580 568792 361632 568812
rect 361632 568792 361634 568812
rect 361578 557796 361634 557832
rect 361578 557776 361580 557796
rect 361580 557776 361632 557796
rect 361632 557776 361634 557796
rect 361762 546760 361818 546816
rect 361762 535744 361818 535800
rect 361762 524728 361818 524784
rect 3790 501744 3846 501800
rect 3698 423544 3754 423600
rect 361762 513712 361818 513768
rect 361762 502696 361818 502752
rect 361762 491680 361818 491736
rect 361762 480664 361818 480720
rect 361762 469648 361818 469704
rect 361762 458632 361818 458688
rect 361578 447616 361634 447672
rect 362222 436600 362278 436656
rect 362314 425584 362370 425640
rect 361578 414568 361634 414624
rect 3974 410488 4030 410544
rect 361578 403552 361634 403608
rect 3790 397432 3846 397488
rect 3606 358400 3662 358456
rect 3514 345344 3570 345400
rect 3422 306176 3478 306232
rect 3330 149776 3386 149832
rect 3238 136720 3294 136776
rect 3606 293120 3662 293176
rect 3606 267144 3662 267200
rect 3514 254088 3570 254144
rect 3422 71576 3478 71632
rect 3698 241032 3754 241088
rect 3606 58520 3662 58576
rect 361578 392536 361634 392592
rect 361578 381520 361634 381576
rect 3974 371320 4030 371376
rect 3882 319232 3938 319288
rect 3882 214920 3938 214976
rect 3790 201864 3846 201920
rect 361578 370504 361634 370560
rect 362222 359488 362278 359544
rect 361762 348472 361818 348528
rect 361762 337456 361818 337512
rect 362222 326440 362278 326496
rect 361762 315424 361818 315480
rect 3974 188808 4030 188864
rect 4066 162832 4122 162888
rect 19338 49544 19394 49600
rect 3422 45484 3478 45520
rect 3422 45464 3424 45484
rect 3424 45464 3476 45484
rect 3476 45464 3478 45484
rect 20902 59880 20958 59936
rect 21454 59880 21510 59936
rect 20902 49408 20958 49464
rect 27618 44920 27674 44976
rect 6918 44784 6974 44840
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 1674 3440 1730 3496
rect 570 3304 626 3360
rect 5262 3848 5318 3904
rect 6458 3712 6514 3768
rect 8758 3576 8814 3632
rect 26238 39208 26294 39264
rect 121458 39344 121514 39400
rect 361762 304408 361818 304464
rect 359646 46280 359702 46336
rect 361762 293392 361818 293448
rect 361762 282376 361818 282432
rect 361762 271360 361818 271416
rect 361762 260344 361818 260400
rect 361762 249328 361818 249384
rect 361762 238312 361818 238368
rect 361762 227296 361818 227352
rect 361578 216316 361580 216336
rect 361580 216316 361632 216336
rect 361632 216316 361634 216336
rect 361578 216280 361634 216316
rect 361762 205264 361818 205320
rect 361670 194248 361726 194304
rect 361670 183232 361726 183288
rect 361762 172216 361818 172272
rect 361762 161200 361818 161256
rect 361762 139168 361818 139224
rect 361210 46416 361266 46472
rect 361578 128188 361580 128208
rect 361580 128188 361632 128208
rect 361632 128188 361634 128208
rect 361578 128152 361634 128188
rect 361578 117136 361634 117192
rect 361578 106120 361634 106176
rect 361762 95140 361764 95160
rect 361764 95140 361816 95160
rect 361816 95140 361818 95160
rect 361762 95104 361818 95140
rect 361762 84124 361764 84144
rect 361764 84124 361816 84144
rect 361816 84124 361818 84144
rect 361762 84088 361818 84124
rect 361762 73108 361764 73128
rect 361764 73108 361816 73128
rect 361816 73108 361818 73128
rect 361762 73072 361818 73108
rect 361762 62076 361818 62112
rect 361762 62056 361764 62076
rect 361764 62056 361816 62076
rect 361816 62056 361818 62076
rect 361762 51040 361818 51096
rect 362406 150184 362462 150240
rect 362222 3848 362278 3904
rect 368202 44920 368258 44976
rect 378782 294480 378838 294536
rect 370870 289040 370926 289096
rect 376390 291760 376446 291816
rect 381634 294752 381690 294808
rect 381818 294616 381874 294672
rect 420274 684528 420330 684584
rect 442906 420144 442962 420200
rect 424138 335416 424194 335472
rect 420734 334464 420790 334520
rect 428094 334464 428150 334520
rect 429198 332968 429254 333024
rect 395342 300464 395398 300520
rect 392582 300056 392638 300112
rect 389822 297336 389878 297392
rect 367742 3712 367798 3768
rect 392582 3576 392638 3632
rect 395526 300192 395582 300248
rect 395710 300328 395766 300384
rect 403898 302776 403954 302832
rect 432602 332832 432658 332888
rect 421378 162696 421434 162752
rect 426162 162696 426218 162752
rect 428646 162696 428702 162752
rect 432694 325488 432750 325544
rect 432602 318144 432658 318200
rect 432970 329160 433026 329216
rect 432786 321816 432842 321872
rect 432694 314472 432750 314528
rect 432602 310800 432658 310856
rect 432418 307128 432474 307184
rect 444194 422864 444250 422920
rect 444286 421912 444342 421968
rect 445390 683304 445446 683360
rect 445206 321680 445262 321736
rect 446310 682760 446366 682816
rect 445666 387640 445722 387696
rect 446310 321544 446366 321600
rect 446586 319640 446642 319696
rect 446862 683168 446918 683224
rect 446770 320048 446826 320104
rect 447966 514392 448022 514448
rect 447414 512760 447470 512816
rect 447966 505144 448022 505200
rect 447138 383580 447194 383616
rect 447138 383560 447140 383580
rect 447140 383560 447192 383580
rect 447192 383560 447194 383580
rect 447138 382200 447194 382256
rect 447138 380840 447194 380896
rect 447138 378800 447194 378856
rect 447138 377440 447194 377496
rect 447138 376080 447194 376136
rect 447138 374720 447194 374776
rect 447138 373360 447194 373416
rect 447138 372000 447194 372056
rect 447138 370640 447194 370696
rect 447138 369280 447194 369336
rect 447138 367920 447194 367976
rect 447138 365880 447194 365936
rect 447138 364520 447194 364576
rect 447138 363160 447194 363216
rect 447138 361800 447194 361856
rect 447138 361120 447194 361176
rect 447138 359080 447194 359136
rect 447138 350920 447194 350976
rect 447138 347520 447194 347576
rect 447322 382880 447378 382936
rect 447322 381520 447378 381576
rect 447322 379480 447378 379536
rect 447322 376760 447378 376816
rect 447322 375400 447378 375456
rect 447322 374040 447378 374096
rect 447322 372680 447378 372736
rect 447322 371320 447378 371376
rect 447322 369960 447378 370016
rect 447322 368600 447378 368656
rect 447322 367240 447378 367296
rect 447322 366560 447378 366616
rect 447322 365200 447378 365256
rect 447322 363840 447378 363896
rect 447322 362480 447378 362536
rect 447322 360440 447378 360496
rect 447322 359760 447378 359816
rect 447322 344120 447378 344176
rect 447230 342080 447286 342136
rect 447138 341400 447194 341456
rect 447138 340720 447194 340776
rect 447230 340040 447286 340096
rect 447230 339360 447286 339416
rect 447138 338680 447194 338736
rect 447230 338000 447286 338056
rect 447138 337320 447194 337376
rect 447230 336640 447286 336696
rect 447138 335960 447194 336016
rect 447230 334600 447286 334656
rect 447138 333920 447194 333976
rect 447230 333240 447286 333296
rect 447138 331880 447194 331936
rect 447230 331200 447286 331256
rect 447138 330556 447140 330576
rect 447140 330556 447192 330576
rect 447192 330556 447194 330576
rect 447138 330520 447194 330556
rect 447138 329160 447194 329216
rect 448150 516704 448206 516760
rect 448334 512760 448390 512816
rect 448518 514392 448574 514448
rect 448150 507728 448206 507784
rect 448058 501880 448114 501936
rect 447506 380160 447562 380216
rect 447506 378120 447562 378176
rect 447874 353640 447930 353696
rect 447782 352280 447838 352336
rect 447506 343440 447562 343496
rect 447506 335280 447562 335336
rect 447414 332560 447470 332616
rect 447414 328480 447470 328536
rect 447598 329840 447654 329896
rect 447506 327800 447562 327856
rect 447414 326440 447470 326496
rect 447966 325760 448022 325816
rect 448426 510448 448482 510504
rect 448334 503376 448390 503432
rect 448426 358400 448482 358456
rect 449070 386960 449126 387016
rect 448978 357720 449034 357776
rect 449070 355680 449126 355736
rect 448426 344800 448482 344856
rect 448426 332560 448482 332616
rect 448334 328480 448390 328536
rect 448242 327120 448298 327176
rect 448242 325080 448298 325136
rect 449806 503376 449862 503432
rect 449898 496068 449900 496088
rect 449900 496068 449952 496088
rect 449952 496068 449954 496088
rect 449898 496032 449954 496068
rect 449438 387096 449494 387152
rect 449530 385600 449586 385656
rect 449438 354320 449494 354376
rect 449622 356360 449678 356416
rect 449806 357040 449862 357096
rect 449714 355000 449770 355056
rect 449898 351056 449954 351112
rect 449714 350240 449770 350296
rect 449622 345480 449678 345536
rect 449530 324400 449586 324456
rect 449806 343440 449862 343496
rect 449990 349968 450046 350024
rect 450266 353232 450322 353288
rect 450358 348608 450414 348664
rect 450174 347248 450230 347304
rect 450082 346296 450138 346352
rect 478510 700440 478566 700496
rect 494794 700304 494850 700360
rect 527178 699760 527234 699816
rect 462318 669840 462374 669896
rect 457810 667936 457866 667992
rect 457718 653248 457774 653304
rect 457626 650800 457682 650856
rect 457534 645904 457590 645960
rect 457442 621424 457498 621480
rect 457350 616528 457406 616584
rect 457258 609184 457314 609240
rect 458086 660592 458142 660648
rect 457994 658144 458050 658200
rect 457902 641008 457958 641064
rect 459190 655696 459246 655752
rect 459098 648352 459154 648408
rect 459006 643456 459062 643512
rect 458914 638560 458970 638616
rect 458822 618976 458878 619032
rect 458638 611632 458694 611688
rect 458914 598168 458970 598224
rect 459466 631216 459522 631272
rect 459282 628768 459338 628824
rect 459190 601840 459246 601896
rect 459098 599528 459154 599584
rect 459006 596944 459062 597000
rect 458730 596808 458786 596864
rect 459374 626320 459430 626376
rect 459558 623804 459614 623860
rect 459650 614080 459706 614136
rect 459742 606668 459798 606724
rect 459834 604220 459890 604276
rect 459466 522280 459522 522336
rect 450634 516296 450690 516352
rect 462962 517520 463018 517576
rect 467194 519424 467250 519480
rect 491850 516180 491906 516216
rect 491850 516160 491852 516180
rect 491852 516160 491904 516180
rect 491904 516160 491906 516180
rect 494150 516704 494206 516760
rect 494150 515888 494206 515944
rect 494334 516704 494390 516760
rect 494150 512488 494206 512544
rect 494058 508816 494114 508872
rect 483846 496848 483902 496904
rect 486422 496848 486478 496904
rect 487986 453872 488042 453928
rect 473358 393896 473414 393952
rect 472898 392536 472954 392592
rect 472162 389000 472218 389056
rect 474370 389000 474426 389056
rect 475842 389000 475898 389056
rect 477314 389000 477370 389056
rect 479522 389000 479578 389056
rect 494242 505164 494298 505200
rect 494242 505144 494244 505164
rect 494244 505144 494296 505164
rect 494296 505144 494298 505164
rect 494702 501200 494758 501256
rect 509514 375536 509570 375592
rect 509330 370096 509386 370152
rect 450634 349016 450690 349072
rect 409234 44784 409290 44840
rect 451738 158208 451794 158264
rect 453302 316920 453358 316976
rect 452106 155488 452162 155544
rect 452198 154128 452254 154184
rect 452106 152768 452162 152824
rect 452014 148688 452070 148744
rect 452106 140528 452162 140584
rect 452106 132404 452108 132424
rect 452108 132404 452160 132424
rect 452160 132404 452162 132424
rect 452106 132368 452162 132404
rect 452566 156884 452568 156904
rect 452568 156884 452620 156904
rect 452620 156884 452622 156904
rect 452566 156848 452622 156884
rect 452566 151444 452568 151464
rect 452568 151444 452620 151464
rect 452620 151444 452622 151464
rect 452566 151408 452622 151444
rect 452474 150048 452530 150104
rect 452566 147364 452568 147384
rect 452568 147364 452620 147384
rect 452620 147364 452622 147384
rect 452566 147328 452622 147364
rect 452566 145968 452622 146024
rect 452566 144644 452568 144664
rect 452568 144644 452620 144664
rect 452620 144644 452622 144664
rect 452566 144608 452622 144644
rect 452566 143284 452568 143304
rect 452568 143284 452620 143304
rect 452620 143284 452622 143304
rect 452566 143248 452622 143284
rect 452566 141924 452568 141944
rect 452568 141924 452620 141944
rect 452620 141924 452622 141944
rect 452566 141888 452622 141924
rect 452566 139168 452622 139224
rect 452566 137844 452568 137864
rect 452568 137844 452620 137864
rect 452620 137844 452622 137864
rect 452566 137808 452622 137844
rect 452566 136484 452568 136504
rect 452568 136484 452620 136504
rect 452620 136484 452622 136504
rect 452566 136448 452622 136484
rect 452566 135124 452568 135144
rect 452568 135124 452620 135144
rect 452620 135124 452622 135144
rect 452566 135088 452622 135124
rect 452474 133764 452476 133784
rect 452476 133764 452528 133784
rect 452528 133764 452530 133784
rect 452474 133728 452530 133764
rect 452566 131044 452568 131064
rect 452568 131044 452620 131064
rect 452620 131044 452622 131064
rect 452566 131008 452622 131044
rect 452382 129648 452438 129704
rect 452290 128288 452346 128344
rect 452198 126948 452254 126984
rect 452198 126928 452200 126948
rect 452200 126928 452252 126948
rect 452252 126928 452254 126948
rect 451922 125568 451978 125624
rect 451738 124208 451794 124264
rect 451738 122848 451794 122904
rect 451738 121488 451794 121544
rect 450726 3440 450782 3496
rect 454958 317192 455014 317248
rect 454682 316648 454738 316704
rect 456154 46552 456210 46608
rect 460202 321952 460258 322008
rect 460018 321408 460074 321464
rect 456798 262656 456854 262712
rect 456798 248784 456854 248840
rect 456798 221040 456854 221096
rect 456890 207168 456946 207224
rect 458086 234912 458142 234968
rect 458730 207168 458786 207224
rect 458914 46824 458970 46880
rect 459098 46688 459154 46744
rect 461674 321136 461730 321192
rect 462226 321816 462282 321872
rect 471610 319776 471666 319832
rect 472714 319640 472770 319696
rect 472162 319504 472218 319560
rect 482374 321272 482430 321328
rect 482926 321680 482982 321736
rect 483202 320048 483258 320104
rect 482650 319912 482706 319968
rect 483754 321544 483810 321600
rect 495806 315288 495862 315344
rect 502246 319368 502302 319424
rect 507214 322224 507270 322280
rect 509422 357584 509478 357640
rect 510710 365608 510766 365664
rect 509606 357584 509662 357640
rect 510802 355816 510858 355872
rect 509790 348336 509846 348392
rect 509698 343984 509754 344040
rect 509698 323312 509754 323368
rect 509514 322088 509570 322144
rect 509882 342352 509938 342408
rect 509790 322904 509846 322960
rect 509974 334192 510030 334248
rect 510066 331880 510122 331936
rect 510158 330248 510214 330304
rect 510894 354184 510950 354240
rect 510986 347656 511042 347712
rect 511078 346024 511134 346080
rect 511170 335688 511226 335744
rect 511998 380316 512054 380352
rect 511998 380296 512000 380316
rect 512000 380296 512052 380316
rect 512052 380296 512054 380316
rect 512734 384648 512790 384704
rect 513286 384104 513342 384160
rect 513010 383560 513066 383616
rect 512458 383036 512514 383072
rect 512458 383016 512460 383036
rect 512460 383016 512512 383036
rect 512512 383016 512514 383036
rect 512274 382472 512330 382528
rect 512458 381928 512514 381984
rect 512182 378664 512238 378720
rect 512274 378120 512330 378176
rect 512090 377576 512146 377632
rect 511998 376488 512054 376544
rect 512090 372700 512146 372736
rect 512090 372680 512092 372700
rect 512092 372680 512144 372700
rect 512144 372680 512146 372700
rect 512090 371592 512146 371648
rect 511998 367260 512054 367296
rect 511998 367240 512000 367260
rect 512000 367240 512052 367260
rect 512052 367240 512054 367260
rect 511998 364540 512054 364576
rect 511998 364520 512000 364540
rect 512000 364520 512052 364540
rect 512052 364520 512054 364540
rect 512182 368328 512238 368384
rect 511538 354728 511594 354784
rect 511906 325760 511962 325816
rect 511906 322224 511962 322280
rect 512090 363976 512146 364032
rect 512090 363432 512146 363488
rect 513286 381384 513342 381440
rect 512826 380840 512882 380896
rect 513286 379752 513342 379808
rect 513286 379208 513342 379264
rect 513194 377032 513250 377088
rect 513286 375944 513342 376000
rect 512366 374856 512422 374912
rect 512458 374312 512514 374368
rect 512642 373788 512698 373824
rect 512642 373768 512644 373788
rect 512644 373768 512696 373788
rect 512696 373768 512698 373788
rect 513286 373224 513342 373280
rect 512458 372136 512514 372192
rect 513286 371048 513342 371104
rect 512734 369980 512790 370016
rect 512734 369960 512736 369980
rect 512736 369960 512788 369980
rect 512788 369960 512790 369980
rect 513286 369416 513342 369472
rect 513470 368872 513526 368928
rect 512642 367784 512698 367840
rect 513194 366696 513250 366752
rect 513286 366152 513342 366208
rect 513286 365064 513342 365120
rect 513194 362888 513250 362944
rect 512366 362364 512422 362400
rect 512366 362344 512368 362364
rect 512368 362344 512420 362364
rect 512420 362344 512422 362364
rect 513286 361800 513342 361856
rect 512826 361256 512882 361312
rect 512366 360712 512422 360768
rect 513286 360168 513342 360224
rect 512918 359624 512974 359680
rect 512366 359080 512422 359136
rect 512458 358536 512514 358592
rect 512366 353660 512422 353696
rect 512366 353640 512368 353660
rect 512368 353640 512420 353660
rect 512420 353640 512422 353660
rect 512366 352552 512422 352608
rect 512366 350940 512422 350976
rect 512366 350920 512368 350940
rect 512368 350920 512420 350940
rect 512420 350920 512422 350940
rect 512366 349308 512422 349344
rect 512366 349288 512368 349308
rect 512368 349288 512420 349308
rect 512420 349288 512422 349308
rect 512366 345480 512422 345536
rect 512918 356360 512974 356416
rect 513286 355272 513342 355328
rect 512826 353116 512882 353152
rect 512826 353096 512828 353116
rect 512828 353096 512880 353116
rect 512880 353096 512882 353116
rect 513286 352028 513342 352064
rect 513286 352008 513288 352028
rect 513288 352008 513340 352028
rect 513340 352008 513342 352028
rect 513010 351464 513066 351520
rect 513194 350376 513250 350432
rect 513010 349832 513066 349888
rect 513010 348200 513066 348256
rect 513286 347112 513342 347168
rect 513102 346588 513158 346624
rect 513102 346568 513104 346588
rect 513104 346568 513156 346588
rect 513156 346568 513158 346588
rect 512550 344936 512606 344992
rect 512642 343848 512698 343904
rect 513010 343304 513066 343360
rect 513286 342252 513288 342272
rect 513288 342252 513340 342272
rect 513340 342252 513342 342272
rect 513286 342216 513342 342252
rect 513010 341672 513066 341728
rect 513286 341128 513342 341184
rect 513194 340584 513250 340640
rect 513102 339532 513104 339552
rect 513104 339532 513156 339552
rect 513156 339532 513158 339552
rect 513102 339496 513158 339532
rect 513286 340040 513342 340096
rect 512826 338952 512882 339008
rect 512642 338408 512698 338464
rect 513286 337864 513342 337920
rect 512642 337320 512698 337376
rect 513286 336776 513342 336832
rect 513286 336232 513342 336288
rect 512734 334600 512790 334656
rect 512918 332424 512974 332480
rect 512734 329160 512790 329216
rect 512826 325352 512882 325408
rect 513562 356904 513618 356960
rect 516966 316784 517022 316840
rect 519542 465704 519598 465760
rect 559654 699760 559710 699816
rect 580170 697176 580226 697232
rect 557538 442856 557594 442912
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580354 644000 580410 644056
rect 580170 630808 580226 630864
rect 580262 617480 580318 617536
rect 580170 590960 580226 591016
rect 579894 564304 579950 564360
rect 580170 537784 580226 537840
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580354 577632 580410 577688
rect 580446 524456 580502 524512
rect 580538 511264 580594 511320
rect 580630 458088 580686 458144
rect 580722 431568 580778 431624
rect 580814 418240 580870 418296
rect 529294 261568 529350 261624
rect 530122 226208 530178 226264
rect 529938 209208 529994 209264
rect 531318 243616 531374 243672
rect 539322 137672 539378 137728
rect 539506 135904 539562 135960
rect 539690 113192 539746 113248
rect 539598 86808 539654 86864
rect 537482 40976 537538 41032
rect 539966 108704 540022 108760
rect 540334 123120 540390 123176
rect 540242 121080 540298 121136
rect 540150 114960 540206 115016
rect 540058 104624 540114 104680
rect 539874 99184 539930 99240
rect 541070 119040 541126 119096
rect 541530 117000 541586 117056
rect 541438 110880 541494 110936
rect 541346 106800 541402 106856
rect 541254 102720 541310 102776
rect 542450 100680 542506 100736
rect 542542 96600 542598 96656
rect 541162 92520 541218 92576
rect 542726 133320 542782 133376
rect 542818 94560 542874 94616
rect 542634 90480 542690 90536
rect 543278 137808 543334 137864
rect 543186 131280 543242 131336
rect 543094 129240 543150 129296
rect 543278 127200 543334 127256
rect 543002 125160 543058 125216
rect 542910 88440 542966 88496
rect 540978 82320 541034 82376
rect 540610 48864 540666 48920
rect 539782 33632 539838 33688
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580262 258848 580318 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 578882 205672 578938 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 454682 3304 454738 3360
<< metal3 >>
rect 202781 700498 202847 700501
rect 449566 700498 449572 700500
rect 202781 700496 449572 700498
rect 202781 700440 202786 700496
rect 202842 700440 449572 700496
rect 202781 700438 449572 700440
rect 202781 700435 202847 700438
rect 449566 700436 449572 700438
rect 449636 700436 449642 700500
rect 451774 700436 451780 700500
rect 451844 700498 451850 700500
rect 478505 700498 478571 700501
rect 451844 700496 478571 700498
rect 451844 700440 478510 700496
rect 478566 700440 478571 700496
rect 451844 700438 478571 700440
rect 451844 700436 451850 700438
rect 478505 700435 478571 700438
rect 40493 700362 40559 700365
rect 447726 700362 447732 700364
rect 40493 700360 447732 700362
rect 40493 700304 40498 700360
rect 40554 700304 447732 700360
rect 40493 700302 447732 700304
rect 40493 700299 40559 700302
rect 447726 700300 447732 700302
rect 447796 700300 447802 700364
rect 455086 700300 455092 700364
rect 455156 700362 455162 700364
rect 494789 700362 494855 700365
rect 455156 700360 494855 700362
rect 455156 700304 494794 700360
rect 494850 700304 494855 700360
rect 455156 700302 494855 700304
rect 455156 700300 455162 700302
rect 494789 700299 494855 700302
rect 527173 699820 527239 699821
rect 527173 699818 527220 699820
rect 527128 699816 527220 699818
rect 527128 699760 527178 699816
rect 527128 699758 527220 699760
rect 527173 699756 527220 699758
rect 527284 699756 527290 699820
rect 556286 699756 556292 699820
rect 556356 699818 556362 699820
rect 559649 699818 559715 699821
rect 556356 699816 559715 699818
rect 556356 699760 559654 699816
rect 559710 699760 559715 699816
rect 556356 699758 559715 699760
rect 556356 699756 556362 699758
rect 527173 699755 527239 699756
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect 153193 692066 153259 692069
rect 450486 692066 450492 692068
rect 153193 692064 450492 692066
rect 153193 692008 153198 692064
rect 153254 692008 450492 692064
rect 153193 692006 450492 692008
rect 153193 692003 153259 692006
rect 450486 692004 450492 692006
rect 450556 692004 450562 692068
rect 282913 690706 282979 690709
rect 444230 690706 444236 690708
rect 282913 690704 444236 690706
rect 282913 690648 282918 690704
rect 282974 690648 444236 690704
rect 282913 690646 444236 690648
rect 282913 690643 282979 690646
rect 444230 690644 444236 690646
rect 444300 690644 444306 690708
rect 136633 689346 136699 689349
rect 450670 689346 450676 689348
rect 136633 689344 450676 689346
rect 136633 689288 136638 689344
rect 136694 689288 450676 689344
rect 136633 689286 450676 689288
rect 136633 689283 136699 689286
rect 450670 689284 450676 689286
rect 450740 689284 450746 689348
rect 22686 684524 22692 684588
rect 22756 684586 22762 684588
rect 420269 684586 420335 684589
rect 22756 684584 420335 684586
rect 22756 684528 420274 684584
rect 420330 684528 420335 684584
rect 22756 684526 420335 684528
rect 22756 684524 22762 684526
rect 420269 684523 420335 684526
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 3550 683300 3556 683364
rect 3620 683362 3626 683364
rect 445385 683362 445451 683365
rect 3620 683360 445451 683362
rect 3620 683304 445390 683360
rect 445446 683304 445451 683360
rect 3620 683302 445451 683304
rect 3620 683300 3626 683302
rect 445385 683299 445451 683302
rect 3734 683164 3740 683228
rect 3804 683226 3810 683228
rect 446857 683226 446923 683229
rect 3804 683224 446923 683226
rect 3804 683168 446862 683224
rect 446918 683168 446923 683224
rect 3804 683166 446923 683168
rect 3804 683164 3810 683166
rect 446857 683163 446923 683166
rect 3366 682756 3372 682820
rect 3436 682818 3442 682820
rect 446305 682818 446371 682821
rect 3436 682816 446371 682818
rect 3436 682760 446310 682816
rect 446366 682760 446371 682816
rect 3436 682758 446371 682760
rect 3436 682756 3442 682758
rect 446305 682755 446371 682758
rect 361757 679010 361823 679013
rect 359812 679008 361823 679010
rect 359812 678952 361762 679008
rect 361818 678952 361823 679008
rect 359812 678950 361823 678952
rect 361757 678947 361823 678950
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 3509 669898 3575 669901
rect 22686 669898 22692 669900
rect 3509 669896 22692 669898
rect 3509 669840 3514 669896
rect 3570 669840 22692 669896
rect 3509 669838 22692 669840
rect 3509 669835 3575 669838
rect 22686 669836 22692 669838
rect 22756 669836 22762 669900
rect 453246 669836 453252 669900
rect 453316 669898 453322 669900
rect 462313 669898 462379 669901
rect 453316 669896 462379 669898
rect 453316 669840 462318 669896
rect 462374 669840 462379 669896
rect 453316 669838 462379 669840
rect 453316 669836 453322 669838
rect 462313 669835 462379 669838
rect 361757 667994 361823 667997
rect 359812 667992 361823 667994
rect 359812 667936 361762 667992
rect 361818 667936 361823 667992
rect 359812 667934 361823 667936
rect 361757 667931 361823 667934
rect 457805 667994 457871 667997
rect 457805 667992 460092 667994
rect 457805 667936 457810 667992
rect 457866 667936 460092 667992
rect 457805 667934 460092 667936
rect 457805 667931 457871 667934
rect 458030 665484 458036 665548
rect 458100 665546 458106 665548
rect 458100 665486 460092 665546
rect 458100 665484 458106 665486
rect 457846 663036 457852 663100
rect 457916 663098 457922 663100
rect 457916 663038 460092 663098
rect 457916 663036 457922 663038
rect 458081 660650 458147 660653
rect 458081 660648 460092 660650
rect 458081 660592 458086 660648
rect 458142 660592 460092 660648
rect 458081 660590 460092 660592
rect 458081 660587 458147 660590
rect -960 658202 480 658292
rect 3734 658202 3740 658204
rect -960 658142 3740 658202
rect -960 658052 480 658142
rect 3734 658140 3740 658142
rect 3804 658140 3810 658204
rect 457989 658202 458055 658205
rect 457989 658200 460092 658202
rect 457989 658144 457994 658200
rect 458050 658144 460092 658200
rect 457989 658142 460092 658144
rect 457989 658139 458055 658142
rect 583520 657236 584960 657476
rect 361757 656978 361823 656981
rect 359812 656976 361823 656978
rect 359812 656920 361762 656976
rect 361818 656920 361823 656976
rect 359812 656918 361823 656920
rect 361757 656915 361823 656918
rect 459185 655754 459251 655757
rect 459185 655752 460092 655754
rect 459185 655696 459190 655752
rect 459246 655696 460092 655752
rect 459185 655694 460092 655696
rect 459185 655691 459251 655694
rect 457713 653306 457779 653309
rect 457713 653304 460092 653306
rect 457713 653248 457718 653304
rect 457774 653248 460092 653304
rect 457713 653246 460092 653248
rect 457713 653243 457779 653246
rect 457621 650858 457687 650861
rect 457621 650856 460092 650858
rect 457621 650800 457626 650856
rect 457682 650800 460092 650856
rect 457621 650798 460092 650800
rect 457621 650795 457687 650798
rect 459093 648410 459159 648413
rect 459093 648408 460092 648410
rect 459093 648352 459098 648408
rect 459154 648352 460092 648408
rect 459093 648350 460092 648352
rect 459093 648347 459159 648350
rect 361757 645962 361823 645965
rect 359812 645960 361823 645962
rect 359812 645904 361762 645960
rect 361818 645904 361823 645960
rect 359812 645902 361823 645904
rect 361757 645899 361823 645902
rect 457529 645962 457595 645965
rect 457529 645960 460092 645962
rect 457529 645904 457534 645960
rect 457590 645904 460092 645960
rect 457529 645902 460092 645904
rect 457529 645899 457595 645902
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect 459001 643514 459067 643517
rect 459001 643512 460092 643514
rect 459001 643456 459006 643512
rect 459062 643456 460092 643512
rect 459001 643454 460092 643456
rect 459001 643451 459067 643454
rect 457897 641066 457963 641069
rect 457897 641064 460092 641066
rect 457897 641008 457902 641064
rect 457958 641008 460092 641064
rect 457897 641006 460092 641008
rect 457897 641003 457963 641006
rect 458909 638618 458975 638621
rect 458909 638616 460092 638618
rect 458909 638560 458914 638616
rect 458970 638560 460092 638616
rect 458909 638558 460092 638560
rect 458909 638555 458975 638558
rect 458950 636108 458956 636172
rect 459020 636170 459026 636172
rect 459020 636110 460092 636170
rect 459020 636108 459026 636110
rect 361573 634946 361639 634949
rect 359812 634944 361639 634946
rect 359812 634888 361578 634944
rect 361634 634888 361639 634944
rect 359812 634886 361639 634888
rect 361573 634883 361639 634886
rect 459134 633660 459140 633724
rect 459204 633722 459210 633724
rect 459204 633662 460092 633722
rect 459204 633660 459210 633662
rect -960 632090 480 632180
rect 3693 632090 3759 632093
rect -960 632088 3759 632090
rect -960 632032 3698 632088
rect 3754 632032 3759 632088
rect -960 632030 3759 632032
rect -960 631940 480 632030
rect 3693 632027 3759 632030
rect 459461 631274 459527 631277
rect 459461 631272 460092 631274
rect 459461 631216 459466 631272
rect 459522 631216 460092 631272
rect 459461 631214 460092 631216
rect 459461 631211 459527 631214
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 459277 628826 459343 628829
rect 459277 628824 460092 628826
rect 459277 628768 459282 628824
rect 459338 628768 460092 628824
rect 459277 628766 460092 628768
rect 459277 628763 459343 628766
rect 459369 626378 459435 626381
rect 459369 626376 460092 626378
rect 459369 626320 459374 626376
rect 459430 626320 460092 626376
rect 459369 626318 460092 626320
rect 459369 626315 459435 626318
rect 361573 623930 361639 623933
rect 359812 623928 361639 623930
rect 359812 623872 361578 623928
rect 361634 623872 361639 623928
rect 359812 623870 361639 623872
rect 361573 623867 361639 623870
rect 459553 623862 459619 623865
rect 459553 623860 460092 623862
rect 459553 623804 459558 623860
rect 459614 623804 460092 623860
rect 459553 623802 460092 623804
rect 459553 623799 459619 623802
rect 457437 621482 457503 621485
rect 457437 621480 460092 621482
rect 457437 621424 457442 621480
rect 457498 621424 460092 621480
rect 457437 621422 460092 621424
rect 457437 621419 457503 621422
rect -960 619170 480 619260
rect 3550 619170 3556 619172
rect -960 619110 3556 619170
rect -960 619020 480 619110
rect 3550 619108 3556 619110
rect 3620 619108 3626 619172
rect 458817 619034 458883 619037
rect 458817 619032 460092 619034
rect 458817 618976 458822 619032
rect 458878 618976 460092 619032
rect 458817 618974 460092 618976
rect 458817 618971 458883 618974
rect 580257 617538 580323 617541
rect 583520 617538 584960 617628
rect 580257 617536 584960 617538
rect 580257 617480 580262 617536
rect 580318 617480 584960 617536
rect 580257 617478 584960 617480
rect 580257 617475 580323 617478
rect 583520 617388 584960 617478
rect 457345 616586 457411 616589
rect 457345 616584 460092 616586
rect 457345 616528 457350 616584
rect 457406 616528 460092 616584
rect 457345 616526 460092 616528
rect 457345 616523 457411 616526
rect 459645 614138 459711 614141
rect 459645 614136 460092 614138
rect 459645 614080 459650 614136
rect 459706 614080 460092 614136
rect 459645 614078 460092 614080
rect 459645 614075 459711 614078
rect 361573 612914 361639 612917
rect 359812 612912 361639 612914
rect 359812 612856 361578 612912
rect 361634 612856 361639 612912
rect 359812 612854 361639 612856
rect 361573 612851 361639 612854
rect 458633 611690 458699 611693
rect 458633 611688 460092 611690
rect 458633 611632 458638 611688
rect 458694 611632 460092 611688
rect 458633 611630 460092 611632
rect 458633 611627 458699 611630
rect 457253 609242 457319 609245
rect 457253 609240 460092 609242
rect 457253 609184 457258 609240
rect 457314 609184 460092 609240
rect 457253 609182 460092 609184
rect 457253 609179 457319 609182
rect 459737 606726 459803 606729
rect 459737 606724 460092 606726
rect 459737 606668 459742 606724
rect 459798 606668 460092 606724
rect 459737 606666 460092 606668
rect 459737 606663 459803 606666
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 459829 604278 459895 604281
rect 459829 604276 460092 604278
rect 459829 604220 459834 604276
rect 459890 604220 460092 604276
rect 459829 604218 460092 604220
rect 459829 604215 459895 604218
rect 583520 604060 584960 604300
rect 361573 601898 361639 601901
rect 359812 601896 361639 601898
rect 359812 601840 361578 601896
rect 361634 601840 361639 601896
rect 359812 601838 361639 601840
rect 361573 601835 361639 601838
rect 459185 601898 459251 601901
rect 459185 601896 460092 601898
rect 459185 601840 459190 601896
rect 459246 601840 460092 601896
rect 459185 601838 460092 601840
rect 459185 601835 459251 601838
rect 459093 599586 459159 599589
rect 478822 599586 478828 599588
rect 459093 599584 478828 599586
rect 459093 599528 459098 599584
rect 459154 599528 478828 599584
rect 459093 599526 478828 599528
rect 459093 599523 459159 599526
rect 478822 599524 478828 599526
rect 478892 599524 478898 599588
rect 458909 598226 458975 598229
rect 474406 598226 474412 598228
rect 458909 598224 474412 598226
rect 458909 598168 458914 598224
rect 458970 598168 474412 598224
rect 458909 598166 474412 598168
rect 458909 598163 458975 598166
rect 474406 598164 474412 598166
rect 474476 598164 474482 598228
rect 459001 597002 459067 597005
rect 474774 597002 474780 597004
rect 459001 597000 474780 597002
rect 459001 596944 459006 597000
rect 459062 596944 474780 597000
rect 459001 596942 474780 596944
rect 459001 596939 459067 596942
rect 474774 596940 474780 596942
rect 474844 596940 474850 597004
rect 458725 596866 458791 596869
rect 476430 596866 476436 596868
rect 458725 596864 476436 596866
rect 458725 596808 458730 596864
rect 458786 596808 476436 596864
rect 458725 596806 476436 596808
rect 458725 596803 458791 596806
rect 476430 596804 476436 596806
rect 476500 596804 476506 596868
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 361757 590882 361823 590885
rect 359812 590880 361823 590882
rect 359812 590824 361762 590880
rect 361818 590824 361823 590880
rect 583520 590868 584960 590958
rect 359812 590822 361823 590824
rect 361757 590819 361823 590822
rect -960 580002 480 580092
rect 3233 580002 3299 580005
rect -960 580000 3299 580002
rect -960 579944 3238 580000
rect 3294 579944 3299 580000
rect -960 579942 3299 579944
rect -960 579852 480 579942
rect 3233 579939 3299 579942
rect 361757 579866 361823 579869
rect 359812 579864 361823 579866
rect 359812 579808 361762 579864
rect 361818 579808 361823 579864
rect 359812 579806 361823 579808
rect 361757 579803 361823 579806
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect 361573 568850 361639 568853
rect 359812 568848 361639 568850
rect 359812 568792 361578 568848
rect 361634 568792 361639 568848
rect 359812 568790 361639 568792
rect 361573 568787 361639 568790
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 579889 564362 579955 564365
rect 583520 564362 584960 564452
rect 579889 564360 584960 564362
rect 579889 564304 579894 564360
rect 579950 564304 584960 564360
rect 579889 564302 584960 564304
rect 579889 564299 579955 564302
rect 583520 564212 584960 564302
rect 361573 557834 361639 557837
rect 359812 557832 361639 557834
rect 359812 557776 361578 557832
rect 361634 557776 361639 557832
rect 359812 557774 361639 557776
rect 361573 557771 361639 557774
rect -960 553890 480 553980
rect 4061 553890 4127 553893
rect -960 553888 4127 553890
rect -960 553832 4066 553888
rect 4122 553832 4127 553888
rect -960 553830 4127 553832
rect -960 553740 480 553830
rect 4061 553827 4127 553830
rect 583520 551020 584960 551260
rect 361757 546818 361823 546821
rect 359812 546816 361823 546818
rect 359812 546760 361762 546816
rect 361818 546760 361823 546816
rect 359812 546758 361823 546760
rect 361757 546755 361823 546758
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 361757 535802 361823 535805
rect 359812 535800 361823 535802
rect 359812 535744 361762 535800
rect 361818 535744 361823 535800
rect 359812 535742 361823 535744
rect 361757 535739 361823 535742
rect -960 527914 480 528004
rect 3969 527914 4035 527917
rect -960 527912 4035 527914
rect -960 527856 3974 527912
rect 4030 527856 4035 527912
rect -960 527854 4035 527856
rect -960 527764 480 527854
rect 3969 527851 4035 527854
rect 361757 524786 361823 524789
rect 359812 524784 361823 524786
rect 359812 524728 361762 524784
rect 361818 524728 361823 524784
rect 359812 524726 361823 524728
rect 361757 524723 361823 524726
rect 580441 524514 580507 524517
rect 583520 524514 584960 524604
rect 580441 524512 584960 524514
rect 580441 524456 580446 524512
rect 580502 524456 584960 524512
rect 580441 524454 584960 524456
rect 580441 524451 580507 524454
rect 583520 524364 584960 524454
rect 459461 522338 459527 522341
rect 472014 522338 472020 522340
rect 459461 522336 472020 522338
rect 459461 522280 459466 522336
rect 459522 522280 472020 522336
rect 459461 522278 472020 522280
rect 459461 522275 459527 522278
rect 472014 522276 472020 522278
rect 472084 522276 472090 522340
rect 457846 519420 457852 519484
rect 457916 519482 457922 519484
rect 467189 519482 467255 519485
rect 457916 519480 467255 519482
rect 457916 519424 467194 519480
rect 467250 519424 467255 519480
rect 457916 519422 467255 519424
rect 457916 519420 457922 519422
rect 467189 519419 467255 519422
rect 458030 517516 458036 517580
rect 458100 517578 458106 517580
rect 462957 517578 463023 517581
rect 458100 517576 463023 517578
rect 458100 517520 462962 517576
rect 463018 517520 463023 517576
rect 458100 517518 463023 517520
rect 458100 517516 458106 517518
rect 462957 517515 463023 517518
rect 448145 516762 448211 516765
rect 494145 516762 494211 516765
rect 494329 516762 494395 516765
rect 448145 516760 494395 516762
rect 448145 516704 448150 516760
rect 448206 516704 494150 516760
rect 494206 516704 494334 516760
rect 494390 516704 494395 516760
rect 448145 516702 494395 516704
rect 448145 516699 448211 516702
rect 494145 516699 494211 516702
rect 494329 516699 494395 516702
rect 450126 516354 450186 516528
rect 450629 516354 450695 516357
rect 450126 516352 450695 516354
rect 450126 516296 450634 516352
rect 450690 516296 450695 516352
rect 450126 516294 450695 516296
rect 448278 516156 448284 516220
rect 448348 516218 448354 516220
rect 450126 516218 450186 516294
rect 450629 516291 450695 516294
rect 448348 516158 450186 516218
rect 491845 516218 491911 516221
rect 491845 516216 491954 516218
rect 491845 516160 491850 516216
rect 491906 516160 491954 516216
rect 448348 516156 448354 516158
rect 491845 516155 491954 516160
rect 491894 515946 491954 516155
rect 494145 515946 494211 515949
rect 491894 515944 494211 515946
rect 491894 515888 494150 515944
rect 494206 515888 494211 515944
rect 491894 515886 494211 515888
rect 494145 515883 494211 515886
rect -960 514858 480 514948
rect 3877 514858 3943 514861
rect -960 514856 3943 514858
rect -960 514800 3882 514856
rect 3938 514800 3943 514856
rect -960 514798 3943 514800
rect -960 514708 480 514798
rect 3877 514795 3943 514798
rect 447961 514450 448027 514453
rect 448513 514450 448579 514453
rect 447961 514448 450186 514450
rect 447961 514392 447966 514448
rect 448022 514392 448518 514448
rect 448574 514392 450186 514448
rect 447961 514390 450186 514392
rect 447961 514387 448027 514390
rect 448513 514387 448579 514390
rect 450126 514352 450186 514390
rect 361757 513770 361823 513773
rect 359812 513768 361823 513770
rect 359812 513712 361762 513768
rect 361818 513712 361823 513768
rect 359812 513710 361823 513712
rect 361757 513707 361823 513710
rect 447409 512818 447475 512821
rect 448329 512818 448395 512821
rect 447409 512816 450186 512818
rect 447409 512760 447414 512816
rect 447470 512760 448334 512816
rect 448390 512760 450186 512816
rect 447409 512758 450186 512760
rect 447409 512755 447475 512758
rect 448329 512755 448395 512758
rect 450126 512176 450186 512758
rect 494145 512546 494211 512549
rect 491894 512544 494211 512546
rect 491894 512488 494150 512544
rect 494206 512488 494211 512544
rect 491894 512486 494211 512488
rect 491894 512448 491954 512486
rect 494145 512483 494211 512486
rect 580533 511322 580599 511325
rect 583520 511322 584960 511412
rect 580533 511320 584960 511322
rect 580533 511264 580538 511320
rect 580594 511264 584960 511320
rect 580533 511262 584960 511264
rect 580533 511259 580599 511262
rect 583520 511172 584960 511262
rect 448421 510506 448487 510509
rect 448421 510504 450186 510506
rect 448421 510448 448426 510504
rect 448482 510448 450186 510504
rect 448421 510446 450186 510448
rect 448421 510443 448487 510446
rect 450126 510000 450186 510446
rect 491894 508874 491954 508912
rect 494053 508874 494119 508877
rect 491894 508872 494119 508874
rect 491894 508816 494058 508872
rect 494114 508816 494119 508872
rect 491894 508814 494119 508816
rect 494053 508811 494119 508814
rect 448145 507786 448211 507789
rect 450126 507786 450186 507824
rect 448145 507784 450186 507786
rect 448145 507728 448150 507784
rect 448206 507728 450186 507784
rect 448145 507726 450186 507728
rect 448145 507723 448211 507726
rect 447961 505202 448027 505205
rect 450126 505202 450186 505648
rect 447961 505200 450186 505202
rect 447961 505144 447966 505200
rect 448022 505144 450186 505200
rect 447961 505142 450186 505144
rect 491894 505202 491954 505376
rect 494237 505202 494303 505205
rect 491894 505200 494303 505202
rect 491894 505144 494242 505200
rect 494298 505144 494303 505200
rect 491894 505142 494303 505144
rect 447961 505139 448027 505142
rect 494237 505139 494303 505142
rect 448329 503434 448395 503437
rect 449801 503434 449867 503437
rect 450126 503434 450186 503472
rect 448329 503432 450186 503434
rect 448329 503376 448334 503432
rect 448390 503376 449806 503432
rect 449862 503376 450186 503432
rect 448329 503374 450186 503376
rect 448329 503371 448395 503374
rect 449801 503371 449867 503374
rect 361757 502754 361823 502757
rect 359812 502752 361823 502754
rect 359812 502696 361762 502752
rect 361818 502696 361823 502752
rect 359812 502694 361823 502696
rect 361757 502691 361823 502694
rect 448053 501938 448119 501941
rect 448053 501936 450186 501938
rect -960 501802 480 501892
rect 448053 501880 448058 501936
rect 448114 501880 450186 501936
rect 448053 501878 450186 501880
rect 448053 501875 448119 501878
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 450126 500986 450186 501878
rect 491894 501258 491954 501840
rect 494697 501258 494763 501261
rect 489870 501256 494763 501258
rect 489870 501200 494702 501256
rect 494758 501200 494763 501256
rect 489870 501198 494763 501200
rect 489870 501122 489930 501198
rect 494697 501195 494763 501198
rect 470550 501062 489930 501122
rect 470550 500986 470610 501062
rect 450126 500926 470610 500986
rect 583520 497844 584960 498084
rect 483054 496844 483060 496908
rect 483124 496906 483130 496908
rect 483841 496906 483907 496909
rect 486417 496908 486483 496909
rect 486366 496906 486372 496908
rect 483124 496904 483907 496906
rect 483124 496848 483846 496904
rect 483902 496848 483907 496904
rect 483124 496846 483907 496848
rect 486326 496846 486372 496906
rect 486436 496904 486483 496908
rect 486478 496848 486483 496904
rect 483124 496844 483130 496846
rect 483841 496843 483907 496846
rect 486366 496844 486372 496846
rect 486436 496844 486483 496848
rect 486417 496843 486483 496844
rect 448278 496028 448284 496092
rect 448348 496090 448354 496092
rect 449893 496090 449959 496093
rect 448348 496088 449959 496090
rect 448348 496032 449898 496088
rect 449954 496032 449959 496088
rect 448348 496030 449959 496032
rect 448348 496028 448354 496030
rect 449893 496027 449959 496030
rect 361757 491738 361823 491741
rect 359812 491736 361823 491738
rect 359812 491680 361762 491736
rect 361818 491680 361823 491736
rect 359812 491678 361823 491680
rect 361757 491675 361823 491678
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 361757 480722 361823 480725
rect 359812 480720 361823 480722
rect 359812 480664 361762 480720
rect 361818 480664 361823 480720
rect 359812 480662 361823 480664
rect 361757 480659 361823 480662
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 361757 469706 361823 469709
rect 359812 469704 361823 469706
rect 359812 469648 361762 469704
rect 361818 469648 361823 469704
rect 359812 469646 361823 469648
rect 361757 469643 361823 469646
rect 519537 465762 519603 465765
rect 527214 465762 527220 465764
rect 519537 465760 527220 465762
rect 519537 465704 519542 465760
rect 519598 465704 527220 465760
rect 519537 465702 527220 465704
rect 519537 465699 519603 465702
rect 527214 465700 527220 465702
rect 527284 465700 527290 465764
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 361757 458690 361823 458693
rect 359812 458688 361823 458690
rect 359812 458632 361762 458688
rect 361818 458632 361823 458688
rect 359812 458630 361823 458632
rect 361757 458627 361823 458630
rect 580625 458146 580691 458149
rect 583520 458146 584960 458236
rect 580625 458144 584960 458146
rect 580625 458088 580630 458144
rect 580686 458088 584960 458144
rect 580625 458086 584960 458088
rect 580625 458083 580691 458086
rect 583520 457996 584960 458086
rect 487102 453868 487108 453932
rect 487172 453930 487178 453932
rect 487981 453930 488047 453933
rect 487172 453928 488047 453930
rect 487172 453872 487986 453928
rect 488042 453872 488047 453928
rect 487172 453870 488047 453872
rect 487172 453868 487178 453870
rect 487981 453867 488047 453870
rect -960 449578 480 449668
rect 3509 449578 3575 449581
rect -960 449576 3575 449578
rect -960 449520 3514 449576
rect 3570 449520 3575 449576
rect -960 449518 3575 449520
rect -960 449428 480 449518
rect 3509 449515 3575 449518
rect 361573 447674 361639 447677
rect 359812 447672 361639 447674
rect 359812 447616 361578 447672
rect 361634 447616 361639 447672
rect 359812 447614 361639 447616
rect 361573 447611 361639 447614
rect 583520 444668 584960 444908
rect 557533 442914 557599 442917
rect 555956 442912 557599 442914
rect 555956 442856 557538 442912
rect 557594 442856 557599 442912
rect 555956 442854 557599 442856
rect 557533 442851 557599 442854
rect -960 436508 480 436748
rect 362217 436658 362283 436661
rect 359812 436656 362283 436658
rect 359812 436600 362222 436656
rect 362278 436600 362283 436656
rect 359812 436598 362283 436600
rect 362217 436595 362283 436598
rect 580717 431626 580783 431629
rect 583520 431626 584960 431716
rect 580717 431624 584960 431626
rect 580717 431568 580722 431624
rect 580778 431568 584960 431624
rect 580717 431566 584960 431568
rect 580717 431563 580783 431566
rect 583520 431476 584960 431566
rect 362309 425642 362375 425645
rect 359812 425640 362375 425642
rect 359812 425584 362314 425640
rect 362370 425584 362375 425640
rect 359812 425582 362375 425584
rect 362309 425579 362375 425582
rect -960 423602 480 423692
rect 3693 423602 3759 423605
rect -960 423600 3759 423602
rect -960 423544 3698 423600
rect 3754 423544 3759 423600
rect -960 423542 3759 423544
rect -960 423452 480 423542
rect 3693 423539 3759 423542
rect 444189 422922 444255 422925
rect 455086 422922 455092 422924
rect 444189 422920 455092 422922
rect 444189 422864 444194 422920
rect 444250 422864 455092 422920
rect 444189 422862 455092 422864
rect 444189 422859 444255 422862
rect 455086 422860 455092 422862
rect 455156 422860 455162 422924
rect 444046 421908 444052 421972
rect 444116 421970 444122 421972
rect 444281 421970 444347 421973
rect 444116 421968 444347 421970
rect 444116 421912 444286 421968
rect 444342 421912 444347 421968
rect 444116 421910 444347 421912
rect 444116 421908 444122 421910
rect 444281 421907 444347 421910
rect 442901 420202 442967 420205
rect 451774 420202 451780 420204
rect 442901 420200 451780 420202
rect 442901 420144 442906 420200
rect 442962 420144 451780 420200
rect 442901 420142 451780 420144
rect 442901 420139 442967 420142
rect 451774 420140 451780 420142
rect 451844 420140 451850 420204
rect 580809 418298 580875 418301
rect 583520 418298 584960 418388
rect 580809 418296 584960 418298
rect 580809 418240 580814 418296
rect 580870 418240 584960 418296
rect 580809 418238 584960 418240
rect 580809 418235 580875 418238
rect 583520 418148 584960 418238
rect 361573 414626 361639 414629
rect 359812 414624 361639 414626
rect 359812 414568 361578 414624
rect 361634 414568 361639 414624
rect 359812 414566 361639 414568
rect 361573 414563 361639 414566
rect -960 410546 480 410636
rect 3969 410546 4035 410549
rect -960 410544 4035 410546
rect -960 410488 3974 410544
rect 4030 410488 4035 410544
rect -960 410486 4035 410488
rect -960 410396 480 410486
rect 3969 410483 4035 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 361573 403610 361639 403613
rect 359812 403608 361639 403610
rect 359812 403552 361578 403608
rect 361634 403552 361639 403608
rect 359812 403550 361639 403552
rect 361573 403547 361639 403550
rect -960 397490 480 397580
rect 3785 397490 3851 397493
rect -960 397488 3851 397490
rect -960 397432 3790 397488
rect 3846 397432 3851 397488
rect -960 397430 3851 397432
rect -960 397340 480 397430
rect 3785 397427 3851 397430
rect 458950 393892 458956 393956
rect 459020 393954 459026 393956
rect 473353 393954 473419 393957
rect 459020 393952 473419 393954
rect 459020 393896 473358 393952
rect 473414 393896 473419 393952
rect 459020 393894 473419 393896
rect 459020 393892 459026 393894
rect 473353 393891 473419 393894
rect 361573 392594 361639 392597
rect 359812 392592 361639 392594
rect 359812 392536 361578 392592
rect 361634 392536 361639 392592
rect 359812 392534 361639 392536
rect 361573 392531 361639 392534
rect 459134 392532 459140 392596
rect 459204 392594 459210 392596
rect 472893 392594 472959 392597
rect 459204 392592 472959 392594
rect 459204 392536 472898 392592
rect 472954 392536 472959 392592
rect 459204 392534 472959 392536
rect 459204 392532 459210 392534
rect 472893 392531 472959 392534
rect 583520 391628 584960 391868
rect 472014 388996 472020 389060
rect 472084 389058 472090 389060
rect 472157 389058 472223 389061
rect 474365 389060 474431 389061
rect 474365 389058 474412 389060
rect 472084 389056 472223 389058
rect 472084 389000 472162 389056
rect 472218 389000 472223 389056
rect 472084 388998 472223 389000
rect 474320 389056 474412 389058
rect 474320 389000 474370 389056
rect 474320 388998 474412 389000
rect 472084 388996 472090 388998
rect 472157 388995 472223 388998
rect 474365 388996 474412 388998
rect 474476 388996 474482 389060
rect 474774 388996 474780 389060
rect 474844 389058 474850 389060
rect 475837 389058 475903 389061
rect 474844 389056 475903 389058
rect 474844 389000 475842 389056
rect 475898 389000 475903 389056
rect 474844 388998 475903 389000
rect 474844 388996 474850 388998
rect 474365 388995 474431 388996
rect 475837 388995 475903 388998
rect 476430 388996 476436 389060
rect 476500 389058 476506 389060
rect 477309 389058 477375 389061
rect 476500 389056 477375 389058
rect 476500 389000 477314 389056
rect 477370 389000 477375 389056
rect 476500 388998 477375 389000
rect 476500 388996 476506 388998
rect 477309 388995 477375 388998
rect 478822 388996 478828 389060
rect 478892 389058 478898 389060
rect 479517 389058 479583 389061
rect 478892 389056 479583 389058
rect 478892 389000 479522 389056
rect 479578 389000 479583 389056
rect 478892 388998 479583 389000
rect 478892 388996 478898 388998
rect 479517 388995 479583 388998
rect 445661 387698 445727 387701
rect 453246 387698 453252 387700
rect 445661 387696 453252 387698
rect 445661 387640 445666 387696
rect 445722 387640 453252 387696
rect 445661 387638 453252 387640
rect 445661 387635 445727 387638
rect 453246 387636 453252 387638
rect 453316 387636 453322 387700
rect 449433 387154 449499 387157
rect 483054 387154 483060 387156
rect 449433 387152 483060 387154
rect 449433 387096 449438 387152
rect 449494 387096 483060 387152
rect 449433 387094 483060 387096
rect 449433 387091 449499 387094
rect 483054 387092 483060 387094
rect 483124 387092 483130 387156
rect 449065 387018 449131 387021
rect 486366 387018 486372 387020
rect 449065 387016 486372 387018
rect 449065 386960 449070 387016
rect 449126 386960 486372 387016
rect 449065 386958 486372 386960
rect 449065 386955 449131 386958
rect 486366 386956 486372 386958
rect 486436 386956 486442 387020
rect 449525 385658 449591 385661
rect 487102 385658 487108 385660
rect 449525 385656 487108 385658
rect 449525 385600 449530 385656
rect 449586 385600 487108 385656
rect 449525 385598 487108 385600
rect 449525 385595 449591 385598
rect 487102 385596 487108 385598
rect 487172 385596 487178 385660
rect 512729 384706 512795 384709
rect 509956 384704 512795 384706
rect 509956 384648 512734 384704
rect 512790 384648 512795 384704
rect 509956 384646 512795 384648
rect 512729 384643 512795 384646
rect -960 384284 480 384524
rect 513281 384162 513347 384165
rect 509956 384160 513347 384162
rect 509956 384104 513286 384160
rect 513342 384104 513347 384160
rect 509956 384102 513347 384104
rect 513281 384099 513347 384102
rect 447133 383618 447199 383621
rect 513005 383618 513071 383621
rect 447133 383616 450156 383618
rect 447133 383560 447138 383616
rect 447194 383560 450156 383616
rect 447133 383558 450156 383560
rect 509956 383616 513071 383618
rect 509956 383560 513010 383616
rect 513066 383560 513071 383616
rect 509956 383558 513071 383560
rect 447133 383555 447199 383558
rect 513005 383555 513071 383558
rect 512453 383074 512519 383077
rect 509956 383072 512519 383074
rect 509956 383016 512458 383072
rect 512514 383016 512519 383072
rect 509956 383014 512519 383016
rect 512453 383011 512519 383014
rect 447317 382938 447383 382941
rect 447317 382936 450156 382938
rect 447317 382880 447322 382936
rect 447378 382880 450156 382936
rect 447317 382878 450156 382880
rect 447317 382875 447383 382878
rect 512269 382530 512335 382533
rect 509956 382528 512335 382530
rect 509956 382472 512274 382528
rect 512330 382472 512335 382528
rect 509956 382470 512335 382472
rect 512269 382467 512335 382470
rect 447133 382258 447199 382261
rect 447133 382256 450156 382258
rect 447133 382200 447138 382256
rect 447194 382200 450156 382256
rect 447133 382198 450156 382200
rect 447133 382195 447199 382198
rect 512453 381986 512519 381989
rect 509956 381984 512519 381986
rect 509956 381928 512458 381984
rect 512514 381928 512519 381984
rect 509956 381926 512519 381928
rect 512453 381923 512519 381926
rect 361573 381578 361639 381581
rect 359812 381576 361639 381578
rect 359812 381520 361578 381576
rect 361634 381520 361639 381576
rect 359812 381518 361639 381520
rect 361573 381515 361639 381518
rect 447317 381578 447383 381581
rect 447317 381576 450156 381578
rect 447317 381520 447322 381576
rect 447378 381520 450156 381576
rect 447317 381518 450156 381520
rect 447317 381515 447383 381518
rect 513281 381442 513347 381445
rect 509956 381440 513347 381442
rect 509956 381384 513286 381440
rect 513342 381384 513347 381440
rect 509956 381382 513347 381384
rect 513281 381379 513347 381382
rect 447133 380898 447199 380901
rect 512821 380898 512887 380901
rect 447133 380896 450156 380898
rect 447133 380840 447138 380896
rect 447194 380840 450156 380896
rect 447133 380838 450156 380840
rect 509956 380896 512887 380898
rect 509956 380840 512826 380896
rect 512882 380840 512887 380896
rect 509956 380838 512887 380840
rect 447133 380835 447199 380838
rect 512821 380835 512887 380838
rect 511993 380354 512059 380357
rect 509956 380352 512059 380354
rect 509956 380296 511998 380352
rect 512054 380296 512059 380352
rect 509956 380294 512059 380296
rect 511993 380291 512059 380294
rect 447501 380218 447567 380221
rect 447501 380216 450156 380218
rect 447501 380160 447506 380216
rect 447562 380160 450156 380216
rect 447501 380158 450156 380160
rect 447501 380155 447567 380158
rect 513281 379810 513347 379813
rect 509956 379808 513347 379810
rect 509956 379752 513286 379808
rect 513342 379752 513347 379808
rect 509956 379750 513347 379752
rect 513281 379747 513347 379750
rect 447317 379538 447383 379541
rect 447317 379536 450156 379538
rect 447317 379480 447322 379536
rect 447378 379480 450156 379536
rect 447317 379478 450156 379480
rect 447317 379475 447383 379478
rect 513281 379266 513347 379269
rect 509956 379264 513347 379266
rect 509956 379208 513286 379264
rect 513342 379208 513347 379264
rect 509956 379206 513347 379208
rect 513281 379203 513347 379206
rect 447133 378858 447199 378861
rect 447133 378856 450156 378858
rect 447133 378800 447138 378856
rect 447194 378800 450156 378856
rect 447133 378798 450156 378800
rect 447133 378795 447199 378798
rect 512177 378722 512243 378725
rect 509956 378720 512243 378722
rect 509956 378664 512182 378720
rect 512238 378664 512243 378720
rect 509956 378662 512243 378664
rect 512177 378659 512243 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 447501 378178 447567 378181
rect 512269 378178 512335 378181
rect 447501 378176 450156 378178
rect 447501 378120 447506 378176
rect 447562 378120 450156 378176
rect 447501 378118 450156 378120
rect 509956 378176 512335 378178
rect 509956 378120 512274 378176
rect 512330 378120 512335 378176
rect 509956 378118 512335 378120
rect 447501 378115 447567 378118
rect 512269 378115 512335 378118
rect 512085 377634 512151 377637
rect 509956 377632 512151 377634
rect 509956 377576 512090 377632
rect 512146 377576 512151 377632
rect 509956 377574 512151 377576
rect 512085 377571 512151 377574
rect 447133 377498 447199 377501
rect 447133 377496 450156 377498
rect 447133 377440 447138 377496
rect 447194 377440 450156 377496
rect 447133 377438 450156 377440
rect 447133 377435 447199 377438
rect 513189 377090 513255 377093
rect 509956 377088 513255 377090
rect 509956 377032 513194 377088
rect 513250 377032 513255 377088
rect 509956 377030 513255 377032
rect 513189 377027 513255 377030
rect 447317 376818 447383 376821
rect 447317 376816 450156 376818
rect 447317 376760 447322 376816
rect 447378 376760 450156 376816
rect 447317 376758 450156 376760
rect 447317 376755 447383 376758
rect 511993 376546 512059 376549
rect 509956 376544 512059 376546
rect 509956 376488 511998 376544
rect 512054 376488 512059 376544
rect 509956 376486 512059 376488
rect 511993 376483 512059 376486
rect 447133 376138 447199 376141
rect 447133 376136 450156 376138
rect 447133 376080 447138 376136
rect 447194 376080 450156 376136
rect 447133 376078 450156 376080
rect 447133 376075 447199 376078
rect 513281 376002 513347 376005
rect 509956 376000 513347 376002
rect 509956 375944 513286 376000
rect 513342 375944 513347 376000
rect 509956 375942 513347 375944
rect 513281 375939 513347 375942
rect 509509 375594 509575 375597
rect 509509 375592 509618 375594
rect 509509 375536 509514 375592
rect 509570 375536 509618 375592
rect 509509 375531 509618 375536
rect 447317 375458 447383 375461
rect 447317 375456 450156 375458
rect 447317 375400 447322 375456
rect 447378 375400 450156 375456
rect 509558 375428 509618 375531
rect 447317 375398 450156 375400
rect 447317 375395 447383 375398
rect 512361 374914 512427 374917
rect 509956 374912 512427 374914
rect 509956 374856 512366 374912
rect 512422 374856 512427 374912
rect 509956 374854 512427 374856
rect 512361 374851 512427 374854
rect 447133 374778 447199 374781
rect 447133 374776 450156 374778
rect 447133 374720 447138 374776
rect 447194 374720 450156 374776
rect 447133 374718 450156 374720
rect 447133 374715 447199 374718
rect 512453 374370 512519 374373
rect 509956 374368 512519 374370
rect 509956 374312 512458 374368
rect 512514 374312 512519 374368
rect 509956 374310 512519 374312
rect 512453 374307 512519 374310
rect 447317 374098 447383 374101
rect 447317 374096 450156 374098
rect 447317 374040 447322 374096
rect 447378 374040 450156 374096
rect 447317 374038 450156 374040
rect 447317 374035 447383 374038
rect 512637 373826 512703 373829
rect 509956 373824 512703 373826
rect 509956 373768 512642 373824
rect 512698 373768 512703 373824
rect 509956 373766 512703 373768
rect 512637 373763 512703 373766
rect 447133 373418 447199 373421
rect 447133 373416 450156 373418
rect 447133 373360 447138 373416
rect 447194 373360 450156 373416
rect 447133 373358 450156 373360
rect 447133 373355 447199 373358
rect 513281 373282 513347 373285
rect 509956 373280 513347 373282
rect 509956 373224 513286 373280
rect 513342 373224 513347 373280
rect 509956 373222 513347 373224
rect 513281 373219 513347 373222
rect 447317 372738 447383 372741
rect 512085 372738 512151 372741
rect 447317 372736 450156 372738
rect 447317 372680 447322 372736
rect 447378 372680 450156 372736
rect 447317 372678 450156 372680
rect 509956 372736 512151 372738
rect 509956 372680 512090 372736
rect 512146 372680 512151 372736
rect 509956 372678 512151 372680
rect 447317 372675 447383 372678
rect 512085 372675 512151 372678
rect 512453 372194 512519 372197
rect 509956 372192 512519 372194
rect 509956 372136 512458 372192
rect 512514 372136 512519 372192
rect 509956 372134 512519 372136
rect 512453 372131 512519 372134
rect 447133 372058 447199 372061
rect 447133 372056 450156 372058
rect 447133 372000 447138 372056
rect 447194 372000 450156 372056
rect 447133 371998 450156 372000
rect 447133 371995 447199 371998
rect 512085 371650 512151 371653
rect 509956 371648 512151 371650
rect 509956 371592 512090 371648
rect 512146 371592 512151 371648
rect 509956 371590 512151 371592
rect 512085 371587 512151 371590
rect -960 371378 480 371468
rect 3969 371378 4035 371381
rect -960 371376 4035 371378
rect -960 371320 3974 371376
rect 4030 371320 4035 371376
rect -960 371318 4035 371320
rect -960 371228 480 371318
rect 3969 371315 4035 371318
rect 447317 371378 447383 371381
rect 447317 371376 450156 371378
rect 447317 371320 447322 371376
rect 447378 371320 450156 371376
rect 447317 371318 450156 371320
rect 447317 371315 447383 371318
rect 513281 371106 513347 371109
rect 509956 371104 513347 371106
rect 509956 371048 513286 371104
rect 513342 371048 513347 371104
rect 509956 371046 513347 371048
rect 513281 371043 513347 371046
rect 447133 370698 447199 370701
rect 447133 370696 450156 370698
rect 447133 370640 447138 370696
rect 447194 370640 450156 370696
rect 447133 370638 450156 370640
rect 447133 370635 447199 370638
rect 361573 370562 361639 370565
rect 359812 370560 361639 370562
rect 359812 370504 361578 370560
rect 361634 370504 361639 370560
rect 359812 370502 361639 370504
rect 361573 370499 361639 370502
rect 509374 370157 509434 370532
rect 509325 370152 509434 370157
rect 509325 370096 509330 370152
rect 509386 370096 509434 370152
rect 509325 370094 509434 370096
rect 509325 370091 509391 370094
rect 447317 370018 447383 370021
rect 512729 370018 512795 370021
rect 447317 370016 450156 370018
rect 447317 369960 447322 370016
rect 447378 369960 450156 370016
rect 447317 369958 450156 369960
rect 509956 370016 512795 370018
rect 509956 369960 512734 370016
rect 512790 369960 512795 370016
rect 509956 369958 512795 369960
rect 447317 369955 447383 369958
rect 512729 369955 512795 369958
rect 513281 369474 513347 369477
rect 509956 369472 513347 369474
rect 509956 369416 513286 369472
rect 513342 369416 513347 369472
rect 509956 369414 513347 369416
rect 513281 369411 513347 369414
rect 447133 369338 447199 369341
rect 447133 369336 450156 369338
rect 447133 369280 447138 369336
rect 447194 369280 450156 369336
rect 447133 369278 450156 369280
rect 447133 369275 447199 369278
rect 513465 368930 513531 368933
rect 509956 368928 513531 368930
rect 509956 368872 513470 368928
rect 513526 368872 513531 368928
rect 509956 368870 513531 368872
rect 513465 368867 513531 368870
rect 447317 368658 447383 368661
rect 447317 368656 450156 368658
rect 447317 368600 447322 368656
rect 447378 368600 450156 368656
rect 447317 368598 450156 368600
rect 447317 368595 447383 368598
rect 512177 368386 512243 368389
rect 509956 368384 512243 368386
rect 509956 368328 512182 368384
rect 512238 368328 512243 368384
rect 509956 368326 512243 368328
rect 512177 368323 512243 368326
rect 447133 367978 447199 367981
rect 447133 367976 450156 367978
rect 447133 367920 447138 367976
rect 447194 367920 450156 367976
rect 447133 367918 450156 367920
rect 447133 367915 447199 367918
rect 512637 367842 512703 367845
rect 509956 367840 512703 367842
rect 509956 367784 512642 367840
rect 512698 367784 512703 367840
rect 509956 367782 512703 367784
rect 512637 367779 512703 367782
rect 447317 367298 447383 367301
rect 511993 367298 512059 367301
rect 447317 367296 450156 367298
rect 447317 367240 447322 367296
rect 447378 367240 450156 367296
rect 447317 367238 450156 367240
rect 509956 367296 512059 367298
rect 509956 367240 511998 367296
rect 512054 367240 512059 367296
rect 509956 367238 512059 367240
rect 447317 367235 447383 367238
rect 511993 367235 512059 367238
rect 513189 366754 513255 366757
rect 509956 366752 513255 366754
rect 509956 366696 513194 366752
rect 513250 366696 513255 366752
rect 509956 366694 513255 366696
rect 513189 366691 513255 366694
rect 447317 366618 447383 366621
rect 447317 366616 450156 366618
rect 447317 366560 447322 366616
rect 447378 366560 450156 366616
rect 447317 366558 450156 366560
rect 447317 366555 447383 366558
rect 513281 366210 513347 366213
rect 509956 366208 513347 366210
rect 509956 366152 513286 366208
rect 513342 366152 513347 366208
rect 509956 366150 513347 366152
rect 513281 366147 513347 366150
rect 447133 365938 447199 365941
rect 447133 365936 450156 365938
rect 447133 365880 447138 365936
rect 447194 365880 450156 365936
rect 447133 365878 450156 365880
rect 447133 365875 447199 365878
rect 510705 365666 510771 365669
rect 509956 365664 510771 365666
rect 509956 365608 510710 365664
rect 510766 365608 510771 365664
rect 509956 365606 510771 365608
rect 510705 365603 510771 365606
rect 447317 365258 447383 365261
rect 447317 365256 450156 365258
rect 447317 365200 447322 365256
rect 447378 365200 450156 365256
rect 447317 365198 450156 365200
rect 447317 365195 447383 365198
rect 513281 365122 513347 365125
rect 509956 365120 513347 365122
rect 509956 365064 513286 365120
rect 513342 365064 513347 365120
rect 509956 365062 513347 365064
rect 513281 365059 513347 365062
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 447133 364578 447199 364581
rect 511993 364578 512059 364581
rect 447133 364576 450156 364578
rect 447133 364520 447138 364576
rect 447194 364520 450156 364576
rect 447133 364518 450156 364520
rect 509956 364576 512059 364578
rect 509956 364520 511998 364576
rect 512054 364520 512059 364576
rect 509956 364518 512059 364520
rect 447133 364515 447199 364518
rect 511993 364515 512059 364518
rect 512085 364034 512151 364037
rect 509956 364032 512151 364034
rect 509956 363976 512090 364032
rect 512146 363976 512151 364032
rect 509956 363974 512151 363976
rect 512085 363971 512151 363974
rect 447317 363898 447383 363901
rect 447317 363896 450156 363898
rect 447317 363840 447322 363896
rect 447378 363840 450156 363896
rect 447317 363838 450156 363840
rect 447317 363835 447383 363838
rect 512085 363490 512151 363493
rect 509956 363488 512151 363490
rect 509956 363432 512090 363488
rect 512146 363432 512151 363488
rect 509956 363430 512151 363432
rect 512085 363427 512151 363430
rect 447133 363218 447199 363221
rect 447133 363216 450156 363218
rect 447133 363160 447138 363216
rect 447194 363160 450156 363216
rect 447133 363158 450156 363160
rect 447133 363155 447199 363158
rect 513189 362946 513255 362949
rect 509956 362944 513255 362946
rect 509956 362888 513194 362944
rect 513250 362888 513255 362944
rect 509956 362886 513255 362888
rect 513189 362883 513255 362886
rect 447317 362538 447383 362541
rect 447317 362536 450156 362538
rect 447317 362480 447322 362536
rect 447378 362480 450156 362536
rect 447317 362478 450156 362480
rect 447317 362475 447383 362478
rect 512361 362402 512427 362405
rect 509956 362400 512427 362402
rect 509956 362344 512366 362400
rect 512422 362344 512427 362400
rect 509956 362342 512427 362344
rect 512361 362339 512427 362342
rect 447133 361858 447199 361861
rect 513281 361858 513347 361861
rect 447133 361856 450156 361858
rect 447133 361800 447138 361856
rect 447194 361800 450156 361856
rect 447133 361798 450156 361800
rect 509956 361856 513347 361858
rect 509956 361800 513286 361856
rect 513342 361800 513347 361856
rect 509956 361798 513347 361800
rect 447133 361795 447199 361798
rect 513281 361795 513347 361798
rect 512821 361314 512887 361317
rect 509956 361312 512887 361314
rect 509956 361256 512826 361312
rect 512882 361256 512887 361312
rect 509956 361254 512887 361256
rect 512821 361251 512887 361254
rect 447133 361178 447199 361181
rect 447133 361176 450156 361178
rect 447133 361120 447138 361176
rect 447194 361120 450156 361176
rect 447133 361118 450156 361120
rect 447133 361115 447199 361118
rect 512361 360770 512427 360773
rect 509956 360768 512427 360770
rect 509956 360712 512366 360768
rect 512422 360712 512427 360768
rect 509956 360710 512427 360712
rect 512361 360707 512427 360710
rect 447317 360498 447383 360501
rect 447317 360496 450156 360498
rect 447317 360440 447322 360496
rect 447378 360440 450156 360496
rect 447317 360438 450156 360440
rect 447317 360435 447383 360438
rect 513281 360226 513347 360229
rect 509956 360224 513347 360226
rect 509956 360168 513286 360224
rect 513342 360168 513347 360224
rect 509956 360166 513347 360168
rect 513281 360163 513347 360166
rect 447317 359818 447383 359821
rect 447317 359816 450156 359818
rect 447317 359760 447322 359816
rect 447378 359760 450156 359816
rect 447317 359758 450156 359760
rect 447317 359755 447383 359758
rect 512913 359682 512979 359685
rect 509956 359680 512979 359682
rect 509956 359624 512918 359680
rect 512974 359624 512979 359680
rect 509956 359622 512979 359624
rect 512913 359619 512979 359622
rect 362217 359546 362283 359549
rect 359812 359544 362283 359546
rect 359812 359488 362222 359544
rect 362278 359488 362283 359544
rect 359812 359486 362283 359488
rect 362217 359483 362283 359486
rect 447133 359138 447199 359141
rect 512361 359138 512427 359141
rect 447133 359136 450156 359138
rect 447133 359080 447138 359136
rect 447194 359080 450156 359136
rect 447133 359078 450156 359080
rect 509956 359136 512427 359138
rect 509956 359080 512366 359136
rect 512422 359080 512427 359136
rect 509956 359078 512427 359080
rect 447133 359075 447199 359078
rect 512361 359075 512427 359078
rect 512453 358594 512519 358597
rect 509956 358592 512519 358594
rect -960 358458 480 358548
rect 509956 358536 512458 358592
rect 512514 358536 512519 358592
rect 509956 358534 512519 358536
rect 512453 358531 512519 358534
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 448421 358458 448487 358461
rect 448421 358456 450156 358458
rect 448421 358400 448426 358456
rect 448482 358400 450156 358456
rect 448421 358398 450156 358400
rect 448421 358395 448487 358398
rect 448973 357778 449039 357781
rect 448973 357776 450156 357778
rect 448973 357720 448978 357776
rect 449034 357720 450156 357776
rect 448973 357718 450156 357720
rect 448973 357715 449039 357718
rect 509558 357645 509618 358020
rect 509417 357642 509483 357645
rect 509374 357640 509483 357642
rect 509374 357584 509422 357640
rect 509478 357584 509483 357640
rect 509374 357579 509483 357584
rect 509558 357640 509667 357645
rect 509558 357584 509606 357640
rect 509662 357584 509667 357640
rect 509558 357582 509667 357584
rect 509601 357579 509667 357582
rect 509374 357476 509434 357579
rect 449801 357098 449867 357101
rect 449801 357096 450156 357098
rect 449801 357040 449806 357096
rect 449862 357040 450156 357096
rect 449801 357038 450156 357040
rect 449801 357035 449867 357038
rect 513557 356962 513623 356965
rect 509956 356960 513623 356962
rect 509956 356904 513562 356960
rect 513618 356904 513623 356960
rect 509956 356902 513623 356904
rect 513557 356899 513623 356902
rect 449617 356418 449683 356421
rect 512913 356418 512979 356421
rect 449617 356416 450156 356418
rect 449617 356360 449622 356416
rect 449678 356360 450156 356416
rect 449617 356358 450156 356360
rect 509956 356416 512979 356418
rect 509956 356360 512918 356416
rect 512974 356360 512979 356416
rect 509956 356358 512979 356360
rect 449617 356355 449683 356358
rect 512913 356355 512979 356358
rect 510797 355874 510863 355877
rect 509956 355872 510863 355874
rect 509956 355816 510802 355872
rect 510858 355816 510863 355872
rect 509956 355814 510863 355816
rect 510797 355811 510863 355814
rect 449065 355738 449131 355741
rect 449065 355736 450156 355738
rect 449065 355680 449070 355736
rect 449126 355680 450156 355736
rect 449065 355678 450156 355680
rect 449065 355675 449131 355678
rect 513281 355330 513347 355333
rect 509956 355328 513347 355330
rect 509956 355272 513286 355328
rect 513342 355272 513347 355328
rect 509956 355270 513347 355272
rect 513281 355267 513347 355270
rect 449709 355058 449775 355061
rect 449709 355056 450156 355058
rect 449709 355000 449714 355056
rect 449770 355000 450156 355056
rect 449709 354998 450156 355000
rect 449709 354995 449775 354998
rect 511533 354786 511599 354789
rect 509956 354784 511599 354786
rect 509956 354728 511538 354784
rect 511594 354728 511599 354784
rect 509956 354726 511599 354728
rect 511533 354723 511599 354726
rect 449433 354378 449499 354381
rect 449433 354376 450156 354378
rect 449433 354320 449438 354376
rect 449494 354320 450156 354376
rect 449433 354318 450156 354320
rect 449433 354315 449499 354318
rect 510889 354242 510955 354245
rect 509956 354240 510955 354242
rect 509956 354184 510894 354240
rect 510950 354184 510955 354240
rect 509956 354182 510955 354184
rect 510889 354179 510955 354182
rect 447869 353698 447935 353701
rect 512361 353698 512427 353701
rect 447869 353696 450156 353698
rect 447869 353640 447874 353696
rect 447930 353640 450156 353696
rect 447869 353638 450156 353640
rect 509956 353696 512427 353698
rect 509956 353640 512366 353696
rect 512422 353640 512427 353696
rect 509956 353638 512427 353640
rect 447869 353635 447935 353638
rect 512361 353635 512427 353638
rect 450261 353290 450327 353293
rect 450261 353288 450370 353290
rect 450261 353232 450266 353288
rect 450322 353232 450370 353288
rect 450261 353227 450370 353232
rect 450310 352988 450370 353227
rect 512821 353154 512887 353157
rect 509956 353152 512887 353154
rect 509956 353096 512826 353152
rect 512882 353096 512887 353152
rect 509956 353094 512887 353096
rect 512821 353091 512887 353094
rect 512361 352610 512427 352613
rect 509956 352608 512427 352610
rect 509956 352552 512366 352608
rect 512422 352552 512427 352608
rect 509956 352550 512427 352552
rect 512361 352547 512427 352550
rect 447777 352338 447843 352341
rect 447777 352336 450156 352338
rect 447777 352280 447782 352336
rect 447838 352280 450156 352336
rect 447777 352278 450156 352280
rect 447777 352275 447843 352278
rect 513281 352066 513347 352069
rect 509956 352064 513347 352066
rect 509956 352008 513286 352064
rect 513342 352008 513347 352064
rect 509956 352006 513347 352008
rect 513281 352003 513347 352006
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 449893 351114 449959 351117
rect 450126 351114 450186 351628
rect 513005 351522 513071 351525
rect 509956 351520 513071 351522
rect 509956 351464 513010 351520
rect 513066 351464 513071 351520
rect 509956 351462 513071 351464
rect 513005 351459 513071 351462
rect 449893 351112 450186 351114
rect 449893 351056 449898 351112
rect 449954 351056 450186 351112
rect 449893 351054 450186 351056
rect 449893 351051 449959 351054
rect 447133 350978 447199 350981
rect 512361 350978 512427 350981
rect 447133 350976 450156 350978
rect 447133 350920 447138 350976
rect 447194 350920 450156 350976
rect 447133 350918 450156 350920
rect 509956 350976 512427 350978
rect 509956 350920 512366 350976
rect 512422 350920 512427 350976
rect 509956 350918 512427 350920
rect 447133 350915 447199 350918
rect 512361 350915 512427 350918
rect 513189 350434 513255 350437
rect 509956 350432 513255 350434
rect 509956 350376 513194 350432
rect 513250 350376 513255 350432
rect 509956 350374 513255 350376
rect 513189 350371 513255 350374
rect 449709 350298 449775 350301
rect 449709 350296 450156 350298
rect 449709 350240 449714 350296
rect 449770 350240 450156 350296
rect 449709 350238 450156 350240
rect 449709 350235 449775 350238
rect 449985 350026 450051 350029
rect 449985 350024 450186 350026
rect 449985 349968 449990 350024
rect 450046 349968 450186 350024
rect 449985 349966 450186 349968
rect 449985 349963 450051 349966
rect 450126 349588 450186 349966
rect 513005 349890 513071 349893
rect 509956 349888 513071 349890
rect 509956 349832 513010 349888
rect 513066 349832 513071 349888
rect 509956 349830 513071 349832
rect 513005 349827 513071 349830
rect 512361 349346 512427 349349
rect 509956 349344 512427 349346
rect 509956 349288 512366 349344
rect 512422 349288 512427 349344
rect 509956 349286 512427 349288
rect 512361 349283 512427 349286
rect 450629 349074 450695 349077
rect 450629 349072 450738 349074
rect 450629 349016 450634 349072
rect 450690 349016 450738 349072
rect 450629 349011 450738 349016
rect 450678 348908 450738 349011
rect 450353 348666 450419 348669
rect 450310 348664 450419 348666
rect 450310 348608 450358 348664
rect 450414 348608 450419 348664
rect 450310 348603 450419 348608
rect 361757 348530 361823 348533
rect 359812 348528 361823 348530
rect 359812 348472 361762 348528
rect 361818 348472 361823 348528
rect 359812 348470 361823 348472
rect 361757 348467 361823 348470
rect 450310 348228 450370 348603
rect 509742 348397 509802 348772
rect 509742 348392 509851 348397
rect 509742 348336 509790 348392
rect 509846 348336 509851 348392
rect 509742 348334 509851 348336
rect 509785 348331 509851 348334
rect 513005 348258 513071 348261
rect 509956 348256 513071 348258
rect 509956 348200 513010 348256
rect 513066 348200 513071 348256
rect 509956 348198 513071 348200
rect 513005 348195 513071 348198
rect 510981 347714 511047 347717
rect 509956 347712 511047 347714
rect 509956 347656 510986 347712
rect 511042 347656 511047 347712
rect 509956 347654 511047 347656
rect 510981 347651 511047 347654
rect 447133 347578 447199 347581
rect 447133 347576 450156 347578
rect 447133 347520 447138 347576
rect 447194 347520 450156 347576
rect 447133 347518 450156 347520
rect 447133 347515 447199 347518
rect 450169 347306 450235 347309
rect 450126 347304 450235 347306
rect 450126 347248 450174 347304
rect 450230 347248 450235 347304
rect 450126 347243 450235 347248
rect 450126 346868 450186 347243
rect 513281 347170 513347 347173
rect 509956 347168 513347 347170
rect 509956 347112 513286 347168
rect 513342 347112 513347 347168
rect 509956 347110 513347 347112
rect 513281 347107 513347 347110
rect 513097 346626 513163 346629
rect 509956 346624 513163 346626
rect 509956 346568 513102 346624
rect 513158 346568 513163 346624
rect 509956 346566 513163 346568
rect 513097 346563 513163 346566
rect 450077 346354 450143 346357
rect 450077 346352 450186 346354
rect 450077 346296 450082 346352
rect 450138 346296 450186 346352
rect 450077 346291 450186 346296
rect 450126 346188 450186 346291
rect 511073 346082 511139 346085
rect 509956 346080 511139 346082
rect 509956 346024 511078 346080
rect 511134 346024 511139 346080
rect 509956 346022 511139 346024
rect 511073 346019 511139 346022
rect 449617 345538 449683 345541
rect 512361 345538 512427 345541
rect 449617 345536 450156 345538
rect -960 345402 480 345492
rect 449617 345480 449622 345536
rect 449678 345480 450156 345536
rect 449617 345478 450156 345480
rect 509956 345536 512427 345538
rect 509956 345480 512366 345536
rect 512422 345480 512427 345536
rect 509956 345478 512427 345480
rect 449617 345475 449683 345478
rect 512361 345475 512427 345478
rect 3509 345402 3575 345405
rect -960 345400 3575 345402
rect -960 345344 3514 345400
rect 3570 345344 3575 345400
rect -960 345342 3575 345344
rect -960 345252 480 345342
rect 3509 345339 3575 345342
rect 512545 344994 512611 344997
rect 509956 344992 512611 344994
rect 509956 344936 512550 344992
rect 512606 344936 512611 344992
rect 509956 344934 512611 344936
rect 512545 344931 512611 344934
rect 448421 344858 448487 344861
rect 448421 344856 450156 344858
rect 448421 344800 448426 344856
rect 448482 344800 450156 344856
rect 448421 344798 450156 344800
rect 448421 344795 448487 344798
rect 447317 344178 447383 344181
rect 447317 344176 450156 344178
rect 447317 344120 447322 344176
rect 447378 344120 450156 344176
rect 447317 344118 450156 344120
rect 447317 344115 447383 344118
rect 509742 344045 509802 344420
rect 509693 344040 509802 344045
rect 509693 343984 509698 344040
rect 509754 343984 509802 344040
rect 509693 343982 509802 343984
rect 509693 343979 509759 343982
rect 512637 343906 512703 343909
rect 509956 343904 512703 343906
rect 509956 343848 512642 343904
rect 512698 343848 512703 343904
rect 509956 343846 512703 343848
rect 512637 343843 512703 343846
rect 447501 343498 447567 343501
rect 449801 343498 449867 343501
rect 447501 343496 450156 343498
rect 447501 343440 447506 343496
rect 447562 343440 449806 343496
rect 449862 343440 450156 343496
rect 447501 343438 450156 343440
rect 447501 343435 447567 343438
rect 449801 343435 449867 343438
rect 513005 343362 513071 343365
rect 509956 343360 513071 343362
rect 509956 343304 513010 343360
rect 513066 343304 513071 343360
rect 509956 343302 513071 343304
rect 513005 343299 513071 343302
rect 509926 342413 509986 342788
rect 509877 342408 509986 342413
rect 509877 342352 509882 342408
rect 509938 342352 509986 342408
rect 509877 342350 509986 342352
rect 509877 342347 509943 342350
rect 513281 342274 513347 342277
rect 509956 342272 513347 342274
rect 509956 342216 513286 342272
rect 513342 342216 513347 342272
rect 509956 342214 513347 342216
rect 513281 342211 513347 342214
rect 447225 342138 447291 342141
rect 447225 342136 450156 342138
rect 447225 342080 447230 342136
rect 447286 342080 450156 342136
rect 447225 342078 450156 342080
rect 447225 342075 447291 342078
rect 513005 341730 513071 341733
rect 509956 341728 513071 341730
rect 509956 341672 513010 341728
rect 513066 341672 513071 341728
rect 509956 341670 513071 341672
rect 513005 341667 513071 341670
rect 447133 341458 447199 341461
rect 447133 341456 450156 341458
rect 447133 341400 447138 341456
rect 447194 341400 450156 341456
rect 447133 341398 450156 341400
rect 447133 341395 447199 341398
rect 513281 341186 513347 341189
rect 509956 341184 513347 341186
rect 509956 341128 513286 341184
rect 513342 341128 513347 341184
rect 509956 341126 513347 341128
rect 513281 341123 513347 341126
rect 447133 340778 447199 340781
rect 447133 340776 450156 340778
rect 447133 340720 447138 340776
rect 447194 340720 450156 340776
rect 447133 340718 450156 340720
rect 447133 340715 447199 340718
rect 513189 340642 513255 340645
rect 509956 340640 513255 340642
rect 509956 340584 513194 340640
rect 513250 340584 513255 340640
rect 509956 340582 513255 340584
rect 513189 340579 513255 340582
rect 447225 340098 447291 340101
rect 513281 340098 513347 340101
rect 447225 340096 450156 340098
rect 447225 340040 447230 340096
rect 447286 340040 450156 340096
rect 447225 340038 450156 340040
rect 509956 340096 513347 340098
rect 509956 340040 513286 340096
rect 513342 340040 513347 340096
rect 509956 340038 513347 340040
rect 447225 340035 447291 340038
rect 513281 340035 513347 340038
rect 513097 339554 513163 339557
rect 509956 339552 513163 339554
rect 509956 339496 513102 339552
rect 513158 339496 513163 339552
rect 509956 339494 513163 339496
rect 513097 339491 513163 339494
rect 447225 339418 447291 339421
rect 447225 339416 450156 339418
rect 447225 339360 447230 339416
rect 447286 339360 450156 339416
rect 447225 339358 450156 339360
rect 447225 339355 447291 339358
rect 512821 339010 512887 339013
rect 509956 339008 512887 339010
rect 509956 338952 512826 339008
rect 512882 338952 512887 339008
rect 509956 338950 512887 338952
rect 512821 338947 512887 338950
rect 447133 338738 447199 338741
rect 447133 338736 450156 338738
rect 447133 338680 447138 338736
rect 447194 338680 450156 338736
rect 447133 338678 450156 338680
rect 447133 338675 447199 338678
rect 512637 338466 512703 338469
rect 509956 338464 512703 338466
rect 509956 338408 512642 338464
rect 512698 338408 512703 338464
rect 583520 338452 584960 338692
rect 509956 338406 512703 338408
rect 512637 338403 512703 338406
rect 447225 338058 447291 338061
rect 447225 338056 450156 338058
rect 447225 338000 447230 338056
rect 447286 338000 450156 338056
rect 447225 337998 450156 338000
rect 447225 337995 447291 337998
rect 513281 337922 513347 337925
rect 509956 337920 513347 337922
rect 509956 337864 513286 337920
rect 513342 337864 513347 337920
rect 509956 337862 513347 337864
rect 513281 337859 513347 337862
rect 361757 337514 361823 337517
rect 359812 337512 361823 337514
rect 359812 337456 361762 337512
rect 361818 337456 361823 337512
rect 359812 337454 361823 337456
rect 361757 337451 361823 337454
rect 447133 337378 447199 337381
rect 512637 337378 512703 337381
rect 447133 337376 450156 337378
rect 447133 337320 447138 337376
rect 447194 337320 450156 337376
rect 447133 337318 450156 337320
rect 509956 337376 512703 337378
rect 509956 337320 512642 337376
rect 512698 337320 512703 337376
rect 509956 337318 512703 337320
rect 447133 337315 447199 337318
rect 512637 337315 512703 337318
rect 513281 336834 513347 336837
rect 509956 336832 513347 336834
rect 509956 336776 513286 336832
rect 513342 336776 513347 336832
rect 509956 336774 513347 336776
rect 513281 336771 513347 336774
rect 447225 336698 447291 336701
rect 447225 336696 450156 336698
rect 447225 336640 447230 336696
rect 447286 336640 450156 336696
rect 447225 336638 450156 336640
rect 447225 336635 447291 336638
rect 513281 336290 513347 336293
rect 509956 336288 513347 336290
rect 509956 336232 513286 336288
rect 513342 336232 513347 336288
rect 509956 336230 513347 336232
rect 513281 336227 513347 336230
rect 447133 336018 447199 336021
rect 447133 336016 450156 336018
rect 447133 335960 447138 336016
rect 447194 335960 450156 336016
rect 447133 335958 450156 335960
rect 447133 335955 447199 335958
rect 511165 335746 511231 335749
rect 509956 335744 511231 335746
rect 509956 335688 511170 335744
rect 511226 335688 511231 335744
rect 509956 335686 511231 335688
rect 511165 335683 511231 335686
rect 424133 335474 424199 335477
rect 425830 335474 425836 335476
rect 424133 335472 425836 335474
rect 424133 335416 424138 335472
rect 424194 335416 425836 335472
rect 424133 335414 425836 335416
rect 424133 335411 424199 335414
rect 425830 335412 425836 335414
rect 425900 335412 425906 335476
rect 447501 335338 447567 335341
rect 447501 335336 450156 335338
rect 447501 335280 447506 335336
rect 447562 335280 450156 335336
rect 447501 335278 450156 335280
rect 447501 335275 447567 335278
rect 518014 335202 518020 335204
rect 509956 335142 518020 335202
rect 518014 335140 518020 335142
rect 518084 335140 518090 335204
rect 447225 334658 447291 334661
rect 512729 334658 512795 334661
rect 447225 334656 450156 334658
rect 447225 334600 447230 334656
rect 447286 334600 450156 334656
rect 447225 334598 450156 334600
rect 509956 334656 512795 334658
rect 509956 334600 512734 334656
rect 512790 334600 512795 334656
rect 509956 334598 512795 334600
rect 447225 334595 447291 334598
rect 512729 334595 512795 334598
rect 420729 334522 420795 334525
rect 421046 334522 421052 334524
rect 420729 334520 421052 334522
rect 420729 334464 420734 334520
rect 420790 334464 421052 334520
rect 420729 334462 421052 334464
rect 420729 334459 420795 334462
rect 421046 334460 421052 334462
rect 421116 334460 421122 334524
rect 428089 334522 428155 334525
rect 428406 334522 428412 334524
rect 428089 334520 428412 334522
rect 428089 334464 428094 334520
rect 428150 334464 428412 334520
rect 428089 334462 428412 334464
rect 428089 334459 428155 334462
rect 428406 334460 428412 334462
rect 428476 334460 428482 334524
rect 509969 334250 510035 334253
rect 509926 334248 510035 334250
rect 509926 334192 509974 334248
rect 510030 334192 510035 334248
rect 509926 334187 510035 334192
rect 509926 334084 509986 334187
rect 447133 333978 447199 333981
rect 447133 333976 450156 333978
rect 447133 333920 447138 333976
rect 447194 333920 450156 333976
rect 447133 333918 450156 333920
rect 447133 333915 447199 333918
rect 511022 333570 511028 333572
rect 509956 333510 511028 333570
rect 511022 333508 511028 333510
rect 511092 333508 511098 333572
rect 447225 333298 447291 333301
rect 447225 333296 450156 333298
rect 447225 333240 447230 333296
rect 447286 333240 450156 333296
rect 447225 333238 450156 333240
rect 447225 333235 447291 333238
rect 425830 332964 425836 333028
rect 425900 333026 425906 333028
rect 429193 333026 429259 333029
rect 515070 333026 515076 333028
rect 425900 333024 429259 333026
rect 425900 332968 429198 333024
rect 429254 332968 429259 333024
rect 425900 332966 429259 332968
rect 509956 332966 515076 333026
rect 425900 332964 425906 332966
rect 429193 332963 429259 332966
rect 515070 332964 515076 332966
rect 515140 332964 515146 333028
rect 432597 332890 432663 332893
rect 429916 332888 432663 332890
rect 429916 332832 432602 332888
rect 432658 332832 432663 332888
rect 429916 332830 432663 332832
rect 432597 332827 432663 332830
rect 447409 332618 447475 332621
rect 448421 332618 448487 332621
rect 447409 332616 450156 332618
rect 447409 332560 447414 332616
rect 447470 332560 448426 332616
rect 448482 332560 450156 332616
rect 447409 332558 450156 332560
rect 447409 332555 447475 332558
rect 448421 332555 448487 332558
rect 512913 332482 512979 332485
rect 509956 332480 512979 332482
rect -960 332196 480 332436
rect 509956 332424 512918 332480
rect 512974 332424 512979 332480
rect 509956 332422 512979 332424
rect 512913 332419 512979 332422
rect 447133 331938 447199 331941
rect 510061 331938 510127 331941
rect 447133 331936 450156 331938
rect 447133 331880 447138 331936
rect 447194 331880 450156 331936
rect 447133 331878 450156 331880
rect 509956 331936 510127 331938
rect 509956 331880 510066 331936
rect 510122 331880 510127 331936
rect 509956 331878 510127 331880
rect 447133 331875 447199 331878
rect 510061 331875 510127 331878
rect 514702 331394 514708 331396
rect 509956 331334 514708 331394
rect 514702 331332 514708 331334
rect 514772 331332 514778 331396
rect 447225 331258 447291 331261
rect 447225 331256 450156 331258
rect 447225 331200 447230 331256
rect 447286 331200 450156 331256
rect 447225 331198 450156 331200
rect 447225 331195 447291 331198
rect 517830 330850 517836 330852
rect 509956 330790 517836 330850
rect 517830 330788 517836 330790
rect 517900 330788 517906 330852
rect 447133 330578 447199 330581
rect 447133 330576 450156 330578
rect 447133 330520 447138 330576
rect 447194 330520 450156 330576
rect 447133 330518 450156 330520
rect 447133 330515 447199 330518
rect 510153 330306 510219 330309
rect 509956 330304 510219 330306
rect 509956 330248 510158 330304
rect 510214 330248 510219 330304
rect 509956 330246 510219 330248
rect 510153 330243 510219 330246
rect 447593 329898 447659 329901
rect 447593 329896 450156 329898
rect 447593 329840 447598 329896
rect 447654 329840 450156 329896
rect 447593 329838 450156 329840
rect 447593 329835 447659 329838
rect 510838 329762 510844 329764
rect 509956 329702 510844 329762
rect 510838 329700 510844 329702
rect 510908 329700 510914 329764
rect 432965 329218 433031 329221
rect 429916 329216 433031 329218
rect 429916 329160 432970 329216
rect 433026 329160 433031 329216
rect 429916 329158 433031 329160
rect 432965 329155 433031 329158
rect 447133 329218 447199 329221
rect 448278 329218 448284 329220
rect 447133 329216 448284 329218
rect 447133 329160 447138 329216
rect 447194 329160 448284 329216
rect 447133 329158 448284 329160
rect 447133 329155 447199 329158
rect 448278 329156 448284 329158
rect 448348 329218 448354 329220
rect 512729 329218 512795 329221
rect 448348 329158 450156 329218
rect 509956 329216 512795 329218
rect 509956 329160 512734 329216
rect 512790 329160 512795 329216
rect 509956 329158 512795 329160
rect 448348 329156 448354 329158
rect 512729 329155 512795 329158
rect 514150 328674 514156 328676
rect 509956 328614 514156 328674
rect 514150 328612 514156 328614
rect 514220 328612 514226 328676
rect 447409 328538 447475 328541
rect 448329 328538 448395 328541
rect 447409 328536 450156 328538
rect 447409 328480 447414 328536
rect 447470 328480 448334 328536
rect 448390 328480 450156 328536
rect 447409 328478 450156 328480
rect 447409 328475 447475 328478
rect 448329 328475 448395 328478
rect 510470 328130 510476 328132
rect 509956 328070 510476 328130
rect 510470 328068 510476 328070
rect 510540 328068 510546 328132
rect 447501 327858 447567 327861
rect 447501 327856 450156 327858
rect 447501 327800 447506 327856
rect 447562 327800 450156 327856
rect 447501 327798 450156 327800
rect 447501 327795 447567 327798
rect 516174 327586 516180 327588
rect 509956 327526 516180 327586
rect 516174 327524 516180 327526
rect 516244 327524 516250 327588
rect 448237 327178 448303 327181
rect 448237 327176 450156 327178
rect 448237 327120 448242 327176
rect 448298 327120 450156 327176
rect 448237 327118 450156 327120
rect 448237 327115 448303 327118
rect 514886 327042 514892 327044
rect 509956 326982 514892 327042
rect 514886 326980 514892 326982
rect 514956 326980 514962 327044
rect 362217 326498 362283 326501
rect 359812 326496 362283 326498
rect 359812 326440 362222 326496
rect 362278 326440 362283 326496
rect 359812 326438 362283 326440
rect 362217 326435 362283 326438
rect 447409 326498 447475 326501
rect 510654 326498 510660 326500
rect 447409 326496 450156 326498
rect 447409 326440 447414 326496
rect 447470 326440 450156 326496
rect 447409 326438 450156 326440
rect 509956 326438 510660 326498
rect 447409 326435 447475 326438
rect 510654 326436 510660 326438
rect 510724 326436 510730 326500
rect 447961 325818 448027 325821
rect 509926 325818 509986 325924
rect 511901 325818 511967 325821
rect 447961 325816 450156 325818
rect 447961 325760 447966 325816
rect 448022 325760 450156 325816
rect 447961 325758 450156 325760
rect 509926 325816 511967 325818
rect 509926 325760 511906 325816
rect 511962 325760 511967 325816
rect 509926 325758 511967 325760
rect 447961 325755 448027 325758
rect 511901 325755 511967 325758
rect 432689 325546 432755 325549
rect 429916 325544 432755 325546
rect 429916 325488 432694 325544
rect 432750 325488 432755 325544
rect 429916 325486 432755 325488
rect 432689 325483 432755 325486
rect 512821 325410 512887 325413
rect 509956 325408 512887 325410
rect 509956 325352 512826 325408
rect 512882 325352 512887 325408
rect 509956 325350 512887 325352
rect 512821 325347 512887 325350
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 448237 325138 448303 325141
rect 448237 325136 450156 325138
rect 448237 325080 448242 325136
rect 448298 325080 450156 325136
rect 583520 325124 584960 325214
rect 448237 325078 450156 325080
rect 448237 325075 448303 325078
rect 514334 324866 514340 324868
rect 509956 324806 514340 324866
rect 514334 324804 514340 324806
rect 514404 324804 514410 324868
rect 449525 324458 449591 324461
rect 449525 324456 450156 324458
rect 449525 324400 449530 324456
rect 449586 324400 450156 324456
rect 449525 324398 450156 324400
rect 449525 324395 449591 324398
rect 510654 324396 510660 324460
rect 510724 324458 510730 324460
rect 511206 324458 511212 324460
rect 510724 324398 511212 324458
rect 510724 324396 510730 324398
rect 511206 324396 511212 324398
rect 511276 324396 511282 324460
rect 510654 324322 510660 324324
rect 509956 324262 510660 324322
rect 510654 324260 510660 324262
rect 510724 324260 510730 324324
rect 509742 323373 509802 323748
rect 509693 323368 509802 323373
rect 509693 323312 509698 323368
rect 509754 323312 509802 323368
rect 509693 323310 509802 323312
rect 509693 323307 509759 323310
rect 509785 322962 509851 322965
rect 509190 322960 509851 322962
rect 509190 322904 509790 322960
rect 509846 322904 509851 322960
rect 509190 322902 509851 322904
rect 508446 322764 508452 322828
rect 508516 322826 508522 322828
rect 509190 322826 509250 322902
rect 509785 322899 509851 322902
rect 508516 322766 509250 322826
rect 508516 322764 508522 322766
rect 509182 322628 509188 322692
rect 509252 322690 509258 322692
rect 509926 322690 509986 323204
rect 509252 322630 509986 322690
rect 509252 322628 509258 322630
rect 507209 322282 507275 322285
rect 511901 322282 511967 322285
rect 507209 322280 511967 322282
rect 507209 322224 507214 322280
rect 507270 322224 511906 322280
rect 511962 322224 511967 322280
rect 507209 322222 511967 322224
rect 507209 322219 507275 322222
rect 511901 322219 511967 322222
rect 509509 322146 509575 322149
rect 466410 322144 509575 322146
rect 466410 322088 509514 322144
rect 509570 322088 509575 322144
rect 466410 322086 509575 322088
rect 460197 322010 460263 322013
rect 466410 322010 466470 322086
rect 509509 322083 509575 322086
rect 460197 322008 466470 322010
rect 460197 321952 460202 322008
rect 460258 321952 466470 322008
rect 460197 321950 466470 321952
rect 460197 321947 460263 321950
rect 432781 321874 432847 321877
rect 429916 321872 432847 321874
rect 429916 321816 432786 321872
rect 432842 321816 432847 321872
rect 429916 321814 432847 321816
rect 432781 321811 432847 321814
rect 447726 321812 447732 321876
rect 447796 321874 447802 321876
rect 462221 321874 462287 321877
rect 447796 321872 462287 321874
rect 447796 321816 462226 321872
rect 462282 321816 462287 321872
rect 447796 321814 462287 321816
rect 447796 321812 447802 321814
rect 462221 321811 462287 321814
rect 445201 321738 445267 321741
rect 482921 321738 482987 321741
rect 445201 321736 482987 321738
rect 445201 321680 445206 321736
rect 445262 321680 482926 321736
rect 482982 321680 482987 321736
rect 445201 321678 482987 321680
rect 445201 321675 445267 321678
rect 482921 321675 482987 321678
rect 446305 321602 446371 321605
rect 483749 321602 483815 321605
rect 446305 321600 483815 321602
rect 446305 321544 446310 321600
rect 446366 321544 483754 321600
rect 483810 321544 483815 321600
rect 446305 321542 483815 321544
rect 446305 321539 446371 321542
rect 483749 321539 483815 321542
rect 460013 321466 460079 321469
rect 556286 321466 556292 321468
rect 460013 321464 556292 321466
rect 460013 321408 460018 321464
rect 460074 321408 556292 321464
rect 460013 321406 556292 321408
rect 460013 321403 460079 321406
rect 556286 321404 556292 321406
rect 556356 321404 556362 321468
rect 449566 321268 449572 321332
rect 449636 321330 449642 321332
rect 482369 321330 482435 321333
rect 449636 321328 482435 321330
rect 449636 321272 482374 321328
rect 482430 321272 482435 321328
rect 449636 321270 482435 321272
rect 449636 321268 449642 321270
rect 482369 321267 482435 321270
rect 444046 321132 444052 321196
rect 444116 321194 444122 321196
rect 461669 321194 461735 321197
rect 444116 321192 461735 321194
rect 444116 321136 461674 321192
rect 461730 321136 461735 321192
rect 444116 321134 461735 321136
rect 444116 321132 444122 321134
rect 461669 321131 461735 321134
rect 446765 320106 446831 320109
rect 483197 320106 483263 320109
rect 446765 320104 483263 320106
rect 446765 320048 446770 320104
rect 446826 320048 483202 320104
rect 483258 320048 483263 320104
rect 446765 320046 483263 320048
rect 446765 320043 446831 320046
rect 483197 320043 483263 320046
rect 450670 319908 450676 319972
rect 450740 319970 450746 319972
rect 482645 319970 482711 319973
rect 450740 319968 482711 319970
rect 450740 319912 482650 319968
rect 482706 319912 482711 319968
rect 450740 319910 482711 319912
rect 450740 319908 450746 319910
rect 482645 319907 482711 319910
rect 444230 319772 444236 319836
rect 444300 319834 444306 319836
rect 471605 319834 471671 319837
rect 444300 319832 471671 319834
rect 444300 319776 471610 319832
rect 471666 319776 471671 319832
rect 444300 319774 471671 319776
rect 444300 319772 444306 319774
rect 471605 319771 471671 319774
rect 446581 319698 446647 319701
rect 472709 319698 472775 319701
rect 446581 319696 472775 319698
rect 446581 319640 446586 319696
rect 446642 319640 472714 319696
rect 472770 319640 472775 319696
rect 446581 319638 472775 319640
rect 446581 319635 446647 319638
rect 472709 319635 472775 319638
rect 450486 319500 450492 319564
rect 450556 319562 450562 319564
rect 472157 319562 472223 319565
rect 450556 319560 472223 319562
rect 450556 319504 472162 319560
rect 472218 319504 472223 319560
rect 450556 319502 472223 319504
rect 450556 319500 450562 319502
rect 472157 319499 472223 319502
rect 502241 319426 502307 319429
rect 538806 319426 538812 319428
rect 502241 319424 538812 319426
rect -960 319290 480 319380
rect 502241 319368 502246 319424
rect 502302 319368 538812 319424
rect 502241 319366 538812 319368
rect 502241 319363 502307 319366
rect 538806 319364 538812 319366
rect 538876 319364 538882 319428
rect 3877 319290 3943 319293
rect -960 319288 3943 319290
rect -960 319232 3882 319288
rect 3938 319232 3943 319288
rect -960 319230 3943 319232
rect -960 319140 480 319230
rect 3877 319227 3943 319230
rect 432597 318202 432663 318205
rect 429916 318200 432663 318202
rect 429916 318144 432602 318200
rect 432658 318144 432663 318200
rect 429916 318142 432663 318144
rect 432597 318139 432663 318142
rect 454953 317250 455019 317253
rect 511206 317250 511212 317252
rect 454953 317248 511212 317250
rect 454953 317192 454958 317248
rect 455014 317192 511212 317248
rect 454953 317190 511212 317192
rect 454953 317187 455019 317190
rect 511206 317188 511212 317190
rect 511276 317188 511282 317252
rect 458950 317052 458956 317116
rect 459020 317114 459026 317116
rect 515070 317114 515076 317116
rect 459020 317054 515076 317114
rect 459020 317052 459026 317054
rect 515070 317052 515076 317054
rect 515140 317052 515146 317116
rect 453297 316978 453363 316981
rect 510654 316978 510660 316980
rect 453297 316976 510660 316978
rect 453297 316920 453302 316976
rect 453358 316920 510660 316976
rect 453297 316918 510660 316920
rect 453297 316915 453363 316918
rect 510654 316916 510660 316918
rect 510724 316916 510730 316980
rect 458766 316780 458772 316844
rect 458836 316842 458842 316844
rect 516961 316842 517027 316845
rect 458836 316840 517027 316842
rect 458836 316784 516966 316840
rect 517022 316784 517027 316840
rect 458836 316782 517027 316784
rect 458836 316780 458842 316782
rect 516961 316779 517027 316782
rect 454677 316706 454743 316709
rect 508998 316706 509004 316708
rect 454677 316704 509004 316706
rect 454677 316648 454682 316704
rect 454738 316648 509004 316704
rect 454677 316646 509004 316648
rect 454677 316643 454743 316646
rect 508998 316644 509004 316646
rect 509068 316644 509074 316708
rect 361757 315482 361823 315485
rect 359812 315480 361823 315482
rect 359812 315424 361762 315480
rect 361818 315424 361823 315480
rect 359812 315422 361823 315424
rect 361757 315419 361823 315422
rect 495801 315346 495867 315349
rect 542670 315346 542676 315348
rect 495801 315344 542676 315346
rect 495801 315288 495806 315344
rect 495862 315288 542676 315344
rect 495801 315286 542676 315288
rect 495801 315283 495867 315286
rect 542670 315284 542676 315286
rect 542740 315284 542746 315348
rect 432689 314530 432755 314533
rect 429916 314528 432755 314530
rect 429916 314472 432694 314528
rect 432750 314472 432755 314528
rect 429916 314470 432755 314472
rect 432689 314467 432755 314470
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 432597 310858 432663 310861
rect 429916 310856 432663 310858
rect 429916 310800 432602 310856
rect 432658 310800 432663 310856
rect 429916 310798 432663 310800
rect 432597 310795 432663 310798
rect 432413 307186 432479 307189
rect 429916 307184 432479 307186
rect 429916 307128 432418 307184
rect 432474 307128 432479 307184
rect 429916 307126 432479 307128
rect 432413 307123 432479 307126
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 361757 304466 361823 304469
rect 359812 304464 361823 304466
rect 359812 304408 361762 304464
rect 361818 304408 361823 304464
rect 359812 304406 361823 304408
rect 361757 304403 361823 304406
rect 403893 302834 403959 302837
rect 510470 302834 510476 302836
rect 403893 302832 510476 302834
rect 403893 302776 403898 302832
rect 403954 302776 510476 302832
rect 403893 302774 510476 302776
rect 403893 302771 403959 302774
rect 510470 302772 510476 302774
rect 510540 302772 510546 302836
rect 395337 300522 395403 300525
rect 510838 300522 510844 300524
rect 395337 300520 510844 300522
rect 395337 300464 395342 300520
rect 395398 300464 510844 300520
rect 395337 300462 510844 300464
rect 395337 300459 395403 300462
rect 510838 300460 510844 300462
rect 510908 300460 510914 300524
rect 395705 300386 395771 300389
rect 514334 300386 514340 300388
rect 395705 300384 514340 300386
rect 395705 300328 395710 300384
rect 395766 300328 514340 300384
rect 395705 300326 514340 300328
rect 395705 300323 395771 300326
rect 514334 300324 514340 300326
rect 514404 300324 514410 300388
rect 395521 300250 395587 300253
rect 514702 300250 514708 300252
rect 395521 300248 514708 300250
rect 395521 300192 395526 300248
rect 395582 300192 514708 300248
rect 395521 300190 514708 300192
rect 395521 300187 395587 300190
rect 514702 300188 514708 300190
rect 514772 300188 514778 300252
rect 392577 300114 392643 300117
rect 514886 300114 514892 300116
rect 392577 300112 514892 300114
rect 392577 300056 392582 300112
rect 392638 300056 514892 300112
rect 392577 300054 514892 300056
rect 392577 300051 392643 300054
rect 514886 300052 514892 300054
rect 514956 300052 514962 300116
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 389817 297394 389883 297397
rect 514150 297394 514156 297396
rect 389817 297392 514156 297394
rect 389817 297336 389822 297392
rect 389878 297336 514156 297392
rect 389817 297334 514156 297336
rect 389817 297331 389883 297334
rect 514150 297332 514156 297334
rect 514220 297332 514226 297396
rect 381629 294810 381695 294813
rect 511022 294810 511028 294812
rect 381629 294808 511028 294810
rect 381629 294752 381634 294808
rect 381690 294752 511028 294808
rect 381629 294750 511028 294752
rect 381629 294747 381695 294750
rect 511022 294748 511028 294750
rect 511092 294748 511098 294812
rect 381813 294674 381879 294677
rect 518014 294674 518020 294676
rect 381813 294672 518020 294674
rect 381813 294616 381818 294672
rect 381874 294616 518020 294672
rect 381813 294614 518020 294616
rect 381813 294611 381879 294614
rect 518014 294612 518020 294614
rect 518084 294612 518090 294676
rect 378777 294538 378843 294541
rect 516174 294538 516180 294540
rect 378777 294536 516180 294538
rect 378777 294480 378782 294536
rect 378838 294480 516180 294536
rect 378777 294478 516180 294480
rect 378777 294475 378843 294478
rect 516174 294476 516180 294478
rect 516244 294476 516250 294540
rect 361757 293450 361823 293453
rect 359812 293448 361823 293450
rect 359812 293392 361762 293448
rect 361818 293392 361823 293448
rect 359812 293390 361823 293392
rect 361757 293387 361823 293390
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 376385 291818 376451 291821
rect 508446 291818 508452 291820
rect 376385 291816 508452 291818
rect 376385 291760 376390 291816
rect 376446 291760 508452 291816
rect 376385 291758 508452 291760
rect 376385 291755 376451 291758
rect 508446 291756 508452 291758
rect 508516 291756 508522 291820
rect 370865 289098 370931 289101
rect 517830 289098 517836 289100
rect 370865 289096 517836 289098
rect 370865 289040 370870 289096
rect 370926 289040 517836 289096
rect 370865 289038 517836 289040
rect 370865 289035 370931 289038
rect 517830 289036 517836 289038
rect 517900 289036 517906 289100
rect 583520 285276 584960 285516
rect 361757 282434 361823 282437
rect 359812 282432 361823 282434
rect 359812 282376 361762 282432
rect 361818 282376 361823 282432
rect 359812 282374 361823 282376
rect 361757 282371 361823 282374
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 361757 271418 361823 271421
rect 359812 271416 361823 271418
rect 359812 271360 361762 271416
rect 361818 271360 361823 271416
rect 359812 271358 361823 271360
rect 361757 271355 361823 271358
rect -960 267202 480 267292
rect 3601 267202 3667 267205
rect -960 267200 3667 267202
rect -960 267144 3606 267200
rect 3662 267144 3667 267200
rect -960 267142 3667 267144
rect -960 267052 480 267142
rect 3601 267139 3667 267142
rect 456793 262714 456859 262717
rect 456793 262712 460092 262714
rect 456793 262656 456798 262712
rect 456854 262656 460092 262712
rect 456793 262654 460092 262656
rect 456793 262651 456859 262654
rect 529289 261626 529355 261629
rect 529289 261624 529490 261626
rect 529289 261568 529294 261624
rect 529350 261568 529490 261624
rect 529289 261566 529490 261568
rect 529289 261563 529355 261566
rect 529430 261052 529490 261566
rect 361757 260402 361823 260405
rect 359812 260400 361823 260402
rect 359812 260344 361762 260400
rect 361818 260344 361823 260400
rect 359812 260342 361823 260344
rect 361757 260339 361823 260342
rect 580257 258906 580323 258909
rect 583520 258906 584960 258996
rect 580257 258904 584960 258906
rect 580257 258848 580262 258904
rect 580318 258848 584960 258904
rect 580257 258846 584960 258848
rect 580257 258843 580323 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 361757 249386 361823 249389
rect 359812 249384 361823 249386
rect 359812 249328 361762 249384
rect 361818 249328 361823 249384
rect 359812 249326 361823 249328
rect 361757 249323 361823 249326
rect 456793 248842 456859 248845
rect 456793 248840 460092 248842
rect 456793 248784 456798 248840
rect 456854 248784 460092 248840
rect 456793 248782 460092 248784
rect 456793 248779 456859 248782
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 531313 243674 531379 243677
rect 529828 243672 531379 243674
rect 529828 243616 531318 243672
rect 531374 243616 531379 243672
rect 529828 243614 531379 243616
rect 531313 243611 531379 243614
rect -960 241090 480 241180
rect 3693 241090 3759 241093
rect -960 241088 3759 241090
rect -960 241032 3698 241088
rect 3754 241032 3759 241088
rect -960 241030 3759 241032
rect -960 240940 480 241030
rect 3693 241027 3759 241030
rect 361757 238370 361823 238373
rect 359812 238368 361823 238370
rect 359812 238312 361762 238368
rect 361818 238312 361823 238368
rect 359812 238310 361823 238312
rect 361757 238307 361823 238310
rect 458081 234970 458147 234973
rect 458081 234968 460092 234970
rect 458081 234912 458086 234968
rect 458142 234912 460092 234968
rect 458081 234910 460092 234912
rect 458081 234907 458147 234910
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 361757 227354 361823 227357
rect 359812 227352 361823 227354
rect 359812 227296 361762 227352
rect 361818 227296 361823 227352
rect 359812 227294 361823 227296
rect 361757 227291 361823 227294
rect 530117 226266 530183 226269
rect 529828 226264 530183 226266
rect 529828 226208 530122 226264
rect 530178 226208 530183 226264
rect 529828 226206 530183 226208
rect 530117 226203 530183 226206
rect 456793 221098 456859 221101
rect 456793 221096 460092 221098
rect 456793 221040 456798 221096
rect 456854 221040 460092 221096
rect 456793 221038 460092 221040
rect 456793 221035 456859 221038
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 361573 216338 361639 216341
rect 359812 216336 361639 216338
rect 359812 216280 361578 216336
rect 361634 216280 361639 216336
rect 359812 216278 361639 216280
rect 361573 216275 361639 216278
rect -960 214978 480 215068
rect 3877 214978 3943 214981
rect -960 214976 3943 214978
rect -960 214920 3882 214976
rect 3938 214920 3943 214976
rect -960 214918 3943 214920
rect -960 214828 480 214918
rect 3877 214915 3943 214918
rect 529933 209266 529999 209269
rect 529798 209264 529999 209266
rect 529798 209208 529938 209264
rect 529994 209208 529999 209264
rect 529798 209206 529999 209208
rect 529798 208828 529858 209206
rect 529933 209203 529999 209206
rect 456885 207226 456951 207229
rect 458725 207226 458791 207229
rect 456885 207224 460092 207226
rect 456885 207168 456890 207224
rect 456946 207168 458730 207224
rect 458786 207168 460092 207224
rect 456885 207166 460092 207168
rect 456885 207163 456951 207166
rect 458725 207163 458791 207166
rect 578877 205730 578943 205733
rect 583520 205730 584960 205820
rect 578877 205728 584960 205730
rect 578877 205672 578882 205728
rect 578938 205672 584960 205728
rect 578877 205670 584960 205672
rect 578877 205667 578943 205670
rect 583520 205580 584960 205670
rect 361757 205322 361823 205325
rect 359812 205320 361823 205322
rect 359812 205264 361762 205320
rect 361818 205264 361823 205320
rect 359812 205262 361823 205264
rect 361757 205259 361823 205262
rect -960 201922 480 202012
rect 3785 201922 3851 201925
rect -960 201920 3851 201922
rect -960 201864 3790 201920
rect 3846 201864 3851 201920
rect -960 201862 3851 201864
rect -960 201772 480 201862
rect 3785 201859 3851 201862
rect 361665 194306 361731 194309
rect 359812 194304 361731 194306
rect 359812 194248 361670 194304
rect 361726 194248 361731 194304
rect 359812 194246 361731 194248
rect 361665 194243 361731 194246
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3969 188866 4035 188869
rect -960 188864 4035 188866
rect -960 188808 3974 188864
rect 4030 188808 4035 188864
rect -960 188806 4035 188808
rect -960 188716 480 188806
rect 3969 188803 4035 188806
rect 361665 183290 361731 183293
rect 359812 183288 361731 183290
rect 359812 183232 361670 183288
rect 361726 183232 361731 183288
rect 359812 183230 361731 183232
rect 361665 183227 361731 183230
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 361757 172274 361823 172277
rect 359812 172272 361823 172274
rect 359812 172216 361762 172272
rect 361818 172216 361823 172272
rect 359812 172214 361823 172216
rect 361757 172211 361823 172214
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 4061 162890 4127 162893
rect -960 162888 4127 162890
rect -960 162832 4066 162888
rect 4122 162832 4127 162888
rect -960 162830 4127 162832
rect -960 162740 480 162830
rect 4061 162827 4127 162830
rect 421046 162692 421052 162756
rect 421116 162754 421122 162756
rect 421373 162754 421439 162757
rect 421116 162752 421439 162754
rect 421116 162696 421378 162752
rect 421434 162696 421439 162752
rect 421116 162694 421439 162696
rect 421116 162692 421122 162694
rect 421373 162691 421439 162694
rect 425830 162692 425836 162756
rect 425900 162754 425906 162756
rect 426157 162754 426223 162757
rect 425900 162752 426223 162754
rect 425900 162696 426162 162752
rect 426218 162696 426223 162752
rect 425900 162694 426223 162696
rect 425900 162692 425906 162694
rect 426157 162691 426223 162694
rect 428406 162692 428412 162756
rect 428476 162754 428482 162756
rect 428641 162754 428707 162757
rect 428476 162752 428707 162754
rect 428476 162696 428646 162752
rect 428702 162696 428707 162752
rect 428476 162694 428707 162696
rect 428476 162692 428482 162694
rect 428641 162691 428707 162694
rect 361757 161258 361823 161261
rect 359812 161256 361823 161258
rect 359812 161200 361762 161256
rect 361818 161200 361823 161256
rect 359812 161198 361823 161200
rect 361757 161195 361823 161198
rect 451733 158266 451799 158269
rect 449788 158264 451799 158266
rect 449788 158208 451738 158264
rect 451794 158208 451799 158264
rect 449788 158206 451799 158208
rect 451733 158203 451799 158206
rect 452561 156906 452627 156909
rect 449788 156904 452627 156906
rect 449788 156848 452566 156904
rect 452622 156848 452627 156904
rect 449788 156846 452627 156848
rect 452561 156843 452627 156846
rect 452101 155546 452167 155549
rect 449788 155544 452167 155546
rect 449788 155488 452106 155544
rect 452162 155488 452167 155544
rect 449788 155486 452167 155488
rect 452101 155483 452167 155486
rect 452193 154186 452259 154189
rect 449788 154184 452259 154186
rect 449788 154128 452198 154184
rect 452254 154128 452259 154184
rect 449788 154126 452259 154128
rect 452193 154123 452259 154126
rect 452101 152826 452167 152829
rect 449788 152824 452167 152826
rect 449788 152768 452106 152824
rect 452162 152768 452167 152824
rect 449788 152766 452167 152768
rect 452101 152763 452167 152766
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 452561 151466 452627 151469
rect 449788 151464 452627 151466
rect 449788 151408 452566 151464
rect 452622 151408 452627 151464
rect 449788 151406 452627 151408
rect 452561 151403 452627 151406
rect 362401 150242 362467 150245
rect 359812 150240 362467 150242
rect 359812 150184 362406 150240
rect 362462 150184 362467 150240
rect 359812 150182 362467 150184
rect 362401 150179 362467 150182
rect 452469 150106 452535 150109
rect 449788 150104 452535 150106
rect 449788 150048 452474 150104
rect 452530 150048 452535 150104
rect 449788 150046 452535 150048
rect 452469 150043 452535 150046
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 452009 148746 452075 148749
rect 449788 148744 452075 148746
rect 449788 148688 452014 148744
rect 452070 148688 452075 148744
rect 449788 148686 452075 148688
rect 452009 148683 452075 148686
rect 452561 147386 452627 147389
rect 449788 147384 452627 147386
rect 449788 147328 452566 147384
rect 452622 147328 452627 147384
rect 449788 147326 452627 147328
rect 452561 147323 452627 147326
rect 452561 146026 452627 146029
rect 449788 146024 452627 146026
rect 449788 145968 452566 146024
rect 452622 145968 452627 146024
rect 449788 145966 452627 145968
rect 452561 145963 452627 145966
rect 452561 144666 452627 144669
rect 449788 144664 452627 144666
rect 449788 144608 452566 144664
rect 452622 144608 452627 144664
rect 449788 144606 452627 144608
rect 452561 144603 452627 144606
rect 452561 143306 452627 143309
rect 449788 143304 452627 143306
rect 449788 143248 452566 143304
rect 452622 143248 452627 143304
rect 449788 143246 452627 143248
rect 452561 143243 452627 143246
rect 452561 141946 452627 141949
rect 449788 141944 452627 141946
rect 449788 141888 452566 141944
rect 452622 141888 452627 141944
rect 449788 141886 452627 141888
rect 452561 141883 452627 141886
rect 452101 140586 452167 140589
rect 449788 140584 452167 140586
rect 449788 140528 452106 140584
rect 452162 140528 452167 140584
rect 449788 140526 452167 140528
rect 452101 140523 452167 140526
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 361757 139226 361823 139229
rect 452561 139226 452627 139229
rect 359812 139224 361823 139226
rect 359812 139168 361762 139224
rect 361818 139168 361823 139224
rect 359812 139166 361823 139168
rect 449788 139224 452627 139226
rect 449788 139168 452566 139224
rect 452622 139168 452627 139224
rect 583520 139212 584960 139302
rect 449788 139166 452627 139168
rect 361757 139163 361823 139166
rect 452561 139163 452627 139166
rect 452561 137866 452627 137869
rect 449788 137864 452627 137866
rect 449788 137808 452566 137864
rect 452622 137808 452627 137864
rect 449788 137806 452627 137808
rect 452561 137803 452627 137806
rect 538806 137804 538812 137868
rect 538876 137866 538882 137868
rect 543273 137866 543339 137869
rect 538876 137864 543339 137866
rect 538876 137808 543278 137864
rect 543334 137808 543339 137864
rect 538876 137806 543339 137808
rect 538876 137804 538882 137806
rect 543273 137803 543339 137806
rect 539317 137730 539383 137733
rect 539317 137728 539426 137730
rect 539317 137672 539322 137728
rect 539378 137672 539426 137728
rect 539317 137667 539426 137672
rect 539366 137428 539426 137667
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 452561 136506 452627 136509
rect 449788 136504 452627 136506
rect 449788 136448 452566 136504
rect 452622 136448 452627 136504
rect 449788 136446 452627 136448
rect 452561 136443 452627 136446
rect 539501 135962 539567 135965
rect 539501 135960 539610 135962
rect 539501 135904 539506 135960
rect 539562 135904 539610 135960
rect 539501 135899 539610 135904
rect 539550 135388 539610 135899
rect 452561 135146 452627 135149
rect 449788 135144 452627 135146
rect 449788 135088 452566 135144
rect 452622 135088 452627 135144
rect 449788 135086 452627 135088
rect 452561 135083 452627 135086
rect 452469 133786 452535 133789
rect 449788 133784 452535 133786
rect 449788 133728 452474 133784
rect 452530 133728 452535 133784
rect 449788 133726 452535 133728
rect 452469 133723 452535 133726
rect 542721 133378 542787 133381
rect 539948 133376 542787 133378
rect 539948 133320 542726 133376
rect 542782 133320 542787 133376
rect 539948 133318 542787 133320
rect 542721 133315 542787 133318
rect 452101 132426 452167 132429
rect 449788 132424 452167 132426
rect 449788 132368 452106 132424
rect 452162 132368 452167 132424
rect 449788 132366 452167 132368
rect 452101 132363 452167 132366
rect 543181 131338 543247 131341
rect 539948 131336 543247 131338
rect 539948 131280 543186 131336
rect 543242 131280 543247 131336
rect 539948 131278 543247 131280
rect 543181 131275 543247 131278
rect 452561 131066 452627 131069
rect 449788 131064 452627 131066
rect 449788 131008 452566 131064
rect 452622 131008 452627 131064
rect 449788 131006 452627 131008
rect 452561 131003 452627 131006
rect 452377 129706 452443 129709
rect 449788 129704 452443 129706
rect 449788 129648 452382 129704
rect 452438 129648 452443 129704
rect 449788 129646 452443 129648
rect 452377 129643 452443 129646
rect 543089 129298 543155 129301
rect 539948 129296 543155 129298
rect 539948 129240 543094 129296
rect 543150 129240 543155 129296
rect 539948 129238 543155 129240
rect 543089 129235 543155 129238
rect 452285 128346 452351 128349
rect 449788 128344 452351 128346
rect 449788 128288 452290 128344
rect 452346 128288 452351 128344
rect 449788 128286 452351 128288
rect 452285 128283 452351 128286
rect 361573 128210 361639 128213
rect 359812 128208 361639 128210
rect 359812 128152 361578 128208
rect 361634 128152 361639 128208
rect 359812 128150 361639 128152
rect 361573 128147 361639 128150
rect 543273 127258 543339 127261
rect 539948 127256 543339 127258
rect 539948 127200 543278 127256
rect 543334 127200 543339 127256
rect 539948 127198 543339 127200
rect 543273 127195 543339 127198
rect 452193 126986 452259 126989
rect 449788 126984 452259 126986
rect 449788 126928 452198 126984
rect 452254 126928 452259 126984
rect 449788 126926 452259 126928
rect 452193 126923 452259 126926
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 451917 125626 451983 125629
rect 449788 125624 451983 125626
rect 449788 125568 451922 125624
rect 451978 125568 451983 125624
rect 449788 125566 451983 125568
rect 451917 125563 451983 125566
rect 542997 125218 543063 125221
rect 539948 125216 543063 125218
rect 539948 125160 543002 125216
rect 543058 125160 543063 125216
rect 539948 125158 543063 125160
rect 542997 125155 543063 125158
rect 451733 124266 451799 124269
rect 449788 124264 451799 124266
rect 449788 124208 451738 124264
rect 451794 124208 451799 124264
rect 449788 124206 451799 124208
rect 451733 124203 451799 124206
rect -960 123572 480 123812
rect 540329 123178 540395 123181
rect 539948 123176 540395 123178
rect 539948 123120 540334 123176
rect 540390 123120 540395 123176
rect 539948 123118 540395 123120
rect 540329 123115 540395 123118
rect 451733 122906 451799 122909
rect 449788 122904 451799 122906
rect 449788 122848 451738 122904
rect 451794 122848 451799 122904
rect 449788 122846 451799 122848
rect 451733 122843 451799 122846
rect 451733 121546 451799 121549
rect 449788 121544 451799 121546
rect 449788 121488 451738 121544
rect 451794 121488 451799 121544
rect 449788 121486 451799 121488
rect 451733 121483 451799 121486
rect 540237 121138 540303 121141
rect 539948 121136 540303 121138
rect 539948 121080 540242 121136
rect 540298 121080 540303 121136
rect 539948 121078 540303 121080
rect 540237 121075 540303 121078
rect 541065 119098 541131 119101
rect 539948 119096 541131 119098
rect 539948 119040 541070 119096
rect 541126 119040 541131 119096
rect 539948 119038 541131 119040
rect 541065 119035 541131 119038
rect 361573 117194 361639 117197
rect 359812 117192 361639 117194
rect 359812 117136 361578 117192
rect 361634 117136 361639 117192
rect 359812 117134 361639 117136
rect 361573 117131 361639 117134
rect 541525 117058 541591 117061
rect 539948 117056 541591 117058
rect 539948 117000 541530 117056
rect 541586 117000 541591 117056
rect 539948 116998 541591 117000
rect 541525 116995 541591 116998
rect 540145 115018 540211 115021
rect 539948 115016 540211 115018
rect 539948 114960 540150 115016
rect 540206 114960 540211 115016
rect 539948 114958 540211 114960
rect 540145 114955 540211 114958
rect 539685 113250 539751 113253
rect 539685 113248 539794 113250
rect 539685 113192 539690 113248
rect 539746 113192 539794 113248
rect 539685 113187 539794 113192
rect 539734 112948 539794 113187
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 541433 110938 541499 110941
rect 539948 110936 541499 110938
rect 539948 110880 541438 110936
rect 541494 110880 541499 110936
rect 539948 110878 541499 110880
rect 541433 110875 541499 110878
rect -960 110666 480 110756
rect 3366 110666 3372 110668
rect -960 110606 3372 110666
rect -960 110516 480 110606
rect 3366 110604 3372 110606
rect 3436 110604 3442 110668
rect 539918 108765 539978 108868
rect 539918 108760 540027 108765
rect 539918 108704 539966 108760
rect 540022 108704 540027 108760
rect 539918 108702 540027 108704
rect 539961 108699 540027 108702
rect 541341 106858 541407 106861
rect 539948 106856 541407 106858
rect 539948 106800 541346 106856
rect 541402 106800 541407 106856
rect 539948 106798 541407 106800
rect 541341 106795 541407 106798
rect 361573 106178 361639 106181
rect 359812 106176 361639 106178
rect 359812 106120 361578 106176
rect 361634 106120 361639 106176
rect 359812 106118 361639 106120
rect 361573 106115 361639 106118
rect 539918 104682 539978 104788
rect 540053 104682 540119 104685
rect 539918 104680 540119 104682
rect 539918 104624 540058 104680
rect 540114 104624 540119 104680
rect 539918 104622 540119 104624
rect 540053 104619 540119 104622
rect 541249 102778 541315 102781
rect 539948 102776 541315 102778
rect 539948 102720 541254 102776
rect 541310 102720 541315 102776
rect 539948 102718 541315 102720
rect 541249 102715 541315 102718
rect 542445 100738 542511 100741
rect 539948 100736 542511 100738
rect 539948 100680 542450 100736
rect 542506 100680 542511 100736
rect 539948 100678 542511 100680
rect 542445 100675 542511 100678
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 539869 99242 539935 99245
rect 539869 99240 539978 99242
rect 539869 99184 539874 99240
rect 539930 99184 539978 99240
rect 539869 99179 539978 99184
rect 539918 98668 539978 99179
rect -960 97610 480 97700
rect 3550 97610 3556 97612
rect -960 97550 3556 97610
rect -960 97460 480 97550
rect 3550 97548 3556 97550
rect 3620 97548 3626 97612
rect 542537 96658 542603 96661
rect 539948 96656 542603 96658
rect 539948 96600 542542 96656
rect 542598 96600 542603 96656
rect 539948 96598 542603 96600
rect 542537 96595 542603 96598
rect 361757 95162 361823 95165
rect 359812 95160 361823 95162
rect 359812 95104 361762 95160
rect 361818 95104 361823 95160
rect 359812 95102 361823 95104
rect 361757 95099 361823 95102
rect 542813 94618 542879 94621
rect 539948 94616 542879 94618
rect 539948 94560 542818 94616
rect 542874 94560 542879 94616
rect 539948 94558 542879 94560
rect 542813 94555 542879 94558
rect 541157 92578 541223 92581
rect 539948 92576 541223 92578
rect 539948 92520 541162 92576
rect 541218 92520 541223 92576
rect 539948 92518 541223 92520
rect 541157 92515 541223 92518
rect 542629 90538 542695 90541
rect 539948 90536 542695 90538
rect 539948 90480 542634 90536
rect 542690 90480 542695 90536
rect 539948 90478 542695 90480
rect 542629 90475 542695 90478
rect 542905 88498 542971 88501
rect 539948 88496 542971 88498
rect 539948 88440 542910 88496
rect 542966 88440 542971 88496
rect 539948 88438 542971 88440
rect 542905 88435 542971 88438
rect 539593 86866 539659 86869
rect 539550 86864 539659 86866
rect 539550 86808 539598 86864
rect 539654 86808 539659 86864
rect 539550 86803 539659 86808
rect 539550 86428 539610 86803
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3734 84690 3740 84692
rect -960 84630 3740 84690
rect -960 84540 480 84630
rect 3734 84628 3740 84630
rect 3804 84628 3810 84692
rect 542670 84418 542676 84420
rect 539948 84358 542676 84418
rect 542670 84356 542676 84358
rect 542740 84356 542746 84420
rect 361757 84146 361823 84149
rect 359812 84144 361823 84146
rect 359812 84088 361762 84144
rect 361818 84088 361823 84144
rect 359812 84086 361823 84088
rect 361757 84083 361823 84086
rect 540973 82378 541039 82381
rect 539948 82376 541039 82378
rect 539948 82320 540978 82376
rect 541034 82320 541039 82376
rect 539948 82318 541039 82320
rect 540973 82315 541039 82318
rect 361757 73130 361823 73133
rect 359812 73128 361823 73130
rect 359812 73072 361762 73128
rect 361818 73072 361823 73128
rect 359812 73070 361823 73072
rect 361757 73067 361823 73070
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 361757 62114 361823 62117
rect 359812 62112 361823 62114
rect 359812 62056 361762 62112
rect 361818 62056 361823 62112
rect 359812 62054 361823 62056
rect 361757 62051 361823 62054
rect 20897 59938 20963 59941
rect 21449 59938 21515 59941
rect 20897 59936 21515 59938
rect 20897 59880 20902 59936
rect 20958 59880 21454 59936
rect 21510 59880 21515 59936
rect 20897 59878 21515 59880
rect 20897 59875 20963 59878
rect 21449 59875 21515 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 361757 51098 361823 51101
rect 359812 51096 361823 51098
rect 359812 51040 361762 51096
rect 361818 51040 361823 51096
rect 359812 51038 361823 51040
rect 361757 51035 361823 51038
rect 19333 49602 19399 49605
rect 22134 49602 22140 49604
rect 19333 49600 22140 49602
rect 19333 49544 19338 49600
rect 19394 49544 22140 49600
rect 19333 49542 22140 49544
rect 19333 49539 19399 49542
rect 22134 49540 22140 49542
rect 22204 49540 22210 49604
rect 20897 49466 20963 49469
rect 22318 49466 22324 49468
rect 20897 49464 22324 49466
rect 20897 49408 20902 49464
rect 20958 49408 22324 49464
rect 20897 49406 22324 49408
rect 20897 49403 20963 49406
rect 22318 49404 22324 49406
rect 22388 49404 22394 49468
rect 540605 48922 540671 48925
rect 540605 48920 540714 48922
rect 540605 48864 540610 48920
rect 540666 48864 540714 48920
rect 540605 48859 540714 48864
rect 540654 48348 540714 48859
rect 3366 46820 3372 46884
rect 3436 46882 3442 46884
rect 458909 46882 458975 46885
rect 3436 46880 458975 46882
rect 3436 46824 458914 46880
rect 458970 46824 458975 46880
rect 3436 46822 458975 46824
rect 3436 46820 3442 46822
rect 458909 46819 458975 46822
rect 3550 46684 3556 46748
rect 3620 46746 3626 46748
rect 459093 46746 459159 46749
rect 3620 46744 459159 46746
rect 3620 46688 459098 46744
rect 459154 46688 459159 46744
rect 3620 46686 459159 46688
rect 3620 46684 3626 46686
rect 459093 46683 459159 46686
rect 3734 46548 3740 46612
rect 3804 46610 3810 46612
rect 456149 46610 456215 46613
rect 3804 46608 456215 46610
rect 3804 46552 456154 46608
rect 456210 46552 456215 46608
rect 3804 46550 456215 46552
rect 3804 46548 3810 46550
rect 456149 46547 456215 46550
rect 22134 46412 22140 46476
rect 22204 46474 22210 46476
rect 361205 46474 361271 46477
rect 22204 46472 361271 46474
rect 22204 46416 361210 46472
rect 361266 46416 361271 46472
rect 22204 46414 361271 46416
rect 22204 46412 22210 46414
rect 361205 46411 361271 46414
rect 22318 46276 22324 46340
rect 22388 46338 22394 46340
rect 359641 46338 359707 46341
rect 22388 46336 359707 46338
rect 22388 46280 359646 46336
rect 359702 46280 359707 46336
rect 22388 46278 359707 46280
rect 22388 46276 22394 46278
rect 359641 46275 359707 46278
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 27613 44978 27679 44981
rect 368197 44978 368263 44981
rect 27613 44976 368263 44978
rect 27613 44920 27618 44976
rect 27674 44920 368202 44976
rect 368258 44920 368263 44976
rect 27613 44918 368263 44920
rect 27613 44915 27679 44918
rect 368197 44915 368263 44918
rect 6913 44842 6979 44845
rect 409229 44842 409295 44845
rect 6913 44840 409295 44842
rect 6913 44784 6918 44840
rect 6974 44784 409234 44840
rect 409290 44784 409295 44840
rect 6913 44782 409295 44784
rect 6913 44779 6979 44782
rect 409229 44779 409295 44782
rect 537477 41034 537543 41037
rect 537477 41032 540132 41034
rect 537477 40976 537482 41032
rect 537538 40976 540132 41032
rect 537477 40974 540132 40976
rect 537477 40971 537543 40974
rect 121453 39402 121519 39405
rect 458766 39402 458772 39404
rect 121453 39400 458772 39402
rect 121453 39344 121458 39400
rect 121514 39344 458772 39400
rect 121453 39342 458772 39344
rect 121453 39339 121519 39342
rect 458766 39340 458772 39342
rect 458836 39340 458842 39404
rect 26233 39266 26299 39269
rect 458950 39266 458956 39268
rect 26233 39264 458956 39266
rect 26233 39208 26238 39264
rect 26294 39208 458956 39264
rect 26233 39206 458956 39208
rect 26233 39203 26299 39206
rect 458950 39204 458956 39206
rect 459020 39204 459026 39268
rect 539777 33690 539843 33693
rect 539777 33688 540132 33690
rect 539777 33632 539782 33688
rect 539838 33632 540132 33688
rect 539777 33630 540132 33632
rect 539777 33627 539843 33630
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 5257 3906 5323 3909
rect 362217 3906 362283 3909
rect 5257 3904 362283 3906
rect 5257 3848 5262 3904
rect 5318 3848 362222 3904
rect 362278 3848 362283 3904
rect 5257 3846 362283 3848
rect 5257 3843 5323 3846
rect 362217 3843 362283 3846
rect 6453 3770 6519 3773
rect 367737 3770 367803 3773
rect 6453 3768 367803 3770
rect 6453 3712 6458 3768
rect 6514 3712 367742 3768
rect 367798 3712 367803 3768
rect 6453 3710 367803 3712
rect 6453 3707 6519 3710
rect 367737 3707 367803 3710
rect 8753 3634 8819 3637
rect 392577 3634 392643 3637
rect 8753 3632 392643 3634
rect 8753 3576 8758 3632
rect 8814 3576 392582 3632
rect 392638 3576 392643 3632
rect 8753 3574 392643 3576
rect 8753 3571 8819 3574
rect 392577 3571 392643 3574
rect 1669 3498 1735 3501
rect 450721 3498 450787 3501
rect 1669 3496 450787 3498
rect 1669 3440 1674 3496
rect 1730 3440 450726 3496
rect 450782 3440 450787 3496
rect 1669 3438 450787 3440
rect 1669 3435 1735 3438
rect 450721 3435 450787 3438
rect 565 3362 631 3365
rect 454677 3362 454743 3365
rect 565 3360 454743 3362
rect 565 3304 570 3360
rect 626 3304 454682 3360
rect 454738 3304 454743 3360
rect 565 3302 454743 3304
rect 565 3299 631 3302
rect 454677 3299 454743 3302
<< via3 >>
rect 449572 700436 449636 700500
rect 451780 700436 451844 700500
rect 447732 700300 447796 700364
rect 455092 700300 455156 700364
rect 527220 699816 527284 699820
rect 527220 699760 527234 699816
rect 527234 699760 527284 699816
rect 527220 699756 527284 699760
rect 556292 699756 556356 699820
rect 450492 692004 450556 692068
rect 444236 690644 444300 690708
rect 450676 689284 450740 689348
rect 22692 684524 22756 684588
rect 3556 683300 3620 683364
rect 3740 683164 3804 683228
rect 3372 682756 3436 682820
rect 22692 669836 22756 669900
rect 453252 669836 453316 669900
rect 458036 665484 458100 665548
rect 457852 663036 457916 663100
rect 3740 658140 3804 658204
rect 458956 636108 459020 636172
rect 459140 633660 459204 633724
rect 3556 619108 3620 619172
rect 3372 606052 3436 606116
rect 478828 599524 478892 599588
rect 474412 598164 474476 598228
rect 474780 596940 474844 597004
rect 476436 596804 476500 596868
rect 472020 522276 472084 522340
rect 457852 519420 457916 519484
rect 458036 517516 458100 517580
rect 448284 516156 448348 516220
rect 483060 496844 483124 496908
rect 486372 496904 486436 496908
rect 486372 496848 486422 496904
rect 486422 496848 486436 496904
rect 486372 496844 486436 496848
rect 448284 496028 448348 496092
rect 527220 465700 527284 465764
rect 487108 453868 487172 453932
rect 455092 422860 455156 422924
rect 444052 421908 444116 421972
rect 451780 420140 451844 420204
rect 458956 393892 459020 393956
rect 459140 392532 459204 392596
rect 472020 388996 472084 389060
rect 474412 389056 474476 389060
rect 474412 389000 474426 389056
rect 474426 389000 474476 389056
rect 474412 388996 474476 389000
rect 474780 388996 474844 389060
rect 476436 388996 476500 389060
rect 478828 388996 478892 389060
rect 453252 387636 453316 387700
rect 483060 387092 483124 387156
rect 486372 386956 486436 387020
rect 487108 385596 487172 385660
rect 425836 335412 425900 335476
rect 518020 335140 518084 335204
rect 421052 334460 421116 334524
rect 428412 334460 428476 334524
rect 511028 333508 511092 333572
rect 425836 332964 425900 333028
rect 515076 332964 515140 333028
rect 514708 331332 514772 331396
rect 517836 330788 517900 330852
rect 510844 329700 510908 329764
rect 448284 329156 448348 329220
rect 514156 328612 514220 328676
rect 510476 328068 510540 328132
rect 516180 327524 516244 327588
rect 514892 326980 514956 327044
rect 510660 326436 510724 326500
rect 514340 324804 514404 324868
rect 510660 324396 510724 324460
rect 511212 324396 511276 324460
rect 510660 324260 510724 324324
rect 508452 322764 508516 322828
rect 509188 322628 509252 322692
rect 447732 321812 447796 321876
rect 556292 321404 556356 321468
rect 449572 321268 449636 321332
rect 444052 321132 444116 321196
rect 450676 319908 450740 319972
rect 444236 319772 444300 319836
rect 450492 319500 450556 319564
rect 538812 319364 538876 319428
rect 511212 317188 511276 317252
rect 458956 317052 459020 317116
rect 515076 317052 515140 317116
rect 510660 316916 510724 316980
rect 458772 316780 458836 316844
rect 509004 316644 509068 316708
rect 542676 315284 542740 315348
rect 510476 302772 510540 302836
rect 510844 300460 510908 300524
rect 514340 300324 514404 300388
rect 514708 300188 514772 300252
rect 514892 300052 514956 300116
rect 514156 297332 514220 297396
rect 511028 294748 511092 294812
rect 518020 294612 518084 294676
rect 516180 294476 516244 294540
rect 508452 291756 508516 291820
rect 517836 289036 517900 289100
rect 421052 162692 421116 162756
rect 425836 162692 425900 162756
rect 428412 162692 428476 162756
rect 538812 137804 538876 137868
rect 3372 110604 3436 110668
rect 3556 97548 3620 97612
rect 3740 84628 3804 84692
rect 542676 84356 542740 84420
rect 22140 49540 22204 49604
rect 22324 49404 22388 49468
rect 3372 46820 3436 46884
rect 3556 46684 3620 46748
rect 3740 46548 3804 46612
rect 22140 46412 22204 46476
rect 22324 46276 22388 46340
rect 458772 39340 458836 39404
rect 458956 39204 459020 39268
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 3555 683364 3621 683365
rect 3555 683300 3556 683364
rect 3620 683300 3621 683364
rect 3555 683299 3621 683300
rect 3371 682820 3437 682821
rect 3371 682756 3372 682820
rect 3436 682756 3437 682820
rect 3371 682755 3437 682756
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 3374 606117 3434 682755
rect 3558 619173 3618 683299
rect 3739 683228 3805 683229
rect 3739 683164 3740 683228
rect 3804 683164 3805 683228
rect 3739 683163 3805 683164
rect 3742 658205 3802 683163
rect 3739 658204 3805 658205
rect 3739 658140 3740 658204
rect 3804 658140 3805 658204
rect 3739 658139 3805 658140
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3555 619172 3621 619173
rect 3555 619108 3556 619172
rect 3620 619108 3621 619172
rect 3555 619107 3621 619108
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 3374 46885 3434 110603
rect 3555 97612 3621 97613
rect 3555 97548 3556 97612
rect 3620 97548 3621 97612
rect 3555 97547 3621 97548
rect 3371 46884 3437 46885
rect 3371 46820 3372 46884
rect 3436 46820 3437 46884
rect 3371 46819 3437 46820
rect 3558 46749 3618 97547
rect 3739 84692 3805 84693
rect 3739 84628 3740 84692
rect 3804 84628 3805 84692
rect 3739 84627 3805 84628
rect 3555 46748 3621 46749
rect 3555 46684 3556 46748
rect 3620 46684 3621 46748
rect 3555 46683 3621 46684
rect 3742 46613 3802 84627
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3739 46612 3805 46613
rect 3739 46548 3740 46612
rect 3804 46548 3805 46612
rect 3739 46547 3805 46548
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 22691 684588 22757 684589
rect 22691 684524 22692 684588
rect 22756 684524 22757 684588
rect 22691 684523 22757 684524
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 22694 669901 22754 684523
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 22691 669900 22757 669901
rect 22691 669836 22692 669900
rect 22756 669836 22757 669900
rect 22691 669835 22757 669836
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 24208 651454 24528 651486
rect 24208 651218 24250 651454
rect 24486 651218 24528 651454
rect 24208 651134 24528 651218
rect 24208 650898 24250 651134
rect 24486 650898 24528 651134
rect 24208 650866 24528 650898
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 674393 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 674393 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 674393 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 674393 49574 698058
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 674393 64454 676938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 674393 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 674393 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 674393 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 674393 85574 698058
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 674393 100454 676938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 674393 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 674393 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 674393 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 674393 121574 698058
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 674393 136454 676938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 674393 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 674393 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 674393 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 674393 157574 698058
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 674393 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 674393 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 674393 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 674393 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 684676 193574 698058
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 674393 208454 676938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 674393 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 674393 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 674393 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 674393 229574 698058
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 674393 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 674393 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 674393 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 674393 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 674393 265574 698058
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 674393 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 674393 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 674393 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 674393 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 684676 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 674393 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 674393 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 674393 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 674393 337574 698058
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 674393 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 39568 655174 39888 655206
rect 39568 654938 39610 655174
rect 39846 654938 39888 655174
rect 39568 654854 39888 654938
rect 39568 654618 39610 654854
rect 39846 654618 39888 654854
rect 39568 654586 39888 654618
rect 70288 655174 70608 655206
rect 70288 654938 70330 655174
rect 70566 654938 70608 655174
rect 70288 654854 70608 654938
rect 70288 654618 70330 654854
rect 70566 654618 70608 654854
rect 70288 654586 70608 654618
rect 101008 655174 101328 655206
rect 101008 654938 101050 655174
rect 101286 654938 101328 655174
rect 101008 654854 101328 654938
rect 101008 654618 101050 654854
rect 101286 654618 101328 654854
rect 101008 654586 101328 654618
rect 131728 655174 132048 655206
rect 131728 654938 131770 655174
rect 132006 654938 132048 655174
rect 131728 654854 132048 654938
rect 131728 654618 131770 654854
rect 132006 654618 132048 654854
rect 131728 654586 132048 654618
rect 162448 655174 162768 655206
rect 162448 654938 162490 655174
rect 162726 654938 162768 655174
rect 162448 654854 162768 654938
rect 162448 654618 162490 654854
rect 162726 654618 162768 654854
rect 162448 654586 162768 654618
rect 193168 655174 193488 655206
rect 193168 654938 193210 655174
rect 193446 654938 193488 655174
rect 193168 654854 193488 654938
rect 193168 654618 193210 654854
rect 193446 654618 193488 654854
rect 193168 654586 193488 654618
rect 223888 655174 224208 655206
rect 223888 654938 223930 655174
rect 224166 654938 224208 655174
rect 223888 654854 224208 654938
rect 223888 654618 223930 654854
rect 224166 654618 224208 654854
rect 223888 654586 224208 654618
rect 254608 655174 254928 655206
rect 254608 654938 254650 655174
rect 254886 654938 254928 655174
rect 254608 654854 254928 654938
rect 254608 654618 254650 654854
rect 254886 654618 254928 654854
rect 254608 654586 254928 654618
rect 285328 655174 285648 655206
rect 285328 654938 285370 655174
rect 285606 654938 285648 655174
rect 285328 654854 285648 654938
rect 285328 654618 285370 654854
rect 285606 654618 285648 654854
rect 285328 654586 285648 654618
rect 316048 655174 316368 655206
rect 316048 654938 316090 655174
rect 316326 654938 316368 655174
rect 316048 654854 316368 654938
rect 316048 654618 316090 654854
rect 316326 654618 316368 654854
rect 316048 654586 316368 654618
rect 346768 655174 347088 655206
rect 346768 654938 346810 655174
rect 347046 654938 347088 655174
rect 346768 654854 347088 654938
rect 346768 654618 346810 654854
rect 347046 654618 347088 654854
rect 346768 654586 347088 654618
rect 54928 651454 55248 651486
rect 54928 651218 54970 651454
rect 55206 651218 55248 651454
rect 54928 651134 55248 651218
rect 54928 650898 54970 651134
rect 55206 650898 55248 651134
rect 54928 650866 55248 650898
rect 85648 651454 85968 651486
rect 85648 651218 85690 651454
rect 85926 651218 85968 651454
rect 85648 651134 85968 651218
rect 85648 650898 85690 651134
rect 85926 650898 85968 651134
rect 85648 650866 85968 650898
rect 116368 651454 116688 651486
rect 116368 651218 116410 651454
rect 116646 651218 116688 651454
rect 116368 651134 116688 651218
rect 116368 650898 116410 651134
rect 116646 650898 116688 651134
rect 116368 650866 116688 650898
rect 147088 651454 147408 651486
rect 147088 651218 147130 651454
rect 147366 651218 147408 651454
rect 147088 651134 147408 651218
rect 147088 650898 147130 651134
rect 147366 650898 147408 651134
rect 147088 650866 147408 650898
rect 177808 651454 178128 651486
rect 177808 651218 177850 651454
rect 178086 651218 178128 651454
rect 177808 651134 178128 651218
rect 177808 650898 177850 651134
rect 178086 650898 178128 651134
rect 177808 650866 178128 650898
rect 208528 651454 208848 651486
rect 208528 651218 208570 651454
rect 208806 651218 208848 651454
rect 208528 651134 208848 651218
rect 208528 650898 208570 651134
rect 208806 650898 208848 651134
rect 208528 650866 208848 650898
rect 239248 651454 239568 651486
rect 239248 651218 239290 651454
rect 239526 651218 239568 651454
rect 239248 651134 239568 651218
rect 239248 650898 239290 651134
rect 239526 650898 239568 651134
rect 239248 650866 239568 650898
rect 269968 651454 270288 651486
rect 269968 651218 270010 651454
rect 270246 651218 270288 651454
rect 269968 651134 270288 651218
rect 269968 650898 270010 651134
rect 270246 650898 270288 651134
rect 269968 650866 270288 650898
rect 300688 651454 301008 651486
rect 300688 651218 300730 651454
rect 300966 651218 301008 651454
rect 300688 651134 301008 651218
rect 300688 650898 300730 651134
rect 300966 650898 301008 651134
rect 300688 650866 301008 650898
rect 331408 651454 331728 651486
rect 331408 651218 331450 651454
rect 331686 651218 331728 651454
rect 331408 651134 331728 651218
rect 331408 650898 331450 651134
rect 331686 650898 331728 651134
rect 331408 650866 331728 650898
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 24208 615454 24528 615486
rect 24208 615218 24250 615454
rect 24486 615218 24528 615454
rect 24208 615134 24528 615218
rect 24208 614898 24250 615134
rect 24486 614898 24528 615134
rect 24208 614866 24528 614898
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 27834 605494 28454 640938
rect 39568 619174 39888 619206
rect 39568 618938 39610 619174
rect 39846 618938 39888 619174
rect 39568 618854 39888 618938
rect 39568 618618 39610 618854
rect 39846 618618 39888 618854
rect 39568 618586 39888 618618
rect 70288 619174 70608 619206
rect 70288 618938 70330 619174
rect 70566 618938 70608 619174
rect 70288 618854 70608 618938
rect 70288 618618 70330 618854
rect 70566 618618 70608 618854
rect 70288 618586 70608 618618
rect 101008 619174 101328 619206
rect 101008 618938 101050 619174
rect 101286 618938 101328 619174
rect 101008 618854 101328 618938
rect 101008 618618 101050 618854
rect 101286 618618 101328 618854
rect 101008 618586 101328 618618
rect 131728 619174 132048 619206
rect 131728 618938 131770 619174
rect 132006 618938 132048 619174
rect 131728 618854 132048 618938
rect 131728 618618 131770 618854
rect 132006 618618 132048 618854
rect 131728 618586 132048 618618
rect 162448 619174 162768 619206
rect 162448 618938 162490 619174
rect 162726 618938 162768 619174
rect 162448 618854 162768 618938
rect 162448 618618 162490 618854
rect 162726 618618 162768 618854
rect 162448 618586 162768 618618
rect 193168 619174 193488 619206
rect 193168 618938 193210 619174
rect 193446 618938 193488 619174
rect 193168 618854 193488 618938
rect 193168 618618 193210 618854
rect 193446 618618 193488 618854
rect 193168 618586 193488 618618
rect 223888 619174 224208 619206
rect 223888 618938 223930 619174
rect 224166 618938 224208 619174
rect 223888 618854 224208 618938
rect 223888 618618 223930 618854
rect 224166 618618 224208 618854
rect 223888 618586 224208 618618
rect 254608 619174 254928 619206
rect 254608 618938 254650 619174
rect 254886 618938 254928 619174
rect 254608 618854 254928 618938
rect 254608 618618 254650 618854
rect 254886 618618 254928 618854
rect 254608 618586 254928 618618
rect 285328 619174 285648 619206
rect 285328 618938 285370 619174
rect 285606 618938 285648 619174
rect 285328 618854 285648 618938
rect 285328 618618 285370 618854
rect 285606 618618 285648 618854
rect 285328 618586 285648 618618
rect 316048 619174 316368 619206
rect 316048 618938 316090 619174
rect 316326 618938 316368 619174
rect 316048 618854 316368 618938
rect 316048 618618 316090 618854
rect 316326 618618 316368 618854
rect 316048 618586 316368 618618
rect 346768 619174 347088 619206
rect 346768 618938 346810 619174
rect 347046 618938 347088 619174
rect 346768 618854 347088 618938
rect 346768 618618 346810 618854
rect 347046 618618 347088 618854
rect 346768 618586 347088 618618
rect 54928 615454 55248 615486
rect 54928 615218 54970 615454
rect 55206 615218 55248 615454
rect 54928 615134 55248 615218
rect 54928 614898 54970 615134
rect 55206 614898 55248 615134
rect 54928 614866 55248 614898
rect 85648 615454 85968 615486
rect 85648 615218 85690 615454
rect 85926 615218 85968 615454
rect 85648 615134 85968 615218
rect 85648 614898 85690 615134
rect 85926 614898 85968 615134
rect 85648 614866 85968 614898
rect 116368 615454 116688 615486
rect 116368 615218 116410 615454
rect 116646 615218 116688 615454
rect 116368 615134 116688 615218
rect 116368 614898 116410 615134
rect 116646 614898 116688 615134
rect 116368 614866 116688 614898
rect 147088 615454 147408 615486
rect 147088 615218 147130 615454
rect 147366 615218 147408 615454
rect 147088 615134 147408 615218
rect 147088 614898 147130 615134
rect 147366 614898 147408 615134
rect 147088 614866 147408 614898
rect 177808 615454 178128 615486
rect 177808 615218 177850 615454
rect 178086 615218 178128 615454
rect 177808 615134 178128 615218
rect 177808 614898 177850 615134
rect 178086 614898 178128 615134
rect 177808 614866 178128 614898
rect 208528 615454 208848 615486
rect 208528 615218 208570 615454
rect 208806 615218 208848 615454
rect 208528 615134 208848 615218
rect 208528 614898 208570 615134
rect 208806 614898 208848 615134
rect 208528 614866 208848 614898
rect 239248 615454 239568 615486
rect 239248 615218 239290 615454
rect 239526 615218 239568 615454
rect 239248 615134 239568 615218
rect 239248 614898 239290 615134
rect 239526 614898 239568 615134
rect 239248 614866 239568 614898
rect 269968 615454 270288 615486
rect 269968 615218 270010 615454
rect 270246 615218 270288 615454
rect 269968 615134 270288 615218
rect 269968 614898 270010 615134
rect 270246 614898 270288 615134
rect 269968 614866 270288 614898
rect 300688 615454 301008 615486
rect 300688 615218 300730 615454
rect 300966 615218 301008 615454
rect 300688 615134 301008 615218
rect 300688 614898 300730 615134
rect 300966 614898 301008 615134
rect 300688 614866 301008 614898
rect 331408 615454 331728 615486
rect 331408 615218 331450 615454
rect 331686 615218 331728 615454
rect 331408 615134 331728 615218
rect 331408 614898 331450 615134
rect 331686 614898 331728 615134
rect 331408 614866 331728 614898
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 24208 579454 24528 579486
rect 24208 579218 24250 579454
rect 24486 579218 24528 579454
rect 24208 579134 24528 579218
rect 24208 578898 24250 579134
rect 24486 578898 24528 579134
rect 24208 578866 24528 578898
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 27834 569494 28454 604938
rect 39568 583174 39888 583206
rect 39568 582938 39610 583174
rect 39846 582938 39888 583174
rect 39568 582854 39888 582938
rect 39568 582618 39610 582854
rect 39846 582618 39888 582854
rect 39568 582586 39888 582618
rect 70288 583174 70608 583206
rect 70288 582938 70330 583174
rect 70566 582938 70608 583174
rect 70288 582854 70608 582938
rect 70288 582618 70330 582854
rect 70566 582618 70608 582854
rect 70288 582586 70608 582618
rect 101008 583174 101328 583206
rect 101008 582938 101050 583174
rect 101286 582938 101328 583174
rect 101008 582854 101328 582938
rect 101008 582618 101050 582854
rect 101286 582618 101328 582854
rect 101008 582586 101328 582618
rect 131728 583174 132048 583206
rect 131728 582938 131770 583174
rect 132006 582938 132048 583174
rect 131728 582854 132048 582938
rect 131728 582618 131770 582854
rect 132006 582618 132048 582854
rect 131728 582586 132048 582618
rect 162448 583174 162768 583206
rect 162448 582938 162490 583174
rect 162726 582938 162768 583174
rect 162448 582854 162768 582938
rect 162448 582618 162490 582854
rect 162726 582618 162768 582854
rect 162448 582586 162768 582618
rect 193168 583174 193488 583206
rect 193168 582938 193210 583174
rect 193446 582938 193488 583174
rect 193168 582854 193488 582938
rect 193168 582618 193210 582854
rect 193446 582618 193488 582854
rect 193168 582586 193488 582618
rect 223888 583174 224208 583206
rect 223888 582938 223930 583174
rect 224166 582938 224208 583174
rect 223888 582854 224208 582938
rect 223888 582618 223930 582854
rect 224166 582618 224208 582854
rect 223888 582586 224208 582618
rect 254608 583174 254928 583206
rect 254608 582938 254650 583174
rect 254886 582938 254928 583174
rect 254608 582854 254928 582938
rect 254608 582618 254650 582854
rect 254886 582618 254928 582854
rect 254608 582586 254928 582618
rect 285328 583174 285648 583206
rect 285328 582938 285370 583174
rect 285606 582938 285648 583174
rect 285328 582854 285648 582938
rect 285328 582618 285370 582854
rect 285606 582618 285648 582854
rect 285328 582586 285648 582618
rect 316048 583174 316368 583206
rect 316048 582938 316090 583174
rect 316326 582938 316368 583174
rect 316048 582854 316368 582938
rect 316048 582618 316090 582854
rect 316326 582618 316368 582854
rect 316048 582586 316368 582618
rect 346768 583174 347088 583206
rect 346768 582938 346810 583174
rect 347046 582938 347088 583174
rect 346768 582854 347088 582938
rect 346768 582618 346810 582854
rect 347046 582618 347088 582854
rect 346768 582586 347088 582618
rect 54928 579454 55248 579486
rect 54928 579218 54970 579454
rect 55206 579218 55248 579454
rect 54928 579134 55248 579218
rect 54928 578898 54970 579134
rect 55206 578898 55248 579134
rect 54928 578866 55248 578898
rect 85648 579454 85968 579486
rect 85648 579218 85690 579454
rect 85926 579218 85968 579454
rect 85648 579134 85968 579218
rect 85648 578898 85690 579134
rect 85926 578898 85968 579134
rect 85648 578866 85968 578898
rect 116368 579454 116688 579486
rect 116368 579218 116410 579454
rect 116646 579218 116688 579454
rect 116368 579134 116688 579218
rect 116368 578898 116410 579134
rect 116646 578898 116688 579134
rect 116368 578866 116688 578898
rect 147088 579454 147408 579486
rect 147088 579218 147130 579454
rect 147366 579218 147408 579454
rect 147088 579134 147408 579218
rect 147088 578898 147130 579134
rect 147366 578898 147408 579134
rect 147088 578866 147408 578898
rect 177808 579454 178128 579486
rect 177808 579218 177850 579454
rect 178086 579218 178128 579454
rect 177808 579134 178128 579218
rect 177808 578898 177850 579134
rect 178086 578898 178128 579134
rect 177808 578866 178128 578898
rect 208528 579454 208848 579486
rect 208528 579218 208570 579454
rect 208806 579218 208848 579454
rect 208528 579134 208848 579218
rect 208528 578898 208570 579134
rect 208806 578898 208848 579134
rect 208528 578866 208848 578898
rect 239248 579454 239568 579486
rect 239248 579218 239290 579454
rect 239526 579218 239568 579454
rect 239248 579134 239568 579218
rect 239248 578898 239290 579134
rect 239526 578898 239568 579134
rect 239248 578866 239568 578898
rect 269968 579454 270288 579486
rect 269968 579218 270010 579454
rect 270246 579218 270288 579454
rect 269968 579134 270288 579218
rect 269968 578898 270010 579134
rect 270246 578898 270288 579134
rect 269968 578866 270288 578898
rect 300688 579454 301008 579486
rect 300688 579218 300730 579454
rect 300966 579218 301008 579454
rect 300688 579134 301008 579218
rect 300688 578898 300730 579134
rect 300966 578898 301008 579134
rect 300688 578866 301008 578898
rect 331408 579454 331728 579486
rect 331408 579218 331450 579454
rect 331686 579218 331728 579454
rect 331408 579134 331728 579218
rect 331408 578898 331450 579134
rect 331686 578898 331728 579134
rect 331408 578866 331728 578898
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 24208 543454 24528 543486
rect 24208 543218 24250 543454
rect 24486 543218 24528 543454
rect 24208 543134 24528 543218
rect 24208 542898 24250 543134
rect 24486 542898 24528 543134
rect 24208 542866 24528 542898
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 27834 533494 28454 568938
rect 39568 547174 39888 547206
rect 39568 546938 39610 547174
rect 39846 546938 39888 547174
rect 39568 546854 39888 546938
rect 39568 546618 39610 546854
rect 39846 546618 39888 546854
rect 39568 546586 39888 546618
rect 70288 547174 70608 547206
rect 70288 546938 70330 547174
rect 70566 546938 70608 547174
rect 70288 546854 70608 546938
rect 70288 546618 70330 546854
rect 70566 546618 70608 546854
rect 70288 546586 70608 546618
rect 101008 547174 101328 547206
rect 101008 546938 101050 547174
rect 101286 546938 101328 547174
rect 101008 546854 101328 546938
rect 101008 546618 101050 546854
rect 101286 546618 101328 546854
rect 101008 546586 101328 546618
rect 131728 547174 132048 547206
rect 131728 546938 131770 547174
rect 132006 546938 132048 547174
rect 131728 546854 132048 546938
rect 131728 546618 131770 546854
rect 132006 546618 132048 546854
rect 131728 546586 132048 546618
rect 162448 547174 162768 547206
rect 162448 546938 162490 547174
rect 162726 546938 162768 547174
rect 162448 546854 162768 546938
rect 162448 546618 162490 546854
rect 162726 546618 162768 546854
rect 162448 546586 162768 546618
rect 193168 547174 193488 547206
rect 193168 546938 193210 547174
rect 193446 546938 193488 547174
rect 193168 546854 193488 546938
rect 193168 546618 193210 546854
rect 193446 546618 193488 546854
rect 193168 546586 193488 546618
rect 223888 547174 224208 547206
rect 223888 546938 223930 547174
rect 224166 546938 224208 547174
rect 223888 546854 224208 546938
rect 223888 546618 223930 546854
rect 224166 546618 224208 546854
rect 223888 546586 224208 546618
rect 254608 547174 254928 547206
rect 254608 546938 254650 547174
rect 254886 546938 254928 547174
rect 254608 546854 254928 546938
rect 254608 546618 254650 546854
rect 254886 546618 254928 546854
rect 254608 546586 254928 546618
rect 285328 547174 285648 547206
rect 285328 546938 285370 547174
rect 285606 546938 285648 547174
rect 285328 546854 285648 546938
rect 285328 546618 285370 546854
rect 285606 546618 285648 546854
rect 285328 546586 285648 546618
rect 316048 547174 316368 547206
rect 316048 546938 316090 547174
rect 316326 546938 316368 547174
rect 316048 546854 316368 546938
rect 316048 546618 316090 546854
rect 316326 546618 316368 546854
rect 316048 546586 316368 546618
rect 346768 547174 347088 547206
rect 346768 546938 346810 547174
rect 347046 546938 347088 547174
rect 346768 546854 347088 546938
rect 346768 546618 346810 546854
rect 347046 546618 347088 546854
rect 346768 546586 347088 546618
rect 54928 543454 55248 543486
rect 54928 543218 54970 543454
rect 55206 543218 55248 543454
rect 54928 543134 55248 543218
rect 54928 542898 54970 543134
rect 55206 542898 55248 543134
rect 54928 542866 55248 542898
rect 85648 543454 85968 543486
rect 85648 543218 85690 543454
rect 85926 543218 85968 543454
rect 85648 543134 85968 543218
rect 85648 542898 85690 543134
rect 85926 542898 85968 543134
rect 85648 542866 85968 542898
rect 116368 543454 116688 543486
rect 116368 543218 116410 543454
rect 116646 543218 116688 543454
rect 116368 543134 116688 543218
rect 116368 542898 116410 543134
rect 116646 542898 116688 543134
rect 116368 542866 116688 542898
rect 147088 543454 147408 543486
rect 147088 543218 147130 543454
rect 147366 543218 147408 543454
rect 147088 543134 147408 543218
rect 147088 542898 147130 543134
rect 147366 542898 147408 543134
rect 147088 542866 147408 542898
rect 177808 543454 178128 543486
rect 177808 543218 177850 543454
rect 178086 543218 178128 543454
rect 177808 543134 178128 543218
rect 177808 542898 177850 543134
rect 178086 542898 178128 543134
rect 177808 542866 178128 542898
rect 208528 543454 208848 543486
rect 208528 543218 208570 543454
rect 208806 543218 208848 543454
rect 208528 543134 208848 543218
rect 208528 542898 208570 543134
rect 208806 542898 208848 543134
rect 208528 542866 208848 542898
rect 239248 543454 239568 543486
rect 239248 543218 239290 543454
rect 239526 543218 239568 543454
rect 239248 543134 239568 543218
rect 239248 542898 239290 543134
rect 239526 542898 239568 543134
rect 239248 542866 239568 542898
rect 269968 543454 270288 543486
rect 269968 543218 270010 543454
rect 270246 543218 270288 543454
rect 269968 543134 270288 543218
rect 269968 542898 270010 543134
rect 270246 542898 270288 543134
rect 269968 542866 270288 542898
rect 300688 543454 301008 543486
rect 300688 543218 300730 543454
rect 300966 543218 301008 543454
rect 300688 543134 301008 543218
rect 300688 542898 300730 543134
rect 300966 542898 301008 543134
rect 300688 542866 301008 542898
rect 331408 543454 331728 543486
rect 331408 543218 331450 543454
rect 331686 543218 331728 543454
rect 331408 543134 331728 543218
rect 331408 542898 331450 543134
rect 331686 542898 331728 543134
rect 331408 542866 331728 542898
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 24208 507454 24528 507486
rect 24208 507218 24250 507454
rect 24486 507218 24528 507454
rect 24208 507134 24528 507218
rect 24208 506898 24250 507134
rect 24486 506898 24528 507134
rect 24208 506866 24528 506898
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 27834 497494 28454 532938
rect 39568 511174 39888 511206
rect 39568 510938 39610 511174
rect 39846 510938 39888 511174
rect 39568 510854 39888 510938
rect 39568 510618 39610 510854
rect 39846 510618 39888 510854
rect 39568 510586 39888 510618
rect 70288 511174 70608 511206
rect 70288 510938 70330 511174
rect 70566 510938 70608 511174
rect 70288 510854 70608 510938
rect 70288 510618 70330 510854
rect 70566 510618 70608 510854
rect 70288 510586 70608 510618
rect 101008 511174 101328 511206
rect 101008 510938 101050 511174
rect 101286 510938 101328 511174
rect 101008 510854 101328 510938
rect 101008 510618 101050 510854
rect 101286 510618 101328 510854
rect 101008 510586 101328 510618
rect 131728 511174 132048 511206
rect 131728 510938 131770 511174
rect 132006 510938 132048 511174
rect 131728 510854 132048 510938
rect 131728 510618 131770 510854
rect 132006 510618 132048 510854
rect 131728 510586 132048 510618
rect 162448 511174 162768 511206
rect 162448 510938 162490 511174
rect 162726 510938 162768 511174
rect 162448 510854 162768 510938
rect 162448 510618 162490 510854
rect 162726 510618 162768 510854
rect 162448 510586 162768 510618
rect 193168 511174 193488 511206
rect 193168 510938 193210 511174
rect 193446 510938 193488 511174
rect 193168 510854 193488 510938
rect 193168 510618 193210 510854
rect 193446 510618 193488 510854
rect 193168 510586 193488 510618
rect 223888 511174 224208 511206
rect 223888 510938 223930 511174
rect 224166 510938 224208 511174
rect 223888 510854 224208 510938
rect 223888 510618 223930 510854
rect 224166 510618 224208 510854
rect 223888 510586 224208 510618
rect 254608 511174 254928 511206
rect 254608 510938 254650 511174
rect 254886 510938 254928 511174
rect 254608 510854 254928 510938
rect 254608 510618 254650 510854
rect 254886 510618 254928 510854
rect 254608 510586 254928 510618
rect 285328 511174 285648 511206
rect 285328 510938 285370 511174
rect 285606 510938 285648 511174
rect 285328 510854 285648 510938
rect 285328 510618 285370 510854
rect 285606 510618 285648 510854
rect 285328 510586 285648 510618
rect 316048 511174 316368 511206
rect 316048 510938 316090 511174
rect 316326 510938 316368 511174
rect 316048 510854 316368 510938
rect 316048 510618 316090 510854
rect 316326 510618 316368 510854
rect 316048 510586 316368 510618
rect 346768 511174 347088 511206
rect 346768 510938 346810 511174
rect 347046 510938 347088 511174
rect 346768 510854 347088 510938
rect 346768 510618 346810 510854
rect 347046 510618 347088 510854
rect 346768 510586 347088 510618
rect 54928 507454 55248 507486
rect 54928 507218 54970 507454
rect 55206 507218 55248 507454
rect 54928 507134 55248 507218
rect 54928 506898 54970 507134
rect 55206 506898 55248 507134
rect 54928 506866 55248 506898
rect 85648 507454 85968 507486
rect 85648 507218 85690 507454
rect 85926 507218 85968 507454
rect 85648 507134 85968 507218
rect 85648 506898 85690 507134
rect 85926 506898 85968 507134
rect 85648 506866 85968 506898
rect 116368 507454 116688 507486
rect 116368 507218 116410 507454
rect 116646 507218 116688 507454
rect 116368 507134 116688 507218
rect 116368 506898 116410 507134
rect 116646 506898 116688 507134
rect 116368 506866 116688 506898
rect 147088 507454 147408 507486
rect 147088 507218 147130 507454
rect 147366 507218 147408 507454
rect 147088 507134 147408 507218
rect 147088 506898 147130 507134
rect 147366 506898 147408 507134
rect 147088 506866 147408 506898
rect 177808 507454 178128 507486
rect 177808 507218 177850 507454
rect 178086 507218 178128 507454
rect 177808 507134 178128 507218
rect 177808 506898 177850 507134
rect 178086 506898 178128 507134
rect 177808 506866 178128 506898
rect 208528 507454 208848 507486
rect 208528 507218 208570 507454
rect 208806 507218 208848 507454
rect 208528 507134 208848 507218
rect 208528 506898 208570 507134
rect 208806 506898 208848 507134
rect 208528 506866 208848 506898
rect 239248 507454 239568 507486
rect 239248 507218 239290 507454
rect 239526 507218 239568 507454
rect 239248 507134 239568 507218
rect 239248 506898 239290 507134
rect 239526 506898 239568 507134
rect 239248 506866 239568 506898
rect 269968 507454 270288 507486
rect 269968 507218 270010 507454
rect 270246 507218 270288 507454
rect 269968 507134 270288 507218
rect 269968 506898 270010 507134
rect 270246 506898 270288 507134
rect 269968 506866 270288 506898
rect 300688 507454 301008 507486
rect 300688 507218 300730 507454
rect 300966 507218 301008 507454
rect 300688 507134 301008 507218
rect 300688 506898 300730 507134
rect 300966 506898 301008 507134
rect 300688 506866 301008 506898
rect 331408 507454 331728 507486
rect 331408 507218 331450 507454
rect 331686 507218 331728 507454
rect 331408 507134 331728 507218
rect 331408 506898 331450 507134
rect 331686 506898 331728 507134
rect 331408 506866 331728 506898
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 24208 471454 24528 471486
rect 24208 471218 24250 471454
rect 24486 471218 24528 471454
rect 24208 471134 24528 471218
rect 24208 470898 24250 471134
rect 24486 470898 24528 471134
rect 24208 470866 24528 470898
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 27834 461494 28454 496938
rect 39568 475174 39888 475206
rect 39568 474938 39610 475174
rect 39846 474938 39888 475174
rect 39568 474854 39888 474938
rect 39568 474618 39610 474854
rect 39846 474618 39888 474854
rect 39568 474586 39888 474618
rect 70288 475174 70608 475206
rect 70288 474938 70330 475174
rect 70566 474938 70608 475174
rect 70288 474854 70608 474938
rect 70288 474618 70330 474854
rect 70566 474618 70608 474854
rect 70288 474586 70608 474618
rect 101008 475174 101328 475206
rect 101008 474938 101050 475174
rect 101286 474938 101328 475174
rect 101008 474854 101328 474938
rect 101008 474618 101050 474854
rect 101286 474618 101328 474854
rect 101008 474586 101328 474618
rect 131728 475174 132048 475206
rect 131728 474938 131770 475174
rect 132006 474938 132048 475174
rect 131728 474854 132048 474938
rect 131728 474618 131770 474854
rect 132006 474618 132048 474854
rect 131728 474586 132048 474618
rect 162448 475174 162768 475206
rect 162448 474938 162490 475174
rect 162726 474938 162768 475174
rect 162448 474854 162768 474938
rect 162448 474618 162490 474854
rect 162726 474618 162768 474854
rect 162448 474586 162768 474618
rect 193168 475174 193488 475206
rect 193168 474938 193210 475174
rect 193446 474938 193488 475174
rect 193168 474854 193488 474938
rect 193168 474618 193210 474854
rect 193446 474618 193488 474854
rect 193168 474586 193488 474618
rect 223888 475174 224208 475206
rect 223888 474938 223930 475174
rect 224166 474938 224208 475174
rect 223888 474854 224208 474938
rect 223888 474618 223930 474854
rect 224166 474618 224208 474854
rect 223888 474586 224208 474618
rect 254608 475174 254928 475206
rect 254608 474938 254650 475174
rect 254886 474938 254928 475174
rect 254608 474854 254928 474938
rect 254608 474618 254650 474854
rect 254886 474618 254928 474854
rect 254608 474586 254928 474618
rect 285328 475174 285648 475206
rect 285328 474938 285370 475174
rect 285606 474938 285648 475174
rect 285328 474854 285648 474938
rect 285328 474618 285370 474854
rect 285606 474618 285648 474854
rect 285328 474586 285648 474618
rect 316048 475174 316368 475206
rect 316048 474938 316090 475174
rect 316326 474938 316368 475174
rect 316048 474854 316368 474938
rect 316048 474618 316090 474854
rect 316326 474618 316368 474854
rect 316048 474586 316368 474618
rect 346768 475174 347088 475206
rect 346768 474938 346810 475174
rect 347046 474938 347088 475174
rect 346768 474854 347088 474938
rect 346768 474618 346810 474854
rect 347046 474618 347088 474854
rect 346768 474586 347088 474618
rect 54928 471454 55248 471486
rect 54928 471218 54970 471454
rect 55206 471218 55248 471454
rect 54928 471134 55248 471218
rect 54928 470898 54970 471134
rect 55206 470898 55248 471134
rect 54928 470866 55248 470898
rect 85648 471454 85968 471486
rect 85648 471218 85690 471454
rect 85926 471218 85968 471454
rect 85648 471134 85968 471218
rect 85648 470898 85690 471134
rect 85926 470898 85968 471134
rect 85648 470866 85968 470898
rect 116368 471454 116688 471486
rect 116368 471218 116410 471454
rect 116646 471218 116688 471454
rect 116368 471134 116688 471218
rect 116368 470898 116410 471134
rect 116646 470898 116688 471134
rect 116368 470866 116688 470898
rect 147088 471454 147408 471486
rect 147088 471218 147130 471454
rect 147366 471218 147408 471454
rect 147088 471134 147408 471218
rect 147088 470898 147130 471134
rect 147366 470898 147408 471134
rect 147088 470866 147408 470898
rect 177808 471454 178128 471486
rect 177808 471218 177850 471454
rect 178086 471218 178128 471454
rect 177808 471134 178128 471218
rect 177808 470898 177850 471134
rect 178086 470898 178128 471134
rect 177808 470866 178128 470898
rect 208528 471454 208848 471486
rect 208528 471218 208570 471454
rect 208806 471218 208848 471454
rect 208528 471134 208848 471218
rect 208528 470898 208570 471134
rect 208806 470898 208848 471134
rect 208528 470866 208848 470898
rect 239248 471454 239568 471486
rect 239248 471218 239290 471454
rect 239526 471218 239568 471454
rect 239248 471134 239568 471218
rect 239248 470898 239290 471134
rect 239526 470898 239568 471134
rect 239248 470866 239568 470898
rect 269968 471454 270288 471486
rect 269968 471218 270010 471454
rect 270246 471218 270288 471454
rect 269968 471134 270288 471218
rect 269968 470898 270010 471134
rect 270246 470898 270288 471134
rect 269968 470866 270288 470898
rect 300688 471454 301008 471486
rect 300688 471218 300730 471454
rect 300966 471218 301008 471454
rect 300688 471134 301008 471218
rect 300688 470898 300730 471134
rect 300966 470898 301008 471134
rect 300688 470866 301008 470898
rect 331408 471454 331728 471486
rect 331408 471218 331450 471454
rect 331686 471218 331728 471454
rect 331408 471134 331728 471218
rect 331408 470898 331450 471134
rect 331686 470898 331728 471134
rect 331408 470866 331728 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 24208 435454 24528 435486
rect 24208 435218 24250 435454
rect 24486 435218 24528 435454
rect 24208 435134 24528 435218
rect 24208 434898 24250 435134
rect 24486 434898 24528 435134
rect 24208 434866 24528 434898
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 27834 425494 28454 460938
rect 39568 439174 39888 439206
rect 39568 438938 39610 439174
rect 39846 438938 39888 439174
rect 39568 438854 39888 438938
rect 39568 438618 39610 438854
rect 39846 438618 39888 438854
rect 39568 438586 39888 438618
rect 70288 439174 70608 439206
rect 70288 438938 70330 439174
rect 70566 438938 70608 439174
rect 70288 438854 70608 438938
rect 70288 438618 70330 438854
rect 70566 438618 70608 438854
rect 70288 438586 70608 438618
rect 101008 439174 101328 439206
rect 101008 438938 101050 439174
rect 101286 438938 101328 439174
rect 101008 438854 101328 438938
rect 101008 438618 101050 438854
rect 101286 438618 101328 438854
rect 101008 438586 101328 438618
rect 131728 439174 132048 439206
rect 131728 438938 131770 439174
rect 132006 438938 132048 439174
rect 131728 438854 132048 438938
rect 131728 438618 131770 438854
rect 132006 438618 132048 438854
rect 131728 438586 132048 438618
rect 162448 439174 162768 439206
rect 162448 438938 162490 439174
rect 162726 438938 162768 439174
rect 162448 438854 162768 438938
rect 162448 438618 162490 438854
rect 162726 438618 162768 438854
rect 162448 438586 162768 438618
rect 193168 439174 193488 439206
rect 193168 438938 193210 439174
rect 193446 438938 193488 439174
rect 193168 438854 193488 438938
rect 193168 438618 193210 438854
rect 193446 438618 193488 438854
rect 193168 438586 193488 438618
rect 223888 439174 224208 439206
rect 223888 438938 223930 439174
rect 224166 438938 224208 439174
rect 223888 438854 224208 438938
rect 223888 438618 223930 438854
rect 224166 438618 224208 438854
rect 223888 438586 224208 438618
rect 254608 439174 254928 439206
rect 254608 438938 254650 439174
rect 254886 438938 254928 439174
rect 254608 438854 254928 438938
rect 254608 438618 254650 438854
rect 254886 438618 254928 438854
rect 254608 438586 254928 438618
rect 285328 439174 285648 439206
rect 285328 438938 285370 439174
rect 285606 438938 285648 439174
rect 285328 438854 285648 438938
rect 285328 438618 285370 438854
rect 285606 438618 285648 438854
rect 285328 438586 285648 438618
rect 316048 439174 316368 439206
rect 316048 438938 316090 439174
rect 316326 438938 316368 439174
rect 316048 438854 316368 438938
rect 316048 438618 316090 438854
rect 316326 438618 316368 438854
rect 316048 438586 316368 438618
rect 346768 439174 347088 439206
rect 346768 438938 346810 439174
rect 347046 438938 347088 439174
rect 346768 438854 347088 438938
rect 346768 438618 346810 438854
rect 347046 438618 347088 438854
rect 346768 438586 347088 438618
rect 54928 435454 55248 435486
rect 54928 435218 54970 435454
rect 55206 435218 55248 435454
rect 54928 435134 55248 435218
rect 54928 434898 54970 435134
rect 55206 434898 55248 435134
rect 54928 434866 55248 434898
rect 85648 435454 85968 435486
rect 85648 435218 85690 435454
rect 85926 435218 85968 435454
rect 85648 435134 85968 435218
rect 85648 434898 85690 435134
rect 85926 434898 85968 435134
rect 85648 434866 85968 434898
rect 116368 435454 116688 435486
rect 116368 435218 116410 435454
rect 116646 435218 116688 435454
rect 116368 435134 116688 435218
rect 116368 434898 116410 435134
rect 116646 434898 116688 435134
rect 116368 434866 116688 434898
rect 147088 435454 147408 435486
rect 147088 435218 147130 435454
rect 147366 435218 147408 435454
rect 147088 435134 147408 435218
rect 147088 434898 147130 435134
rect 147366 434898 147408 435134
rect 147088 434866 147408 434898
rect 177808 435454 178128 435486
rect 177808 435218 177850 435454
rect 178086 435218 178128 435454
rect 177808 435134 178128 435218
rect 177808 434898 177850 435134
rect 178086 434898 178128 435134
rect 177808 434866 178128 434898
rect 208528 435454 208848 435486
rect 208528 435218 208570 435454
rect 208806 435218 208848 435454
rect 208528 435134 208848 435218
rect 208528 434898 208570 435134
rect 208806 434898 208848 435134
rect 208528 434866 208848 434898
rect 239248 435454 239568 435486
rect 239248 435218 239290 435454
rect 239526 435218 239568 435454
rect 239248 435134 239568 435218
rect 239248 434898 239290 435134
rect 239526 434898 239568 435134
rect 239248 434866 239568 434898
rect 269968 435454 270288 435486
rect 269968 435218 270010 435454
rect 270246 435218 270288 435454
rect 269968 435134 270288 435218
rect 269968 434898 270010 435134
rect 270246 434898 270288 435134
rect 269968 434866 270288 434898
rect 300688 435454 301008 435486
rect 300688 435218 300730 435454
rect 300966 435218 301008 435454
rect 300688 435134 301008 435218
rect 300688 434898 300730 435134
rect 300966 434898 301008 435134
rect 300688 434866 301008 434898
rect 331408 435454 331728 435486
rect 331408 435218 331450 435454
rect 331686 435218 331728 435454
rect 331408 435134 331728 435218
rect 331408 434898 331450 435134
rect 331686 434898 331728 435134
rect 331408 434866 331728 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 24208 399454 24528 399486
rect 24208 399218 24250 399454
rect 24486 399218 24528 399454
rect 24208 399134 24528 399218
rect 24208 398898 24250 399134
rect 24486 398898 24528 399134
rect 24208 398866 24528 398898
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 27834 389494 28454 424938
rect 39568 403174 39888 403206
rect 39568 402938 39610 403174
rect 39846 402938 39888 403174
rect 39568 402854 39888 402938
rect 39568 402618 39610 402854
rect 39846 402618 39888 402854
rect 39568 402586 39888 402618
rect 70288 403174 70608 403206
rect 70288 402938 70330 403174
rect 70566 402938 70608 403174
rect 70288 402854 70608 402938
rect 70288 402618 70330 402854
rect 70566 402618 70608 402854
rect 70288 402586 70608 402618
rect 101008 403174 101328 403206
rect 101008 402938 101050 403174
rect 101286 402938 101328 403174
rect 101008 402854 101328 402938
rect 101008 402618 101050 402854
rect 101286 402618 101328 402854
rect 101008 402586 101328 402618
rect 131728 403174 132048 403206
rect 131728 402938 131770 403174
rect 132006 402938 132048 403174
rect 131728 402854 132048 402938
rect 131728 402618 131770 402854
rect 132006 402618 132048 402854
rect 131728 402586 132048 402618
rect 162448 403174 162768 403206
rect 162448 402938 162490 403174
rect 162726 402938 162768 403174
rect 162448 402854 162768 402938
rect 162448 402618 162490 402854
rect 162726 402618 162768 402854
rect 162448 402586 162768 402618
rect 193168 403174 193488 403206
rect 193168 402938 193210 403174
rect 193446 402938 193488 403174
rect 193168 402854 193488 402938
rect 193168 402618 193210 402854
rect 193446 402618 193488 402854
rect 193168 402586 193488 402618
rect 223888 403174 224208 403206
rect 223888 402938 223930 403174
rect 224166 402938 224208 403174
rect 223888 402854 224208 402938
rect 223888 402618 223930 402854
rect 224166 402618 224208 402854
rect 223888 402586 224208 402618
rect 254608 403174 254928 403206
rect 254608 402938 254650 403174
rect 254886 402938 254928 403174
rect 254608 402854 254928 402938
rect 254608 402618 254650 402854
rect 254886 402618 254928 402854
rect 254608 402586 254928 402618
rect 285328 403174 285648 403206
rect 285328 402938 285370 403174
rect 285606 402938 285648 403174
rect 285328 402854 285648 402938
rect 285328 402618 285370 402854
rect 285606 402618 285648 402854
rect 285328 402586 285648 402618
rect 316048 403174 316368 403206
rect 316048 402938 316090 403174
rect 316326 402938 316368 403174
rect 316048 402854 316368 402938
rect 316048 402618 316090 402854
rect 316326 402618 316368 402854
rect 316048 402586 316368 402618
rect 346768 403174 347088 403206
rect 346768 402938 346810 403174
rect 347046 402938 347088 403174
rect 346768 402854 347088 402938
rect 346768 402618 346810 402854
rect 347046 402618 347088 402854
rect 346768 402586 347088 402618
rect 54928 399454 55248 399486
rect 54928 399218 54970 399454
rect 55206 399218 55248 399454
rect 54928 399134 55248 399218
rect 54928 398898 54970 399134
rect 55206 398898 55248 399134
rect 54928 398866 55248 398898
rect 85648 399454 85968 399486
rect 85648 399218 85690 399454
rect 85926 399218 85968 399454
rect 85648 399134 85968 399218
rect 85648 398898 85690 399134
rect 85926 398898 85968 399134
rect 85648 398866 85968 398898
rect 116368 399454 116688 399486
rect 116368 399218 116410 399454
rect 116646 399218 116688 399454
rect 116368 399134 116688 399218
rect 116368 398898 116410 399134
rect 116646 398898 116688 399134
rect 116368 398866 116688 398898
rect 147088 399454 147408 399486
rect 147088 399218 147130 399454
rect 147366 399218 147408 399454
rect 147088 399134 147408 399218
rect 147088 398898 147130 399134
rect 147366 398898 147408 399134
rect 147088 398866 147408 398898
rect 177808 399454 178128 399486
rect 177808 399218 177850 399454
rect 178086 399218 178128 399454
rect 177808 399134 178128 399218
rect 177808 398898 177850 399134
rect 178086 398898 178128 399134
rect 177808 398866 178128 398898
rect 208528 399454 208848 399486
rect 208528 399218 208570 399454
rect 208806 399218 208848 399454
rect 208528 399134 208848 399218
rect 208528 398898 208570 399134
rect 208806 398898 208848 399134
rect 208528 398866 208848 398898
rect 239248 399454 239568 399486
rect 239248 399218 239290 399454
rect 239526 399218 239568 399454
rect 239248 399134 239568 399218
rect 239248 398898 239290 399134
rect 239526 398898 239568 399134
rect 239248 398866 239568 398898
rect 269968 399454 270288 399486
rect 269968 399218 270010 399454
rect 270246 399218 270288 399454
rect 269968 399134 270288 399218
rect 269968 398898 270010 399134
rect 270246 398898 270288 399134
rect 269968 398866 270288 398898
rect 300688 399454 301008 399486
rect 300688 399218 300730 399454
rect 300966 399218 301008 399454
rect 300688 399134 301008 399218
rect 300688 398898 300730 399134
rect 300966 398898 301008 399134
rect 300688 398866 301008 398898
rect 331408 399454 331728 399486
rect 331408 399218 331450 399454
rect 331686 399218 331728 399454
rect 331408 399134 331728 399218
rect 331408 398898 331450 399134
rect 331686 398898 331728 399134
rect 331408 398866 331728 398898
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 24208 363454 24528 363486
rect 24208 363218 24250 363454
rect 24486 363218 24528 363454
rect 24208 363134 24528 363218
rect 24208 362898 24250 363134
rect 24486 362898 24528 363134
rect 24208 362866 24528 362898
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 27834 353494 28454 388938
rect 39568 367174 39888 367206
rect 39568 366938 39610 367174
rect 39846 366938 39888 367174
rect 39568 366854 39888 366938
rect 39568 366618 39610 366854
rect 39846 366618 39888 366854
rect 39568 366586 39888 366618
rect 70288 367174 70608 367206
rect 70288 366938 70330 367174
rect 70566 366938 70608 367174
rect 70288 366854 70608 366938
rect 70288 366618 70330 366854
rect 70566 366618 70608 366854
rect 70288 366586 70608 366618
rect 101008 367174 101328 367206
rect 101008 366938 101050 367174
rect 101286 366938 101328 367174
rect 101008 366854 101328 366938
rect 101008 366618 101050 366854
rect 101286 366618 101328 366854
rect 101008 366586 101328 366618
rect 131728 367174 132048 367206
rect 131728 366938 131770 367174
rect 132006 366938 132048 367174
rect 131728 366854 132048 366938
rect 131728 366618 131770 366854
rect 132006 366618 132048 366854
rect 131728 366586 132048 366618
rect 162448 367174 162768 367206
rect 162448 366938 162490 367174
rect 162726 366938 162768 367174
rect 162448 366854 162768 366938
rect 162448 366618 162490 366854
rect 162726 366618 162768 366854
rect 162448 366586 162768 366618
rect 193168 367174 193488 367206
rect 193168 366938 193210 367174
rect 193446 366938 193488 367174
rect 193168 366854 193488 366938
rect 193168 366618 193210 366854
rect 193446 366618 193488 366854
rect 193168 366586 193488 366618
rect 223888 367174 224208 367206
rect 223888 366938 223930 367174
rect 224166 366938 224208 367174
rect 223888 366854 224208 366938
rect 223888 366618 223930 366854
rect 224166 366618 224208 366854
rect 223888 366586 224208 366618
rect 254608 367174 254928 367206
rect 254608 366938 254650 367174
rect 254886 366938 254928 367174
rect 254608 366854 254928 366938
rect 254608 366618 254650 366854
rect 254886 366618 254928 366854
rect 254608 366586 254928 366618
rect 285328 367174 285648 367206
rect 285328 366938 285370 367174
rect 285606 366938 285648 367174
rect 285328 366854 285648 366938
rect 285328 366618 285370 366854
rect 285606 366618 285648 366854
rect 285328 366586 285648 366618
rect 316048 367174 316368 367206
rect 316048 366938 316090 367174
rect 316326 366938 316368 367174
rect 316048 366854 316368 366938
rect 316048 366618 316090 366854
rect 316326 366618 316368 366854
rect 316048 366586 316368 366618
rect 346768 367174 347088 367206
rect 346768 366938 346810 367174
rect 347046 366938 347088 367174
rect 346768 366854 347088 366938
rect 346768 366618 346810 366854
rect 347046 366618 347088 366854
rect 346768 366586 347088 366618
rect 54928 363454 55248 363486
rect 54928 363218 54970 363454
rect 55206 363218 55248 363454
rect 54928 363134 55248 363218
rect 54928 362898 54970 363134
rect 55206 362898 55248 363134
rect 54928 362866 55248 362898
rect 85648 363454 85968 363486
rect 85648 363218 85690 363454
rect 85926 363218 85968 363454
rect 85648 363134 85968 363218
rect 85648 362898 85690 363134
rect 85926 362898 85968 363134
rect 85648 362866 85968 362898
rect 116368 363454 116688 363486
rect 116368 363218 116410 363454
rect 116646 363218 116688 363454
rect 116368 363134 116688 363218
rect 116368 362898 116410 363134
rect 116646 362898 116688 363134
rect 116368 362866 116688 362898
rect 147088 363454 147408 363486
rect 147088 363218 147130 363454
rect 147366 363218 147408 363454
rect 147088 363134 147408 363218
rect 147088 362898 147130 363134
rect 147366 362898 147408 363134
rect 147088 362866 147408 362898
rect 177808 363454 178128 363486
rect 177808 363218 177850 363454
rect 178086 363218 178128 363454
rect 177808 363134 178128 363218
rect 177808 362898 177850 363134
rect 178086 362898 178128 363134
rect 177808 362866 178128 362898
rect 208528 363454 208848 363486
rect 208528 363218 208570 363454
rect 208806 363218 208848 363454
rect 208528 363134 208848 363218
rect 208528 362898 208570 363134
rect 208806 362898 208848 363134
rect 208528 362866 208848 362898
rect 239248 363454 239568 363486
rect 239248 363218 239290 363454
rect 239526 363218 239568 363454
rect 239248 363134 239568 363218
rect 239248 362898 239290 363134
rect 239526 362898 239568 363134
rect 239248 362866 239568 362898
rect 269968 363454 270288 363486
rect 269968 363218 270010 363454
rect 270246 363218 270288 363454
rect 269968 363134 270288 363218
rect 269968 362898 270010 363134
rect 270246 362898 270288 363134
rect 269968 362866 270288 362898
rect 300688 363454 301008 363486
rect 300688 363218 300730 363454
rect 300966 363218 301008 363454
rect 300688 363134 301008 363218
rect 300688 362898 300730 363134
rect 300966 362898 301008 363134
rect 300688 362866 301008 362898
rect 331408 363454 331728 363486
rect 331408 363218 331450 363454
rect 331686 363218 331728 363454
rect 331408 363134 331728 363218
rect 331408 362898 331450 363134
rect 331686 362898 331728 363134
rect 331408 362866 331728 362898
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 24208 327454 24528 327486
rect 24208 327218 24250 327454
rect 24486 327218 24528 327454
rect 24208 327134 24528 327218
rect 24208 326898 24250 327134
rect 24486 326898 24528 327134
rect 24208 326866 24528 326898
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 27834 317494 28454 352938
rect 39568 331174 39888 331206
rect 39568 330938 39610 331174
rect 39846 330938 39888 331174
rect 39568 330854 39888 330938
rect 39568 330618 39610 330854
rect 39846 330618 39888 330854
rect 39568 330586 39888 330618
rect 70288 331174 70608 331206
rect 70288 330938 70330 331174
rect 70566 330938 70608 331174
rect 70288 330854 70608 330938
rect 70288 330618 70330 330854
rect 70566 330618 70608 330854
rect 70288 330586 70608 330618
rect 101008 331174 101328 331206
rect 101008 330938 101050 331174
rect 101286 330938 101328 331174
rect 101008 330854 101328 330938
rect 101008 330618 101050 330854
rect 101286 330618 101328 330854
rect 101008 330586 101328 330618
rect 131728 331174 132048 331206
rect 131728 330938 131770 331174
rect 132006 330938 132048 331174
rect 131728 330854 132048 330938
rect 131728 330618 131770 330854
rect 132006 330618 132048 330854
rect 131728 330586 132048 330618
rect 162448 331174 162768 331206
rect 162448 330938 162490 331174
rect 162726 330938 162768 331174
rect 162448 330854 162768 330938
rect 162448 330618 162490 330854
rect 162726 330618 162768 330854
rect 162448 330586 162768 330618
rect 193168 331174 193488 331206
rect 193168 330938 193210 331174
rect 193446 330938 193488 331174
rect 193168 330854 193488 330938
rect 193168 330618 193210 330854
rect 193446 330618 193488 330854
rect 193168 330586 193488 330618
rect 223888 331174 224208 331206
rect 223888 330938 223930 331174
rect 224166 330938 224208 331174
rect 223888 330854 224208 330938
rect 223888 330618 223930 330854
rect 224166 330618 224208 330854
rect 223888 330586 224208 330618
rect 254608 331174 254928 331206
rect 254608 330938 254650 331174
rect 254886 330938 254928 331174
rect 254608 330854 254928 330938
rect 254608 330618 254650 330854
rect 254886 330618 254928 330854
rect 254608 330586 254928 330618
rect 285328 331174 285648 331206
rect 285328 330938 285370 331174
rect 285606 330938 285648 331174
rect 285328 330854 285648 330938
rect 285328 330618 285370 330854
rect 285606 330618 285648 330854
rect 285328 330586 285648 330618
rect 316048 331174 316368 331206
rect 316048 330938 316090 331174
rect 316326 330938 316368 331174
rect 316048 330854 316368 330938
rect 316048 330618 316090 330854
rect 316326 330618 316368 330854
rect 316048 330586 316368 330618
rect 346768 331174 347088 331206
rect 346768 330938 346810 331174
rect 347046 330938 347088 331174
rect 346768 330854 347088 330938
rect 346768 330618 346810 330854
rect 347046 330618 347088 330854
rect 346768 330586 347088 330618
rect 54928 327454 55248 327486
rect 54928 327218 54970 327454
rect 55206 327218 55248 327454
rect 54928 327134 55248 327218
rect 54928 326898 54970 327134
rect 55206 326898 55248 327134
rect 54928 326866 55248 326898
rect 85648 327454 85968 327486
rect 85648 327218 85690 327454
rect 85926 327218 85968 327454
rect 85648 327134 85968 327218
rect 85648 326898 85690 327134
rect 85926 326898 85968 327134
rect 85648 326866 85968 326898
rect 116368 327454 116688 327486
rect 116368 327218 116410 327454
rect 116646 327218 116688 327454
rect 116368 327134 116688 327218
rect 116368 326898 116410 327134
rect 116646 326898 116688 327134
rect 116368 326866 116688 326898
rect 147088 327454 147408 327486
rect 147088 327218 147130 327454
rect 147366 327218 147408 327454
rect 147088 327134 147408 327218
rect 147088 326898 147130 327134
rect 147366 326898 147408 327134
rect 147088 326866 147408 326898
rect 177808 327454 178128 327486
rect 177808 327218 177850 327454
rect 178086 327218 178128 327454
rect 177808 327134 178128 327218
rect 177808 326898 177850 327134
rect 178086 326898 178128 327134
rect 177808 326866 178128 326898
rect 208528 327454 208848 327486
rect 208528 327218 208570 327454
rect 208806 327218 208848 327454
rect 208528 327134 208848 327218
rect 208528 326898 208570 327134
rect 208806 326898 208848 327134
rect 208528 326866 208848 326898
rect 239248 327454 239568 327486
rect 239248 327218 239290 327454
rect 239526 327218 239568 327454
rect 239248 327134 239568 327218
rect 239248 326898 239290 327134
rect 239526 326898 239568 327134
rect 239248 326866 239568 326898
rect 269968 327454 270288 327486
rect 269968 327218 270010 327454
rect 270246 327218 270288 327454
rect 269968 327134 270288 327218
rect 269968 326898 270010 327134
rect 270246 326898 270288 327134
rect 269968 326866 270288 326898
rect 300688 327454 301008 327486
rect 300688 327218 300730 327454
rect 300966 327218 301008 327454
rect 300688 327134 301008 327218
rect 300688 326898 300730 327134
rect 300966 326898 301008 327134
rect 300688 326866 301008 326898
rect 331408 327454 331728 327486
rect 331408 327218 331450 327454
rect 331686 327218 331728 327454
rect 331408 327134 331728 327218
rect 331408 326898 331450 327134
rect 331686 326898 331728 327134
rect 331408 326866 331728 326898
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 24208 291454 24528 291486
rect 24208 291218 24250 291454
rect 24486 291218 24528 291454
rect 24208 291134 24528 291218
rect 24208 290898 24250 291134
rect 24486 290898 24528 291134
rect 24208 290866 24528 290898
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 27834 281494 28454 316938
rect 39568 295174 39888 295206
rect 39568 294938 39610 295174
rect 39846 294938 39888 295174
rect 39568 294854 39888 294938
rect 39568 294618 39610 294854
rect 39846 294618 39888 294854
rect 39568 294586 39888 294618
rect 70288 295174 70608 295206
rect 70288 294938 70330 295174
rect 70566 294938 70608 295174
rect 70288 294854 70608 294938
rect 70288 294618 70330 294854
rect 70566 294618 70608 294854
rect 70288 294586 70608 294618
rect 101008 295174 101328 295206
rect 101008 294938 101050 295174
rect 101286 294938 101328 295174
rect 101008 294854 101328 294938
rect 101008 294618 101050 294854
rect 101286 294618 101328 294854
rect 101008 294586 101328 294618
rect 131728 295174 132048 295206
rect 131728 294938 131770 295174
rect 132006 294938 132048 295174
rect 131728 294854 132048 294938
rect 131728 294618 131770 294854
rect 132006 294618 132048 294854
rect 131728 294586 132048 294618
rect 162448 295174 162768 295206
rect 162448 294938 162490 295174
rect 162726 294938 162768 295174
rect 162448 294854 162768 294938
rect 162448 294618 162490 294854
rect 162726 294618 162768 294854
rect 162448 294586 162768 294618
rect 193168 295174 193488 295206
rect 193168 294938 193210 295174
rect 193446 294938 193488 295174
rect 193168 294854 193488 294938
rect 193168 294618 193210 294854
rect 193446 294618 193488 294854
rect 193168 294586 193488 294618
rect 223888 295174 224208 295206
rect 223888 294938 223930 295174
rect 224166 294938 224208 295174
rect 223888 294854 224208 294938
rect 223888 294618 223930 294854
rect 224166 294618 224208 294854
rect 223888 294586 224208 294618
rect 254608 295174 254928 295206
rect 254608 294938 254650 295174
rect 254886 294938 254928 295174
rect 254608 294854 254928 294938
rect 254608 294618 254650 294854
rect 254886 294618 254928 294854
rect 254608 294586 254928 294618
rect 285328 295174 285648 295206
rect 285328 294938 285370 295174
rect 285606 294938 285648 295174
rect 285328 294854 285648 294938
rect 285328 294618 285370 294854
rect 285606 294618 285648 294854
rect 285328 294586 285648 294618
rect 316048 295174 316368 295206
rect 316048 294938 316090 295174
rect 316326 294938 316368 295174
rect 316048 294854 316368 294938
rect 316048 294618 316090 294854
rect 316326 294618 316368 294854
rect 316048 294586 316368 294618
rect 346768 295174 347088 295206
rect 346768 294938 346810 295174
rect 347046 294938 347088 295174
rect 346768 294854 347088 294938
rect 346768 294618 346810 294854
rect 347046 294618 347088 294854
rect 346768 294586 347088 294618
rect 54928 291454 55248 291486
rect 54928 291218 54970 291454
rect 55206 291218 55248 291454
rect 54928 291134 55248 291218
rect 54928 290898 54970 291134
rect 55206 290898 55248 291134
rect 54928 290866 55248 290898
rect 85648 291454 85968 291486
rect 85648 291218 85690 291454
rect 85926 291218 85968 291454
rect 85648 291134 85968 291218
rect 85648 290898 85690 291134
rect 85926 290898 85968 291134
rect 85648 290866 85968 290898
rect 116368 291454 116688 291486
rect 116368 291218 116410 291454
rect 116646 291218 116688 291454
rect 116368 291134 116688 291218
rect 116368 290898 116410 291134
rect 116646 290898 116688 291134
rect 116368 290866 116688 290898
rect 147088 291454 147408 291486
rect 147088 291218 147130 291454
rect 147366 291218 147408 291454
rect 147088 291134 147408 291218
rect 147088 290898 147130 291134
rect 147366 290898 147408 291134
rect 147088 290866 147408 290898
rect 177808 291454 178128 291486
rect 177808 291218 177850 291454
rect 178086 291218 178128 291454
rect 177808 291134 178128 291218
rect 177808 290898 177850 291134
rect 178086 290898 178128 291134
rect 177808 290866 178128 290898
rect 208528 291454 208848 291486
rect 208528 291218 208570 291454
rect 208806 291218 208848 291454
rect 208528 291134 208848 291218
rect 208528 290898 208570 291134
rect 208806 290898 208848 291134
rect 208528 290866 208848 290898
rect 239248 291454 239568 291486
rect 239248 291218 239290 291454
rect 239526 291218 239568 291454
rect 239248 291134 239568 291218
rect 239248 290898 239290 291134
rect 239526 290898 239568 291134
rect 239248 290866 239568 290898
rect 269968 291454 270288 291486
rect 269968 291218 270010 291454
rect 270246 291218 270288 291454
rect 269968 291134 270288 291218
rect 269968 290898 270010 291134
rect 270246 290898 270288 291134
rect 269968 290866 270288 290898
rect 300688 291454 301008 291486
rect 300688 291218 300730 291454
rect 300966 291218 301008 291454
rect 300688 291134 301008 291218
rect 300688 290898 300730 291134
rect 300966 290898 301008 291134
rect 300688 290866 301008 290898
rect 331408 291454 331728 291486
rect 331408 291218 331450 291454
rect 331686 291218 331728 291454
rect 331408 291134 331728 291218
rect 331408 290898 331450 291134
rect 331686 290898 331728 291134
rect 331408 290866 331728 290898
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 24208 255454 24528 255486
rect 24208 255218 24250 255454
rect 24486 255218 24528 255454
rect 24208 255134 24528 255218
rect 24208 254898 24250 255134
rect 24486 254898 24528 255134
rect 24208 254866 24528 254898
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 27834 245494 28454 280938
rect 39568 259174 39888 259206
rect 39568 258938 39610 259174
rect 39846 258938 39888 259174
rect 39568 258854 39888 258938
rect 39568 258618 39610 258854
rect 39846 258618 39888 258854
rect 39568 258586 39888 258618
rect 70288 259174 70608 259206
rect 70288 258938 70330 259174
rect 70566 258938 70608 259174
rect 70288 258854 70608 258938
rect 70288 258618 70330 258854
rect 70566 258618 70608 258854
rect 70288 258586 70608 258618
rect 101008 259174 101328 259206
rect 101008 258938 101050 259174
rect 101286 258938 101328 259174
rect 101008 258854 101328 258938
rect 101008 258618 101050 258854
rect 101286 258618 101328 258854
rect 101008 258586 101328 258618
rect 131728 259174 132048 259206
rect 131728 258938 131770 259174
rect 132006 258938 132048 259174
rect 131728 258854 132048 258938
rect 131728 258618 131770 258854
rect 132006 258618 132048 258854
rect 131728 258586 132048 258618
rect 162448 259174 162768 259206
rect 162448 258938 162490 259174
rect 162726 258938 162768 259174
rect 162448 258854 162768 258938
rect 162448 258618 162490 258854
rect 162726 258618 162768 258854
rect 162448 258586 162768 258618
rect 193168 259174 193488 259206
rect 193168 258938 193210 259174
rect 193446 258938 193488 259174
rect 193168 258854 193488 258938
rect 193168 258618 193210 258854
rect 193446 258618 193488 258854
rect 193168 258586 193488 258618
rect 223888 259174 224208 259206
rect 223888 258938 223930 259174
rect 224166 258938 224208 259174
rect 223888 258854 224208 258938
rect 223888 258618 223930 258854
rect 224166 258618 224208 258854
rect 223888 258586 224208 258618
rect 254608 259174 254928 259206
rect 254608 258938 254650 259174
rect 254886 258938 254928 259174
rect 254608 258854 254928 258938
rect 254608 258618 254650 258854
rect 254886 258618 254928 258854
rect 254608 258586 254928 258618
rect 285328 259174 285648 259206
rect 285328 258938 285370 259174
rect 285606 258938 285648 259174
rect 285328 258854 285648 258938
rect 285328 258618 285370 258854
rect 285606 258618 285648 258854
rect 285328 258586 285648 258618
rect 316048 259174 316368 259206
rect 316048 258938 316090 259174
rect 316326 258938 316368 259174
rect 316048 258854 316368 258938
rect 316048 258618 316090 258854
rect 316326 258618 316368 258854
rect 316048 258586 316368 258618
rect 346768 259174 347088 259206
rect 346768 258938 346810 259174
rect 347046 258938 347088 259174
rect 346768 258854 347088 258938
rect 346768 258618 346810 258854
rect 347046 258618 347088 258854
rect 346768 258586 347088 258618
rect 54928 255454 55248 255486
rect 54928 255218 54970 255454
rect 55206 255218 55248 255454
rect 54928 255134 55248 255218
rect 54928 254898 54970 255134
rect 55206 254898 55248 255134
rect 54928 254866 55248 254898
rect 85648 255454 85968 255486
rect 85648 255218 85690 255454
rect 85926 255218 85968 255454
rect 85648 255134 85968 255218
rect 85648 254898 85690 255134
rect 85926 254898 85968 255134
rect 85648 254866 85968 254898
rect 116368 255454 116688 255486
rect 116368 255218 116410 255454
rect 116646 255218 116688 255454
rect 116368 255134 116688 255218
rect 116368 254898 116410 255134
rect 116646 254898 116688 255134
rect 116368 254866 116688 254898
rect 147088 255454 147408 255486
rect 147088 255218 147130 255454
rect 147366 255218 147408 255454
rect 147088 255134 147408 255218
rect 147088 254898 147130 255134
rect 147366 254898 147408 255134
rect 147088 254866 147408 254898
rect 177808 255454 178128 255486
rect 177808 255218 177850 255454
rect 178086 255218 178128 255454
rect 177808 255134 178128 255218
rect 177808 254898 177850 255134
rect 178086 254898 178128 255134
rect 177808 254866 178128 254898
rect 208528 255454 208848 255486
rect 208528 255218 208570 255454
rect 208806 255218 208848 255454
rect 208528 255134 208848 255218
rect 208528 254898 208570 255134
rect 208806 254898 208848 255134
rect 208528 254866 208848 254898
rect 239248 255454 239568 255486
rect 239248 255218 239290 255454
rect 239526 255218 239568 255454
rect 239248 255134 239568 255218
rect 239248 254898 239290 255134
rect 239526 254898 239568 255134
rect 239248 254866 239568 254898
rect 269968 255454 270288 255486
rect 269968 255218 270010 255454
rect 270246 255218 270288 255454
rect 269968 255134 270288 255218
rect 269968 254898 270010 255134
rect 270246 254898 270288 255134
rect 269968 254866 270288 254898
rect 300688 255454 301008 255486
rect 300688 255218 300730 255454
rect 300966 255218 301008 255454
rect 300688 255134 301008 255218
rect 300688 254898 300730 255134
rect 300966 254898 301008 255134
rect 300688 254866 301008 254898
rect 331408 255454 331728 255486
rect 331408 255218 331450 255454
rect 331686 255218 331728 255454
rect 331408 255134 331728 255218
rect 331408 254898 331450 255134
rect 331686 254898 331728 255134
rect 331408 254866 331728 254898
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 24208 219454 24528 219486
rect 24208 219218 24250 219454
rect 24486 219218 24528 219454
rect 24208 219134 24528 219218
rect 24208 218898 24250 219134
rect 24486 218898 24528 219134
rect 24208 218866 24528 218898
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 27834 209494 28454 244938
rect 39568 223174 39888 223206
rect 39568 222938 39610 223174
rect 39846 222938 39888 223174
rect 39568 222854 39888 222938
rect 39568 222618 39610 222854
rect 39846 222618 39888 222854
rect 39568 222586 39888 222618
rect 70288 223174 70608 223206
rect 70288 222938 70330 223174
rect 70566 222938 70608 223174
rect 70288 222854 70608 222938
rect 70288 222618 70330 222854
rect 70566 222618 70608 222854
rect 70288 222586 70608 222618
rect 101008 223174 101328 223206
rect 101008 222938 101050 223174
rect 101286 222938 101328 223174
rect 101008 222854 101328 222938
rect 101008 222618 101050 222854
rect 101286 222618 101328 222854
rect 101008 222586 101328 222618
rect 131728 223174 132048 223206
rect 131728 222938 131770 223174
rect 132006 222938 132048 223174
rect 131728 222854 132048 222938
rect 131728 222618 131770 222854
rect 132006 222618 132048 222854
rect 131728 222586 132048 222618
rect 162448 223174 162768 223206
rect 162448 222938 162490 223174
rect 162726 222938 162768 223174
rect 162448 222854 162768 222938
rect 162448 222618 162490 222854
rect 162726 222618 162768 222854
rect 162448 222586 162768 222618
rect 193168 223174 193488 223206
rect 193168 222938 193210 223174
rect 193446 222938 193488 223174
rect 193168 222854 193488 222938
rect 193168 222618 193210 222854
rect 193446 222618 193488 222854
rect 193168 222586 193488 222618
rect 223888 223174 224208 223206
rect 223888 222938 223930 223174
rect 224166 222938 224208 223174
rect 223888 222854 224208 222938
rect 223888 222618 223930 222854
rect 224166 222618 224208 222854
rect 223888 222586 224208 222618
rect 254608 223174 254928 223206
rect 254608 222938 254650 223174
rect 254886 222938 254928 223174
rect 254608 222854 254928 222938
rect 254608 222618 254650 222854
rect 254886 222618 254928 222854
rect 254608 222586 254928 222618
rect 285328 223174 285648 223206
rect 285328 222938 285370 223174
rect 285606 222938 285648 223174
rect 285328 222854 285648 222938
rect 285328 222618 285370 222854
rect 285606 222618 285648 222854
rect 285328 222586 285648 222618
rect 316048 223174 316368 223206
rect 316048 222938 316090 223174
rect 316326 222938 316368 223174
rect 316048 222854 316368 222938
rect 316048 222618 316090 222854
rect 316326 222618 316368 222854
rect 316048 222586 316368 222618
rect 346768 223174 347088 223206
rect 346768 222938 346810 223174
rect 347046 222938 347088 223174
rect 346768 222854 347088 222938
rect 346768 222618 346810 222854
rect 347046 222618 347088 222854
rect 346768 222586 347088 222618
rect 54928 219454 55248 219486
rect 54928 219218 54970 219454
rect 55206 219218 55248 219454
rect 54928 219134 55248 219218
rect 54928 218898 54970 219134
rect 55206 218898 55248 219134
rect 54928 218866 55248 218898
rect 85648 219454 85968 219486
rect 85648 219218 85690 219454
rect 85926 219218 85968 219454
rect 85648 219134 85968 219218
rect 85648 218898 85690 219134
rect 85926 218898 85968 219134
rect 85648 218866 85968 218898
rect 116368 219454 116688 219486
rect 116368 219218 116410 219454
rect 116646 219218 116688 219454
rect 116368 219134 116688 219218
rect 116368 218898 116410 219134
rect 116646 218898 116688 219134
rect 116368 218866 116688 218898
rect 147088 219454 147408 219486
rect 147088 219218 147130 219454
rect 147366 219218 147408 219454
rect 147088 219134 147408 219218
rect 147088 218898 147130 219134
rect 147366 218898 147408 219134
rect 147088 218866 147408 218898
rect 177808 219454 178128 219486
rect 177808 219218 177850 219454
rect 178086 219218 178128 219454
rect 177808 219134 178128 219218
rect 177808 218898 177850 219134
rect 178086 218898 178128 219134
rect 177808 218866 178128 218898
rect 208528 219454 208848 219486
rect 208528 219218 208570 219454
rect 208806 219218 208848 219454
rect 208528 219134 208848 219218
rect 208528 218898 208570 219134
rect 208806 218898 208848 219134
rect 208528 218866 208848 218898
rect 239248 219454 239568 219486
rect 239248 219218 239290 219454
rect 239526 219218 239568 219454
rect 239248 219134 239568 219218
rect 239248 218898 239290 219134
rect 239526 218898 239568 219134
rect 239248 218866 239568 218898
rect 269968 219454 270288 219486
rect 269968 219218 270010 219454
rect 270246 219218 270288 219454
rect 269968 219134 270288 219218
rect 269968 218898 270010 219134
rect 270246 218898 270288 219134
rect 269968 218866 270288 218898
rect 300688 219454 301008 219486
rect 300688 219218 300730 219454
rect 300966 219218 301008 219454
rect 300688 219134 301008 219218
rect 300688 218898 300730 219134
rect 300966 218898 301008 219134
rect 300688 218866 301008 218898
rect 331408 219454 331728 219486
rect 331408 219218 331450 219454
rect 331686 219218 331728 219454
rect 331408 219134 331728 219218
rect 331408 218898 331450 219134
rect 331686 218898 331728 219134
rect 331408 218866 331728 218898
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 24208 183454 24528 183486
rect 24208 183218 24250 183454
rect 24486 183218 24528 183454
rect 24208 183134 24528 183218
rect 24208 182898 24250 183134
rect 24486 182898 24528 183134
rect 24208 182866 24528 182898
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 27834 173494 28454 208938
rect 39568 187174 39888 187206
rect 39568 186938 39610 187174
rect 39846 186938 39888 187174
rect 39568 186854 39888 186938
rect 39568 186618 39610 186854
rect 39846 186618 39888 186854
rect 39568 186586 39888 186618
rect 70288 187174 70608 187206
rect 70288 186938 70330 187174
rect 70566 186938 70608 187174
rect 70288 186854 70608 186938
rect 70288 186618 70330 186854
rect 70566 186618 70608 186854
rect 70288 186586 70608 186618
rect 101008 187174 101328 187206
rect 101008 186938 101050 187174
rect 101286 186938 101328 187174
rect 101008 186854 101328 186938
rect 101008 186618 101050 186854
rect 101286 186618 101328 186854
rect 101008 186586 101328 186618
rect 131728 187174 132048 187206
rect 131728 186938 131770 187174
rect 132006 186938 132048 187174
rect 131728 186854 132048 186938
rect 131728 186618 131770 186854
rect 132006 186618 132048 186854
rect 131728 186586 132048 186618
rect 162448 187174 162768 187206
rect 162448 186938 162490 187174
rect 162726 186938 162768 187174
rect 162448 186854 162768 186938
rect 162448 186618 162490 186854
rect 162726 186618 162768 186854
rect 162448 186586 162768 186618
rect 193168 187174 193488 187206
rect 193168 186938 193210 187174
rect 193446 186938 193488 187174
rect 193168 186854 193488 186938
rect 193168 186618 193210 186854
rect 193446 186618 193488 186854
rect 193168 186586 193488 186618
rect 223888 187174 224208 187206
rect 223888 186938 223930 187174
rect 224166 186938 224208 187174
rect 223888 186854 224208 186938
rect 223888 186618 223930 186854
rect 224166 186618 224208 186854
rect 223888 186586 224208 186618
rect 254608 187174 254928 187206
rect 254608 186938 254650 187174
rect 254886 186938 254928 187174
rect 254608 186854 254928 186938
rect 254608 186618 254650 186854
rect 254886 186618 254928 186854
rect 254608 186586 254928 186618
rect 285328 187174 285648 187206
rect 285328 186938 285370 187174
rect 285606 186938 285648 187174
rect 285328 186854 285648 186938
rect 285328 186618 285370 186854
rect 285606 186618 285648 186854
rect 285328 186586 285648 186618
rect 316048 187174 316368 187206
rect 316048 186938 316090 187174
rect 316326 186938 316368 187174
rect 316048 186854 316368 186938
rect 316048 186618 316090 186854
rect 316326 186618 316368 186854
rect 316048 186586 316368 186618
rect 346768 187174 347088 187206
rect 346768 186938 346810 187174
rect 347046 186938 347088 187174
rect 346768 186854 347088 186938
rect 346768 186618 346810 186854
rect 347046 186618 347088 186854
rect 346768 186586 347088 186618
rect 54928 183454 55248 183486
rect 54928 183218 54970 183454
rect 55206 183218 55248 183454
rect 54928 183134 55248 183218
rect 54928 182898 54970 183134
rect 55206 182898 55248 183134
rect 54928 182866 55248 182898
rect 85648 183454 85968 183486
rect 85648 183218 85690 183454
rect 85926 183218 85968 183454
rect 85648 183134 85968 183218
rect 85648 182898 85690 183134
rect 85926 182898 85968 183134
rect 85648 182866 85968 182898
rect 116368 183454 116688 183486
rect 116368 183218 116410 183454
rect 116646 183218 116688 183454
rect 116368 183134 116688 183218
rect 116368 182898 116410 183134
rect 116646 182898 116688 183134
rect 116368 182866 116688 182898
rect 147088 183454 147408 183486
rect 147088 183218 147130 183454
rect 147366 183218 147408 183454
rect 147088 183134 147408 183218
rect 147088 182898 147130 183134
rect 147366 182898 147408 183134
rect 147088 182866 147408 182898
rect 177808 183454 178128 183486
rect 177808 183218 177850 183454
rect 178086 183218 178128 183454
rect 177808 183134 178128 183218
rect 177808 182898 177850 183134
rect 178086 182898 178128 183134
rect 177808 182866 178128 182898
rect 208528 183454 208848 183486
rect 208528 183218 208570 183454
rect 208806 183218 208848 183454
rect 208528 183134 208848 183218
rect 208528 182898 208570 183134
rect 208806 182898 208848 183134
rect 208528 182866 208848 182898
rect 239248 183454 239568 183486
rect 239248 183218 239290 183454
rect 239526 183218 239568 183454
rect 239248 183134 239568 183218
rect 239248 182898 239290 183134
rect 239526 182898 239568 183134
rect 239248 182866 239568 182898
rect 269968 183454 270288 183486
rect 269968 183218 270010 183454
rect 270246 183218 270288 183454
rect 269968 183134 270288 183218
rect 269968 182898 270010 183134
rect 270246 182898 270288 183134
rect 269968 182866 270288 182898
rect 300688 183454 301008 183486
rect 300688 183218 300730 183454
rect 300966 183218 301008 183454
rect 300688 183134 301008 183218
rect 300688 182898 300730 183134
rect 300966 182898 301008 183134
rect 300688 182866 301008 182898
rect 331408 183454 331728 183486
rect 331408 183218 331450 183454
rect 331686 183218 331728 183454
rect 331408 183134 331728 183218
rect 331408 182898 331450 183134
rect 331686 182898 331728 183134
rect 331408 182866 331728 182898
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 24208 147454 24528 147486
rect 24208 147218 24250 147454
rect 24486 147218 24528 147454
rect 24208 147134 24528 147218
rect 24208 146898 24250 147134
rect 24486 146898 24528 147134
rect 24208 146866 24528 146898
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 27834 137494 28454 172938
rect 39568 151174 39888 151206
rect 39568 150938 39610 151174
rect 39846 150938 39888 151174
rect 39568 150854 39888 150938
rect 39568 150618 39610 150854
rect 39846 150618 39888 150854
rect 39568 150586 39888 150618
rect 70288 151174 70608 151206
rect 70288 150938 70330 151174
rect 70566 150938 70608 151174
rect 70288 150854 70608 150938
rect 70288 150618 70330 150854
rect 70566 150618 70608 150854
rect 70288 150586 70608 150618
rect 101008 151174 101328 151206
rect 101008 150938 101050 151174
rect 101286 150938 101328 151174
rect 101008 150854 101328 150938
rect 101008 150618 101050 150854
rect 101286 150618 101328 150854
rect 101008 150586 101328 150618
rect 131728 151174 132048 151206
rect 131728 150938 131770 151174
rect 132006 150938 132048 151174
rect 131728 150854 132048 150938
rect 131728 150618 131770 150854
rect 132006 150618 132048 150854
rect 131728 150586 132048 150618
rect 162448 151174 162768 151206
rect 162448 150938 162490 151174
rect 162726 150938 162768 151174
rect 162448 150854 162768 150938
rect 162448 150618 162490 150854
rect 162726 150618 162768 150854
rect 162448 150586 162768 150618
rect 193168 151174 193488 151206
rect 193168 150938 193210 151174
rect 193446 150938 193488 151174
rect 193168 150854 193488 150938
rect 193168 150618 193210 150854
rect 193446 150618 193488 150854
rect 193168 150586 193488 150618
rect 223888 151174 224208 151206
rect 223888 150938 223930 151174
rect 224166 150938 224208 151174
rect 223888 150854 224208 150938
rect 223888 150618 223930 150854
rect 224166 150618 224208 150854
rect 223888 150586 224208 150618
rect 254608 151174 254928 151206
rect 254608 150938 254650 151174
rect 254886 150938 254928 151174
rect 254608 150854 254928 150938
rect 254608 150618 254650 150854
rect 254886 150618 254928 150854
rect 254608 150586 254928 150618
rect 285328 151174 285648 151206
rect 285328 150938 285370 151174
rect 285606 150938 285648 151174
rect 285328 150854 285648 150938
rect 285328 150618 285370 150854
rect 285606 150618 285648 150854
rect 285328 150586 285648 150618
rect 316048 151174 316368 151206
rect 316048 150938 316090 151174
rect 316326 150938 316368 151174
rect 316048 150854 316368 150938
rect 316048 150618 316090 150854
rect 316326 150618 316368 150854
rect 316048 150586 316368 150618
rect 346768 151174 347088 151206
rect 346768 150938 346810 151174
rect 347046 150938 347088 151174
rect 346768 150854 347088 150938
rect 346768 150618 346810 150854
rect 347046 150618 347088 150854
rect 346768 150586 347088 150618
rect 54928 147454 55248 147486
rect 54928 147218 54970 147454
rect 55206 147218 55248 147454
rect 54928 147134 55248 147218
rect 54928 146898 54970 147134
rect 55206 146898 55248 147134
rect 54928 146866 55248 146898
rect 85648 147454 85968 147486
rect 85648 147218 85690 147454
rect 85926 147218 85968 147454
rect 85648 147134 85968 147218
rect 85648 146898 85690 147134
rect 85926 146898 85968 147134
rect 85648 146866 85968 146898
rect 116368 147454 116688 147486
rect 116368 147218 116410 147454
rect 116646 147218 116688 147454
rect 116368 147134 116688 147218
rect 116368 146898 116410 147134
rect 116646 146898 116688 147134
rect 116368 146866 116688 146898
rect 147088 147454 147408 147486
rect 147088 147218 147130 147454
rect 147366 147218 147408 147454
rect 147088 147134 147408 147218
rect 147088 146898 147130 147134
rect 147366 146898 147408 147134
rect 147088 146866 147408 146898
rect 177808 147454 178128 147486
rect 177808 147218 177850 147454
rect 178086 147218 178128 147454
rect 177808 147134 178128 147218
rect 177808 146898 177850 147134
rect 178086 146898 178128 147134
rect 177808 146866 178128 146898
rect 208528 147454 208848 147486
rect 208528 147218 208570 147454
rect 208806 147218 208848 147454
rect 208528 147134 208848 147218
rect 208528 146898 208570 147134
rect 208806 146898 208848 147134
rect 208528 146866 208848 146898
rect 239248 147454 239568 147486
rect 239248 147218 239290 147454
rect 239526 147218 239568 147454
rect 239248 147134 239568 147218
rect 239248 146898 239290 147134
rect 239526 146898 239568 147134
rect 239248 146866 239568 146898
rect 269968 147454 270288 147486
rect 269968 147218 270010 147454
rect 270246 147218 270288 147454
rect 269968 147134 270288 147218
rect 269968 146898 270010 147134
rect 270246 146898 270288 147134
rect 269968 146866 270288 146898
rect 300688 147454 301008 147486
rect 300688 147218 300730 147454
rect 300966 147218 301008 147454
rect 300688 147134 301008 147218
rect 300688 146898 300730 147134
rect 300966 146898 301008 147134
rect 300688 146866 301008 146898
rect 331408 147454 331728 147486
rect 331408 147218 331450 147454
rect 331686 147218 331728 147454
rect 331408 147134 331728 147218
rect 331408 146898 331450 147134
rect 331686 146898 331728 147134
rect 331408 146866 331728 146898
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 24208 111454 24528 111486
rect 24208 111218 24250 111454
rect 24486 111218 24528 111454
rect 24208 111134 24528 111218
rect 24208 110898 24250 111134
rect 24486 110898 24528 111134
rect 24208 110866 24528 110898
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 27834 101494 28454 136938
rect 39568 115174 39888 115206
rect 39568 114938 39610 115174
rect 39846 114938 39888 115174
rect 39568 114854 39888 114938
rect 39568 114618 39610 114854
rect 39846 114618 39888 114854
rect 39568 114586 39888 114618
rect 70288 115174 70608 115206
rect 70288 114938 70330 115174
rect 70566 114938 70608 115174
rect 70288 114854 70608 114938
rect 70288 114618 70330 114854
rect 70566 114618 70608 114854
rect 70288 114586 70608 114618
rect 101008 115174 101328 115206
rect 101008 114938 101050 115174
rect 101286 114938 101328 115174
rect 101008 114854 101328 114938
rect 101008 114618 101050 114854
rect 101286 114618 101328 114854
rect 101008 114586 101328 114618
rect 131728 115174 132048 115206
rect 131728 114938 131770 115174
rect 132006 114938 132048 115174
rect 131728 114854 132048 114938
rect 131728 114618 131770 114854
rect 132006 114618 132048 114854
rect 131728 114586 132048 114618
rect 162448 115174 162768 115206
rect 162448 114938 162490 115174
rect 162726 114938 162768 115174
rect 162448 114854 162768 114938
rect 162448 114618 162490 114854
rect 162726 114618 162768 114854
rect 162448 114586 162768 114618
rect 193168 115174 193488 115206
rect 193168 114938 193210 115174
rect 193446 114938 193488 115174
rect 193168 114854 193488 114938
rect 193168 114618 193210 114854
rect 193446 114618 193488 114854
rect 193168 114586 193488 114618
rect 223888 115174 224208 115206
rect 223888 114938 223930 115174
rect 224166 114938 224208 115174
rect 223888 114854 224208 114938
rect 223888 114618 223930 114854
rect 224166 114618 224208 114854
rect 223888 114586 224208 114618
rect 254608 115174 254928 115206
rect 254608 114938 254650 115174
rect 254886 114938 254928 115174
rect 254608 114854 254928 114938
rect 254608 114618 254650 114854
rect 254886 114618 254928 114854
rect 254608 114586 254928 114618
rect 285328 115174 285648 115206
rect 285328 114938 285370 115174
rect 285606 114938 285648 115174
rect 285328 114854 285648 114938
rect 285328 114618 285370 114854
rect 285606 114618 285648 114854
rect 285328 114586 285648 114618
rect 316048 115174 316368 115206
rect 316048 114938 316090 115174
rect 316326 114938 316368 115174
rect 316048 114854 316368 114938
rect 316048 114618 316090 114854
rect 316326 114618 316368 114854
rect 316048 114586 316368 114618
rect 346768 115174 347088 115206
rect 346768 114938 346810 115174
rect 347046 114938 347088 115174
rect 346768 114854 347088 114938
rect 346768 114618 346810 114854
rect 347046 114618 347088 114854
rect 346768 114586 347088 114618
rect 54928 111454 55248 111486
rect 54928 111218 54970 111454
rect 55206 111218 55248 111454
rect 54928 111134 55248 111218
rect 54928 110898 54970 111134
rect 55206 110898 55248 111134
rect 54928 110866 55248 110898
rect 85648 111454 85968 111486
rect 85648 111218 85690 111454
rect 85926 111218 85968 111454
rect 85648 111134 85968 111218
rect 85648 110898 85690 111134
rect 85926 110898 85968 111134
rect 85648 110866 85968 110898
rect 116368 111454 116688 111486
rect 116368 111218 116410 111454
rect 116646 111218 116688 111454
rect 116368 111134 116688 111218
rect 116368 110898 116410 111134
rect 116646 110898 116688 111134
rect 116368 110866 116688 110898
rect 147088 111454 147408 111486
rect 147088 111218 147130 111454
rect 147366 111218 147408 111454
rect 147088 111134 147408 111218
rect 147088 110898 147130 111134
rect 147366 110898 147408 111134
rect 147088 110866 147408 110898
rect 177808 111454 178128 111486
rect 177808 111218 177850 111454
rect 178086 111218 178128 111454
rect 177808 111134 178128 111218
rect 177808 110898 177850 111134
rect 178086 110898 178128 111134
rect 177808 110866 178128 110898
rect 208528 111454 208848 111486
rect 208528 111218 208570 111454
rect 208806 111218 208848 111454
rect 208528 111134 208848 111218
rect 208528 110898 208570 111134
rect 208806 110898 208848 111134
rect 208528 110866 208848 110898
rect 239248 111454 239568 111486
rect 239248 111218 239290 111454
rect 239526 111218 239568 111454
rect 239248 111134 239568 111218
rect 239248 110898 239290 111134
rect 239526 110898 239568 111134
rect 239248 110866 239568 110898
rect 269968 111454 270288 111486
rect 269968 111218 270010 111454
rect 270246 111218 270288 111454
rect 269968 111134 270288 111218
rect 269968 110898 270010 111134
rect 270246 110898 270288 111134
rect 269968 110866 270288 110898
rect 300688 111454 301008 111486
rect 300688 111218 300730 111454
rect 300966 111218 301008 111454
rect 300688 111134 301008 111218
rect 300688 110898 300730 111134
rect 300966 110898 301008 111134
rect 300688 110866 301008 110898
rect 331408 111454 331728 111486
rect 331408 111218 331450 111454
rect 331686 111218 331728 111454
rect 331408 111134 331728 111218
rect 331408 110898 331450 111134
rect 331686 110898 331728 111134
rect 331408 110866 331728 110898
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 24208 75454 24528 75486
rect 24208 75218 24250 75454
rect 24486 75218 24528 75454
rect 24208 75134 24528 75218
rect 24208 74898 24250 75134
rect 24486 74898 24528 75134
rect 24208 74866 24528 74898
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 27834 65494 28454 100938
rect 39568 79174 39888 79206
rect 39568 78938 39610 79174
rect 39846 78938 39888 79174
rect 39568 78854 39888 78938
rect 39568 78618 39610 78854
rect 39846 78618 39888 78854
rect 39568 78586 39888 78618
rect 70288 79174 70608 79206
rect 70288 78938 70330 79174
rect 70566 78938 70608 79174
rect 70288 78854 70608 78938
rect 70288 78618 70330 78854
rect 70566 78618 70608 78854
rect 70288 78586 70608 78618
rect 101008 79174 101328 79206
rect 101008 78938 101050 79174
rect 101286 78938 101328 79174
rect 101008 78854 101328 78938
rect 101008 78618 101050 78854
rect 101286 78618 101328 78854
rect 101008 78586 101328 78618
rect 131728 79174 132048 79206
rect 131728 78938 131770 79174
rect 132006 78938 132048 79174
rect 131728 78854 132048 78938
rect 131728 78618 131770 78854
rect 132006 78618 132048 78854
rect 131728 78586 132048 78618
rect 162448 79174 162768 79206
rect 162448 78938 162490 79174
rect 162726 78938 162768 79174
rect 162448 78854 162768 78938
rect 162448 78618 162490 78854
rect 162726 78618 162768 78854
rect 162448 78586 162768 78618
rect 193168 79174 193488 79206
rect 193168 78938 193210 79174
rect 193446 78938 193488 79174
rect 193168 78854 193488 78938
rect 193168 78618 193210 78854
rect 193446 78618 193488 78854
rect 193168 78586 193488 78618
rect 223888 79174 224208 79206
rect 223888 78938 223930 79174
rect 224166 78938 224208 79174
rect 223888 78854 224208 78938
rect 223888 78618 223930 78854
rect 224166 78618 224208 78854
rect 223888 78586 224208 78618
rect 254608 79174 254928 79206
rect 254608 78938 254650 79174
rect 254886 78938 254928 79174
rect 254608 78854 254928 78938
rect 254608 78618 254650 78854
rect 254886 78618 254928 78854
rect 254608 78586 254928 78618
rect 285328 79174 285648 79206
rect 285328 78938 285370 79174
rect 285606 78938 285648 79174
rect 285328 78854 285648 78938
rect 285328 78618 285370 78854
rect 285606 78618 285648 78854
rect 285328 78586 285648 78618
rect 316048 79174 316368 79206
rect 316048 78938 316090 79174
rect 316326 78938 316368 79174
rect 316048 78854 316368 78938
rect 316048 78618 316090 78854
rect 316326 78618 316368 78854
rect 316048 78586 316368 78618
rect 346768 79174 347088 79206
rect 346768 78938 346810 79174
rect 347046 78938 347088 79174
rect 346768 78854 347088 78938
rect 346768 78618 346810 78854
rect 347046 78618 347088 78854
rect 346768 78586 347088 78618
rect 54928 75454 55248 75486
rect 54928 75218 54970 75454
rect 55206 75218 55248 75454
rect 54928 75134 55248 75218
rect 54928 74898 54970 75134
rect 55206 74898 55248 75134
rect 54928 74866 55248 74898
rect 85648 75454 85968 75486
rect 85648 75218 85690 75454
rect 85926 75218 85968 75454
rect 85648 75134 85968 75218
rect 85648 74898 85690 75134
rect 85926 74898 85968 75134
rect 85648 74866 85968 74898
rect 116368 75454 116688 75486
rect 116368 75218 116410 75454
rect 116646 75218 116688 75454
rect 116368 75134 116688 75218
rect 116368 74898 116410 75134
rect 116646 74898 116688 75134
rect 116368 74866 116688 74898
rect 147088 75454 147408 75486
rect 147088 75218 147130 75454
rect 147366 75218 147408 75454
rect 147088 75134 147408 75218
rect 147088 74898 147130 75134
rect 147366 74898 147408 75134
rect 147088 74866 147408 74898
rect 177808 75454 178128 75486
rect 177808 75218 177850 75454
rect 178086 75218 178128 75454
rect 177808 75134 178128 75218
rect 177808 74898 177850 75134
rect 178086 74898 178128 75134
rect 177808 74866 178128 74898
rect 208528 75454 208848 75486
rect 208528 75218 208570 75454
rect 208806 75218 208848 75454
rect 208528 75134 208848 75218
rect 208528 74898 208570 75134
rect 208806 74898 208848 75134
rect 208528 74866 208848 74898
rect 239248 75454 239568 75486
rect 239248 75218 239290 75454
rect 239526 75218 239568 75454
rect 239248 75134 239568 75218
rect 239248 74898 239290 75134
rect 239526 74898 239568 75134
rect 239248 74866 239568 74898
rect 269968 75454 270288 75486
rect 269968 75218 270010 75454
rect 270246 75218 270288 75454
rect 269968 75134 270288 75218
rect 269968 74898 270010 75134
rect 270246 74898 270288 75134
rect 269968 74866 270288 74898
rect 300688 75454 301008 75486
rect 300688 75218 300730 75454
rect 300966 75218 301008 75454
rect 300688 75134 301008 75218
rect 300688 74898 300730 75134
rect 300966 74898 301008 75134
rect 300688 74866 301008 74898
rect 331408 75454 331728 75486
rect 331408 75218 331450 75454
rect 331686 75218 331728 75454
rect 331408 75134 331728 75218
rect 331408 74898 331450 75134
rect 331686 74898 331728 75134
rect 331408 74866 331728 74898
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 22139 49604 22205 49605
rect 22139 49540 22140 49604
rect 22204 49540 22205 49604
rect 22139 49539 22205 49540
rect 22142 46477 22202 49539
rect 22323 49468 22389 49469
rect 22323 49404 22324 49468
rect 22388 49404 22389 49468
rect 22323 49403 22389 49404
rect 22139 46476 22205 46477
rect 22139 46412 22140 46476
rect 22204 46412 22205 46476
rect 22139 46411 22205 46412
rect 22326 46341 22386 49403
rect 22323 46340 22389 46341
rect 22323 46276 22324 46340
rect 22388 46276 22389 46340
rect 22323 46275 22389 46276
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 25774 24734 45068
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 39454 38414 49367
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 43174 42134 49367
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 46894 45854 49367
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 49367
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 49367
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 49367
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 49367
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 29494 64454 49367
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 49367
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 49367
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 49367
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 49367
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 49367
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 49367
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 25774 96734 49367
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 29494 100454 49367
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 39454 110414 49367
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 43174 114134 49367
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 46894 117854 49367
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 49367
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 49367
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 49367
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 25774 132734 49367
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 29494 136454 49367
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 39454 146414 49367
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 43174 150134 49367
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 46894 153854 49367
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 14614 157574 49367
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 18334 161294 49367
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 22054 165014 49367
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 25774 168734 49367
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 29494 172454 49367
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 39454 182414 49367
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 43174 186134 49367
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 46894 189854 49367
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 14614 193574 45068
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 18334 197294 49367
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 22054 201014 49367
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 25774 204734 49367
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 29494 208454 49367
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 39454 218414 49367
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 43174 222134 49367
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 46894 225854 49367
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 14614 229574 49367
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 49367
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 22054 237014 49367
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 49367
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 29494 244454 49367
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 49367
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 43174 258134 49367
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 46894 261854 49367
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 49367
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 49367
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 49367
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 49367
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 49367
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 49367
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 43174 294134 49367
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 46894 297854 49367
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 45068
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 49367
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 49367
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 49367
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 45068
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 49367
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 43174 330134 49367
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 46894 333854 49367
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 49367
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 49367
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 49367
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 49367
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 49367
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 404417 327454 404737 327486
rect 404417 327218 404459 327454
rect 404695 327218 404737 327454
rect 404417 327134 404737 327218
rect 404417 326898 404459 327134
rect 404695 326898 404737 327134
rect 404417 326866 404737 326898
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 298894 405854 334338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 407890 331174 408210 331206
rect 407890 330938 407932 331174
rect 408168 330938 408210 331174
rect 407890 330854 408210 330938
rect 407890 330618 407932 330854
rect 408168 330618 408210 330854
rect 407890 330586 408210 330618
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 302614 409574 338058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 411363 327454 411683 327486
rect 411363 327218 411405 327454
rect 411641 327218 411683 327454
rect 411363 327134 411683 327218
rect 411363 326898 411405 327134
rect 411641 326898 411683 327134
rect 411363 326866 411683 326898
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 306334 413294 341778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 414836 331174 415156 331206
rect 414836 330938 414878 331174
rect 415114 330938 415156 331174
rect 414836 330854 415156 330938
rect 414836 330618 414878 330854
rect 415114 330618 415156 330854
rect 414836 330586 415156 330618
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 416394 310054 417014 345498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 444412 424454 460938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442833 434414 470898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 444412 438134 474618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 447731 700364 447797 700365
rect 447731 700300 447732 700364
rect 447796 700300 447797 700364
rect 447731 700299 447797 700300
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444235 690708 444301 690709
rect 444235 690644 444236 690708
rect 444300 690644 444301 690708
rect 444235 690643 444301 690644
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442833 441854 478338
rect 426624 439174 426944 439206
rect 426624 438938 426666 439174
rect 426902 438938 426944 439174
rect 426624 438854 426944 438938
rect 426624 438618 426666 438854
rect 426902 438618 426944 438854
rect 426624 438586 426944 438618
rect 432305 439174 432625 439206
rect 432305 438938 432347 439174
rect 432583 438938 432625 439174
rect 432305 438854 432625 438938
rect 432305 438618 432347 438854
rect 432583 438618 432625 438854
rect 432305 438586 432625 438618
rect 437986 439174 438306 439206
rect 437986 438938 438028 439174
rect 438264 438938 438306 439174
rect 437986 438854 438306 438938
rect 437986 438618 438028 438854
rect 438264 438618 438306 438854
rect 437986 438586 438306 438618
rect 443667 439174 443987 439206
rect 443667 438938 443709 439174
rect 443945 438938 443987 439174
rect 443667 438854 443987 438938
rect 443667 438618 443709 438854
rect 443945 438618 443987 438854
rect 443667 438586 443987 438618
rect 423784 435454 424104 435486
rect 423784 435218 423826 435454
rect 424062 435218 424104 435454
rect 423784 435134 424104 435218
rect 423784 434898 423826 435134
rect 424062 434898 424104 435134
rect 423784 434866 424104 434898
rect 429465 435454 429785 435486
rect 429465 435218 429507 435454
rect 429743 435218 429785 435454
rect 429465 435134 429785 435218
rect 429465 434898 429507 435134
rect 429743 434898 429785 435134
rect 429465 434866 429785 434898
rect 435146 435454 435466 435486
rect 435146 435218 435188 435454
rect 435424 435218 435466 435454
rect 435146 435134 435466 435218
rect 435146 434898 435188 435134
rect 435424 434898 435466 435134
rect 435146 434866 435466 434898
rect 440827 435454 441147 435486
rect 440827 435218 440869 435454
rect 441105 435218 441147 435454
rect 440827 435134 441147 435218
rect 440827 434898 440869 435134
rect 441105 434898 441147 435134
rect 440827 434866 441147 434898
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 418309 327454 418629 327486
rect 418309 327218 418351 327454
rect 418587 327218 418629 327454
rect 418309 327134 418629 327218
rect 418309 326898 418351 327134
rect 418587 326898 418629 327134
rect 418309 326866 418629 326898
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 157249 417014 165498
rect 420114 313774 420734 349218
rect 423834 389494 424454 420068
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 421051 334524 421117 334525
rect 421051 334460 421052 334524
rect 421116 334460 421117 334524
rect 421051 334459 421117 334460
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 157249 420734 169218
rect 421054 162757 421114 334459
rect 421782 331174 422102 331206
rect 421782 330938 421824 331174
rect 422060 330938 422102 331174
rect 421782 330854 422102 330938
rect 421782 330618 421824 330854
rect 422060 330618 422102 330854
rect 421782 330586 422102 330618
rect 423834 317494 424454 352938
rect 433794 399454 434414 422599
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 425835 335476 425901 335477
rect 425835 335412 425836 335476
rect 425900 335412 425901 335476
rect 425835 335411 425901 335412
rect 425838 333029 425898 335411
rect 428411 334524 428477 334525
rect 428411 334460 428412 334524
rect 428476 334460 428477 334524
rect 428411 334459 428477 334460
rect 425835 333028 425901 333029
rect 425835 332964 425836 333028
rect 425900 332964 425901 333028
rect 425835 332963 425901 332964
rect 425255 327454 425575 327486
rect 425255 327218 425297 327454
rect 425533 327218 425575 327454
rect 425255 327134 425575 327218
rect 425255 326898 425297 327134
rect 425533 326898 425575 327134
rect 425255 326866 425575 326898
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 421051 162756 421117 162757
rect 421051 162692 421052 162756
rect 421116 162692 421117 162756
rect 421051 162691 421117 162692
rect 423834 157249 424454 172938
rect 425838 162757 425898 332963
rect 428414 162757 428474 334459
rect 428728 331174 429048 331206
rect 428728 330938 428770 331174
rect 429006 330938 429048 331174
rect 428728 330854 429048 330938
rect 428728 330618 428770 330854
rect 429006 330618 429048 330854
rect 428728 330586 429048 330618
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 425835 162756 425901 162757
rect 425835 162692 425836 162756
rect 425900 162692 425901 162756
rect 425835 162691 425901 162692
rect 428411 162756 428477 162757
rect 428411 162692 428412 162756
rect 428476 162692 428477 162756
rect 428411 162691 428477 162692
rect 433794 157249 434414 182898
rect 437514 403174 438134 420068
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 157249 438134 186618
rect 441234 406894 441854 422599
rect 444051 421972 444117 421973
rect 444051 421908 444052 421972
rect 444116 421908 444117 421972
rect 444051 421907 444117 421908
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 444054 321197 444114 421907
rect 444051 321196 444117 321197
rect 444051 321132 444052 321196
rect 444116 321132 444117 321196
rect 444051 321131 444117 321132
rect 444238 319837 444298 690643
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444235 319836 444301 319837
rect 444235 319772 444236 319836
rect 444300 319772 444301 319836
rect 444235 319771 444301 319772
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 157249 441854 190338
rect 444954 302614 445574 338058
rect 447734 321877 447794 700299
rect 448674 666334 449294 708122
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 449571 700500 449637 700501
rect 449571 700436 449572 700500
rect 449636 700436 449637 700500
rect 449571 700435 449637 700436
rect 451779 700500 451845 700501
rect 451779 700436 451780 700500
rect 451844 700436 451845 700500
rect 451779 700435 451845 700436
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448283 516220 448349 516221
rect 448283 516156 448284 516220
rect 448348 516156 448349 516220
rect 448283 516155 448349 516156
rect 448286 496093 448346 516155
rect 448283 496092 448349 496093
rect 448283 496028 448284 496092
rect 448348 496028 448349 496092
rect 448283 496027 448349 496028
rect 448286 329221 448346 496027
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448283 329220 448349 329221
rect 448283 329156 448284 329220
rect 448348 329156 448349 329220
rect 448283 329155 448349 329156
rect 447731 321876 447797 321877
rect 447731 321812 447732 321876
rect 447796 321812 447797 321876
rect 447731 321811 447797 321812
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 159644 445574 194058
rect 448674 306334 449294 341778
rect 449574 321333 449634 700435
rect 450491 692068 450557 692069
rect 450491 692004 450492 692068
rect 450556 692004 450557 692068
rect 450491 692003 450557 692004
rect 449571 321332 449637 321333
rect 449571 321268 449572 321332
rect 449636 321268 449637 321332
rect 449571 321267 449637 321268
rect 450494 319565 450554 692003
rect 450675 689348 450741 689349
rect 450675 689284 450676 689348
rect 450740 689284 450741 689348
rect 450675 689283 450741 689284
rect 450678 319973 450738 689283
rect 451782 420205 451842 700435
rect 452394 670054 453014 709082
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 455091 700364 455157 700365
rect 455091 700300 455092 700364
rect 455156 700300 455157 700364
rect 455091 700299 455157 700300
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 453251 669900 453317 669901
rect 453251 669836 453252 669900
rect 453316 669836 453317 669900
rect 453251 669835 453317 669836
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 517884 453014 525498
rect 452163 507454 452483 507486
rect 452163 507218 452205 507454
rect 452441 507218 452483 507454
rect 452163 507134 452483 507218
rect 452163 506898 452205 507134
rect 452441 506898 452483 507134
rect 452163 506866 452483 506898
rect 452394 490054 453014 500068
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 451779 420204 451845 420205
rect 451779 420140 451780 420204
rect 451844 420140 451845 420204
rect 451779 420139 451845 420140
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 453254 387701 453314 669835
rect 453382 511174 453702 511206
rect 453382 510938 453424 511174
rect 453660 510938 453702 511174
rect 453382 510854 453702 510938
rect 453382 510618 453424 510854
rect 453660 510618 453702 510854
rect 453382 510586 453702 510618
rect 454601 507454 454921 507486
rect 454601 507218 454643 507454
rect 454879 507218 454921 507454
rect 454601 507134 454921 507218
rect 454601 506898 454643 507134
rect 454879 506898 454921 507134
rect 454601 506866 454921 506898
rect 455094 422925 455154 700299
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 668393 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 668393 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 668393 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 668393 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 668393 481574 698058
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 668393 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 668393 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 668393 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 668393 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 668393 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 668393 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 668393 517574 698058
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 527219 699820 527285 699821
rect 527219 699756 527220 699820
rect 527284 699756 527285 699820
rect 527219 699755 527285 699756
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 458035 665548 458101 665549
rect 458035 665484 458036 665548
rect 458100 665484 458101 665548
rect 458035 665483 458101 665484
rect 457851 663100 457917 663101
rect 457851 663036 457852 663100
rect 457916 663036 457917 663100
rect 457851 663035 457917 663036
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 517884 456734 529218
rect 457854 519485 457914 663035
rect 457851 519484 457917 519485
rect 457851 519420 457852 519484
rect 457916 519420 457917 519484
rect 457851 519419 457917 519420
rect 458038 517581 458098 665483
rect 479568 655174 479888 655206
rect 479568 654938 479610 655174
rect 479846 654938 479888 655174
rect 479568 654854 479888 654938
rect 479568 654618 479610 654854
rect 479846 654618 479888 654854
rect 479568 654586 479888 654618
rect 510288 655174 510608 655206
rect 510288 654938 510330 655174
rect 510566 654938 510608 655174
rect 510288 654854 510608 654938
rect 510288 654618 510330 654854
rect 510566 654618 510608 654854
rect 510288 654586 510608 654618
rect 464208 651454 464528 651486
rect 464208 651218 464250 651454
rect 464486 651218 464528 651454
rect 464208 651134 464528 651218
rect 464208 650898 464250 651134
rect 464486 650898 464528 651134
rect 464208 650866 464528 650898
rect 494928 651454 495248 651486
rect 494928 651218 494970 651454
rect 495206 651218 495248 651454
rect 494928 651134 495248 651218
rect 494928 650898 494970 651134
rect 495206 650898 495248 651134
rect 494928 650866 495248 650898
rect 458955 636172 459021 636173
rect 458955 636108 458956 636172
rect 459020 636108 459021 636172
rect 458955 636107 459021 636108
rect 458035 517580 458101 517581
rect 458035 517516 458036 517580
rect 458100 517516 458101 517580
rect 458035 517515 458101 517516
rect 455820 511174 456140 511206
rect 455820 510938 455862 511174
rect 456098 510938 456140 511174
rect 455820 510854 456140 510938
rect 455820 510618 455862 510854
rect 456098 510618 456140 510854
rect 455820 510586 456140 510618
rect 458258 511174 458578 511206
rect 458258 510938 458300 511174
rect 458536 510938 458578 511174
rect 458258 510854 458578 510938
rect 458258 510618 458300 510854
rect 458536 510618 458578 510854
rect 458258 510586 458578 510618
rect 457039 507454 457359 507486
rect 457039 507218 457081 507454
rect 457317 507218 457359 507454
rect 457039 507134 457359 507218
rect 457039 506898 457081 507134
rect 457317 506898 457359 507134
rect 457039 506866 457359 506898
rect 456114 493774 456734 500068
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 455091 422924 455157 422925
rect 455091 422860 455092 422924
rect 455156 422860 455157 422924
rect 455091 422859 455157 422860
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 453251 387700 453317 387701
rect 453251 387636 453252 387700
rect 453316 387636 453317 387700
rect 453251 387635 453317 387636
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 456114 385774 456734 421218
rect 458958 393957 459018 636107
rect 524394 634054 525014 669498
rect 525648 651454 525968 651486
rect 525648 651218 525690 651454
rect 525926 651218 525968 651454
rect 525648 651134 525968 651218
rect 525648 650898 525690 651134
rect 525926 650898 525968 651134
rect 525648 650866 525968 650898
rect 524394 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 525014 634054
rect 524394 633734 525014 633818
rect 459139 633724 459205 633725
rect 459139 633660 459140 633724
rect 459204 633660 459205 633724
rect 459139 633659 459205 633660
rect 458955 393956 459021 393957
rect 458955 393892 458956 393956
rect 459020 393892 459021 393956
rect 458955 393891 459021 393892
rect 459142 392597 459202 633659
rect 524394 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 525014 633734
rect 479568 619174 479888 619206
rect 479568 618938 479610 619174
rect 479846 618938 479888 619174
rect 479568 618854 479888 618938
rect 479568 618618 479610 618854
rect 479846 618618 479888 618854
rect 479568 618586 479888 618618
rect 510288 619174 510608 619206
rect 510288 618938 510330 619174
rect 510566 618938 510608 619174
rect 510288 618854 510608 618938
rect 510288 618618 510330 618854
rect 510566 618618 510608 618854
rect 510288 618586 510608 618618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 478827 599588 478893 599589
rect 478827 599524 478828 599588
rect 478892 599524 478893 599588
rect 478827 599523 478893 599524
rect 459834 569494 460454 598927
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 517884 460454 532938
rect 469794 579454 470414 598927
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 460696 511174 461016 511206
rect 460696 510938 460738 511174
rect 460974 510938 461016 511174
rect 460696 510854 461016 510938
rect 460696 510618 460738 510854
rect 460974 510618 461016 510854
rect 460696 510586 461016 510618
rect 459477 507454 459797 507486
rect 459477 507218 459519 507454
rect 459755 507218 459797 507454
rect 459477 507134 459797 507218
rect 459477 506898 459519 507134
rect 459755 506898 459797 507134
rect 459477 506866 459797 506898
rect 469794 507454 470414 542898
rect 473514 583174 474134 598927
rect 474411 598228 474477 598229
rect 474411 598164 474412 598228
rect 474476 598164 474477 598228
rect 474411 598163 474477 598164
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 472019 522340 472085 522341
rect 472019 522276 472020 522340
rect 472084 522276 472085 522340
rect 472019 522275 472085 522276
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 459834 497494 460454 500068
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459139 392596 459205 392597
rect 459139 392532 459140 392596
rect 459204 392532 459205 392596
rect 459139 392531 459205 392532
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 454208 363454 454528 363486
rect 454208 363218 454250 363454
rect 454486 363218 454528 363454
rect 454208 363134 454528 363218
rect 454208 362898 454250 363134
rect 454486 362898 454528 363134
rect 454208 362866 454528 362898
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 450675 319972 450741 319973
rect 450675 319908 450676 319972
rect 450740 319908 450741 319972
rect 450675 319907 450741 319908
rect 450491 319564 450557 319565
rect 450491 319500 450492 319564
rect 450556 319500 450557 319564
rect 450491 319499 450557 319500
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 429568 151174 429888 151206
rect 429568 150938 429610 151174
rect 429846 150938 429888 151174
rect 429568 150854 429888 150938
rect 429568 150618 429610 150854
rect 429846 150618 429888 150854
rect 429568 150586 429888 150618
rect 414208 147454 414528 147486
rect 414208 147218 414250 147454
rect 414486 147218 414528 147454
rect 414208 147134 414528 147218
rect 414208 146898 414250 147134
rect 414486 146898 414528 147134
rect 414208 146866 414528 146898
rect 444928 147454 445248 147486
rect 444928 147218 444970 147454
rect 445206 147218 445248 147454
rect 444928 147134 445248 147218
rect 444928 146898 444970 147134
rect 445206 146898 445248 147134
rect 444928 146866 445248 146898
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 94054 417014 127767
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 97774 420734 127767
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 101494 424454 127767
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 111454 434414 127767
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 115174 438134 127767
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 118894 441854 127767
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 86614 445574 120068
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 310054 453014 345498
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 454208 327454 454528 327486
rect 454208 327218 454250 327454
rect 454486 327218 454528 327454
rect 454208 327134 454528 327218
rect 454208 326898 454250 327134
rect 454486 326898 454528 327134
rect 454208 326866 454528 326898
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 313774 456734 349218
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 385580 470414 398898
rect 472022 389061 472082 522275
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 453692 474134 474618
rect 473416 435454 473736 435486
rect 473416 435218 473458 435454
rect 473694 435218 473736 435454
rect 473416 435134 473736 435218
rect 473416 434898 473458 435134
rect 473694 434898 473736 435134
rect 473416 434866 473736 434898
rect 474414 389061 474474 598163
rect 474779 597004 474845 597005
rect 474779 596940 474780 597004
rect 474844 596940 474845 597004
rect 474779 596939 474845 596940
rect 474782 389061 474842 596939
rect 476435 596868 476501 596869
rect 476435 596804 476436 596868
rect 476500 596804 476501 596868
rect 476435 596803 476501 596804
rect 475888 439174 476208 439206
rect 475888 438938 475930 439174
rect 476166 438938 476208 439174
rect 475888 438854 476208 438938
rect 475888 438618 475930 438854
rect 476166 438618 476208 438854
rect 475888 438586 476208 438618
rect 476438 389061 476498 596803
rect 477234 586894 477854 598927
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 478361 435454 478681 435486
rect 478361 435218 478403 435454
rect 478639 435218 478681 435454
rect 478361 435134 478681 435218
rect 478361 434898 478403 435134
rect 478639 434898 478681 435134
rect 478361 434866 478681 434898
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 472019 389060 472085 389061
rect 472019 388996 472020 389060
rect 472084 388996 472085 389060
rect 472019 388995 472085 388996
rect 474411 389060 474477 389061
rect 474411 388996 474412 389060
rect 474476 388996 474477 389060
rect 474411 388995 474477 388996
rect 474779 389060 474845 389061
rect 474779 388996 474780 389060
rect 474844 388996 474845 389060
rect 474779 388995 474845 388996
rect 476435 389060 476501 389061
rect 476435 388996 476436 389060
rect 476500 388996 476501 389060
rect 476435 388995 476501 388996
rect 477234 385225 477854 406338
rect 478830 389061 478890 599523
rect 480954 590614 481574 598927
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 484674 594334 485294 598927
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 517884 485294 521778
rect 488394 598054 489014 598927
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 517884 489014 525498
rect 492114 565774 492734 598927
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 483382 511174 483702 511206
rect 483382 510938 483424 511174
rect 483660 510938 483702 511174
rect 483382 510854 483702 510938
rect 483382 510618 483424 510854
rect 483660 510618 483702 510854
rect 483382 510586 483702 510618
rect 485820 511174 486140 511206
rect 485820 510938 485862 511174
rect 486098 510938 486140 511174
rect 485820 510854 486140 510938
rect 485820 510618 485862 510854
rect 486098 510618 486140 510854
rect 485820 510586 486140 510618
rect 488258 511174 488578 511206
rect 488258 510938 488300 511174
rect 488536 510938 488578 511174
rect 488258 510854 488578 510938
rect 488258 510618 488300 510854
rect 488536 510618 488578 510854
rect 488258 510586 488578 510618
rect 490696 511174 491016 511206
rect 490696 510938 490738 511174
rect 490974 510938 491016 511174
rect 490696 510854 491016 510938
rect 490696 510618 490738 510854
rect 490974 510618 491016 510854
rect 490696 510586 491016 510618
rect 482163 507454 482483 507486
rect 482163 507218 482205 507454
rect 482441 507218 482483 507454
rect 482163 507134 482483 507218
rect 482163 506898 482205 507134
rect 482441 506898 482483 507134
rect 482163 506866 482483 506898
rect 484601 507454 484921 507486
rect 484601 507218 484643 507454
rect 484879 507218 484921 507454
rect 484601 507134 484921 507218
rect 484601 506898 484643 507134
rect 484879 506898 484921 507134
rect 484601 506866 484921 506898
rect 487039 507454 487359 507486
rect 487039 507218 487081 507454
rect 487317 507218 487359 507454
rect 487039 507134 487359 507218
rect 487039 506898 487081 507134
rect 487317 506898 487359 507134
rect 487039 506866 487359 506898
rect 489477 507454 489797 507486
rect 489477 507218 489519 507454
rect 489755 507218 489797 507454
rect 489477 507134 489797 507218
rect 489477 506898 489519 507134
rect 489755 506898 489797 507134
rect 489477 506866 489797 506898
rect 483059 496908 483125 496909
rect 483059 496844 483060 496908
rect 483124 496844 483125 496908
rect 483059 496843 483125 496844
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 453692 481574 482058
rect 480833 439174 481153 439206
rect 480833 438938 480875 439174
rect 481111 438938 481153 439174
rect 480833 438854 481153 438938
rect 480833 438618 480875 438854
rect 481111 438618 481153 438854
rect 480833 438586 481153 438618
rect 478827 389060 478893 389061
rect 478827 388996 478828 389060
rect 478892 388996 478893 389060
rect 478827 388995 478893 388996
rect 483062 387157 483122 496843
rect 484674 486334 485294 500068
rect 486371 496908 486437 496909
rect 486371 496844 486372 496908
rect 486436 496844 486437 496908
rect 486371 496843 486437 496844
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 483306 435454 483626 435486
rect 483306 435218 483348 435454
rect 483584 435218 483626 435454
rect 483306 435134 483626 435218
rect 483306 434898 483348 435134
rect 483584 434898 483626 435134
rect 483306 434866 483626 434898
rect 484674 414334 485294 449778
rect 485778 439174 486098 439206
rect 485778 438938 485820 439174
rect 486056 438938 486098 439174
rect 485778 438854 486098 438938
rect 485778 438618 485820 438854
rect 486056 438618 486098 438854
rect 485778 438586 486098 438618
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 483059 387156 483125 387157
rect 483059 387092 483060 387156
rect 483124 387092 483125 387156
rect 483059 387091 483125 387092
rect 484674 385580 485294 413778
rect 486374 387021 486434 496843
rect 488394 490054 489014 500068
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454007 489014 489498
rect 487107 453932 487173 453933
rect 487107 453868 487108 453932
rect 487172 453868 487173 453932
rect 487107 453867 487173 453868
rect 486371 387020 486437 387021
rect 486371 386956 486372 387020
rect 486436 386956 486437 387020
rect 486371 386955 486437 386956
rect 487110 385661 487170 453867
rect 488394 453771 488426 454007
rect 488662 453771 488746 454007
rect 488982 453771 489014 454007
rect 488394 453692 489014 453771
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 490723 439174 491043 439206
rect 490723 438938 490765 439174
rect 491001 438938 491043 439174
rect 490723 438854 491043 438938
rect 490723 438618 490765 438854
rect 491001 438618 491043 438854
rect 490723 438586 491043 438618
rect 488251 435454 488571 435486
rect 488251 435218 488293 435454
rect 488529 435218 488571 435454
rect 488251 435134 488571 435218
rect 488251 434898 488293 435134
rect 488529 434898 488571 435134
rect 488251 434866 488571 434898
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 487107 385660 487173 385661
rect 487107 385596 487108 385660
rect 487172 385596 487173 385660
rect 487107 385595 487173 385596
rect 492114 385225 492734 421218
rect 495834 569494 496454 598927
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 469568 367174 469888 367206
rect 469568 366938 469610 367174
rect 469846 366938 469888 367174
rect 469568 366854 469888 366938
rect 469568 366618 469610 366854
rect 469846 366618 469888 366854
rect 469568 366586 469888 366618
rect 484928 363454 485248 363486
rect 484928 363218 484970 363454
rect 485206 363218 485248 363454
rect 484928 363134 485248 363218
rect 484928 362898 484970 363134
rect 485206 362898 485248 363134
rect 484928 362866 485248 362898
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 495834 353494 496454 388938
rect 505794 579454 506414 598927
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 500288 367174 500608 367206
rect 500288 366938 500330 367174
rect 500566 366938 500608 367174
rect 500288 366854 500608 366938
rect 500288 366618 500330 366854
rect 500566 366618 500608 366854
rect 500288 366586 500608 366618
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 469568 331174 469888 331206
rect 469568 330938 469610 331174
rect 469846 330938 469888 331174
rect 469568 330854 469888 330938
rect 469568 330618 469610 330854
rect 469846 330618 469888 330854
rect 469568 330586 469888 330618
rect 484928 327454 485248 327486
rect 484928 327218 484970 327454
rect 485206 327218 485248 327454
rect 484928 327134 485248 327218
rect 484928 326898 484970 327134
rect 485206 326898 485248 327134
rect 484928 326866 485248 326898
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 458955 317116 459021 317117
rect 458955 317052 458956 317116
rect 459020 317052 459021 317116
rect 458955 317051 459021 317052
rect 458771 316844 458837 316845
rect 458771 316780 458772 316844
rect 458836 316780 458837 316844
rect 458771 316779 458837 316780
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 456114 205774 456734 241218
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 458774 39405 458834 316779
rect 458771 39404 458837 39405
rect 458771 39340 458772 39404
rect 458836 39340 458837 39404
rect 458771 39339 458837 39340
rect 458958 39269 459018 317051
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 477234 298894 477854 322287
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 259417 477854 262338
rect 480954 302614 481574 322287
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 259417 481574 266058
rect 484674 306334 485294 322068
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 259417 485294 269778
rect 488394 310054 489014 322287
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 259417 489014 273498
rect 492114 313774 492734 322287
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 259417 492734 277218
rect 495834 317494 496454 352938
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 500288 331174 500608 331206
rect 500288 330938 500330 331174
rect 500566 330938 500608 331174
rect 500288 330854 500608 330938
rect 500288 330618 500330 330854
rect 500566 330618 500608 330854
rect 500288 330586 500608 330618
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 259417 496454 280938
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 509514 583174 510134 598927
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 513234 586894 513854 598927
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 511027 333572 511093 333573
rect 511027 333508 511028 333572
rect 511092 333508 511093 333572
rect 511027 333507 511093 333508
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 508451 322828 508517 322829
rect 508451 322764 508452 322828
rect 508516 322764 508517 322828
rect 508451 322763 508517 322764
rect 508454 291821 508514 322763
rect 509187 322692 509253 322693
rect 509187 322690 509188 322692
rect 509006 322630 509188 322690
rect 509006 316709 509066 322630
rect 509187 322628 509188 322630
rect 509252 322628 509253 322692
rect 509187 322627 509253 322628
rect 509003 316708 509069 316709
rect 509003 316644 509004 316708
rect 509068 316644 509069 316708
rect 509003 316643 509069 316644
rect 509514 295174 510134 330618
rect 510843 329764 510909 329765
rect 510843 329700 510844 329764
rect 510908 329700 510909 329764
rect 510843 329699 510909 329700
rect 510475 328132 510541 328133
rect 510475 328068 510476 328132
rect 510540 328068 510541 328132
rect 510475 328067 510541 328068
rect 510478 302837 510538 328067
rect 510659 326500 510725 326501
rect 510659 326436 510660 326500
rect 510724 326436 510725 326500
rect 510659 326435 510725 326436
rect 510662 324461 510722 326435
rect 510659 324460 510725 324461
rect 510659 324396 510660 324460
rect 510724 324396 510725 324460
rect 510659 324395 510725 324396
rect 510659 324324 510725 324325
rect 510659 324260 510660 324324
rect 510724 324260 510725 324324
rect 510659 324259 510725 324260
rect 510662 316981 510722 324259
rect 510659 316980 510725 316981
rect 510659 316916 510660 316980
rect 510724 316916 510725 316980
rect 510659 316915 510725 316916
rect 510475 302836 510541 302837
rect 510475 302772 510476 302836
rect 510540 302772 510541 302836
rect 510475 302771 510541 302772
rect 510846 300525 510906 329699
rect 510843 300524 510909 300525
rect 510843 300460 510844 300524
rect 510908 300460 510909 300524
rect 510843 300459 510909 300460
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 511030 294813 511090 333507
rect 511211 324460 511277 324461
rect 511211 324396 511212 324460
rect 511276 324396 511277 324460
rect 511211 324395 511277 324396
rect 511214 317253 511274 324395
rect 511211 317252 511277 317253
rect 511211 317188 511212 317252
rect 511276 317188 511277 317252
rect 511211 317187 511277 317188
rect 513234 298894 513854 334338
rect 516954 590614 517574 598927
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 515075 333028 515141 333029
rect 515075 332964 515076 333028
rect 515140 332964 515141 333028
rect 515075 332963 515141 332964
rect 514707 331396 514773 331397
rect 514707 331332 514708 331396
rect 514772 331332 514773 331396
rect 514707 331331 514773 331332
rect 514155 328676 514221 328677
rect 514155 328612 514156 328676
rect 514220 328612 514221 328676
rect 514155 328611 514221 328612
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 511027 294812 511093 294813
rect 511027 294748 511028 294812
rect 511092 294748 511093 294812
rect 511027 294747 511093 294748
rect 508451 291820 508517 291821
rect 508451 291756 508452 291820
rect 508516 291756 508517 291820
rect 508451 291755 508517 291756
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 259417 506414 290898
rect 509514 259417 510134 294618
rect 513234 262894 513854 298338
rect 514158 297397 514218 328611
rect 514339 324868 514405 324869
rect 514339 324804 514340 324868
rect 514404 324804 514405 324868
rect 514339 324803 514405 324804
rect 514342 300389 514402 324803
rect 514339 300388 514405 300389
rect 514339 300324 514340 300388
rect 514404 300324 514405 300388
rect 514339 300323 514405 300324
rect 514710 300253 514770 331331
rect 514891 327044 514957 327045
rect 514891 326980 514892 327044
rect 514956 326980 514957 327044
rect 514891 326979 514957 326980
rect 514707 300252 514773 300253
rect 514707 300188 514708 300252
rect 514772 300188 514773 300252
rect 514707 300187 514773 300188
rect 514894 300117 514954 326979
rect 515078 317117 515138 332963
rect 516179 327588 516245 327589
rect 516179 327524 516180 327588
rect 516244 327524 516245 327588
rect 516179 327523 516245 327524
rect 515075 317116 515141 317117
rect 515075 317052 515076 317116
rect 515140 317052 515141 317116
rect 515075 317051 515141 317052
rect 514891 300116 514957 300117
rect 514891 300052 514892 300116
rect 514956 300052 514957 300116
rect 514891 300051 514957 300052
rect 514155 297396 514221 297397
rect 514155 297332 514156 297396
rect 514220 297332 514221 297396
rect 514155 297331 514221 297332
rect 516182 294541 516242 327523
rect 516954 302614 517574 338058
rect 520674 594334 521294 598927
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 518019 335204 518085 335205
rect 518019 335140 518020 335204
rect 518084 335140 518085 335204
rect 518019 335139 518085 335140
rect 517835 330852 517901 330853
rect 517835 330788 517836 330852
rect 517900 330788 517901 330852
rect 517835 330787 517901 330788
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516179 294540 516245 294541
rect 516179 294476 516180 294540
rect 516244 294476 516245 294540
rect 516179 294475 516245 294476
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 259417 513854 262338
rect 516954 266614 517574 302058
rect 517838 289101 517898 330787
rect 518022 294677 518082 335139
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 518019 294676 518085 294677
rect 518019 294612 518020 294676
rect 518084 294612 518085 294676
rect 518019 294611 518085 294612
rect 517835 289100 517901 289101
rect 517835 289036 517836 289100
rect 517900 289036 517901 289100
rect 517835 289035 517901 289036
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 259417 517574 266058
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 259417 521294 269778
rect 524394 598054 525014 633498
rect 525648 615454 525968 615486
rect 525648 615218 525690 615454
rect 525926 615218 525968 615454
rect 525648 615134 525968 615218
rect 525648 614898 525690 615134
rect 525926 614898 525968 615134
rect 525648 614866 525968 614898
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 527222 465765 527282 699755
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 637774 528734 673218
rect 528114 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 528734 637774
rect 528114 637454 528734 637538
rect 528114 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 528734 637454
rect 528114 601774 528734 637218
rect 528114 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 528734 601774
rect 528114 601454 528734 601538
rect 528114 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 528734 601454
rect 528114 565774 528734 601218
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 527219 465764 527285 465765
rect 527219 465700 527220 465764
rect 527284 465700 527285 465764
rect 527219 465699 527285 465700
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 525164 435454 525484 435486
rect 525164 435218 525206 435454
rect 525442 435218 525484 435454
rect 525164 435134 525484 435218
rect 525164 434898 525206 435134
rect 525442 434898 525484 435134
rect 525164 434866 525484 434898
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 259417 525014 273498
rect 528114 421774 528734 457218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 641494 532454 676938
rect 531834 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 532454 641494
rect 531834 641174 532454 641258
rect 531834 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 532454 641174
rect 531834 605494 532454 640938
rect 531834 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 532454 605494
rect 531834 605174 532454 605258
rect 531834 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 532454 605174
rect 531834 569494 532454 604938
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 529384 439174 529704 439206
rect 529384 438938 529426 439174
rect 529662 438938 529704 439174
rect 529384 438854 529704 438938
rect 529384 438618 529426 438854
rect 529662 438618 529704 438854
rect 529384 438586 529704 438618
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 259417 528734 277218
rect 531834 425494 532454 460938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 460836 542414 470898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 457897 546134 474618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 537825 439174 538145 439206
rect 537825 438938 537867 439174
rect 538103 438938 538145 439174
rect 537825 438854 538145 438938
rect 537825 438618 537867 438854
rect 538103 438618 538145 438854
rect 537825 438586 538145 438618
rect 545514 439174 546134 446095
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 533605 435454 533925 435486
rect 533605 435218 533647 435454
rect 533883 435218 533925 435454
rect 533605 435134 533925 435218
rect 533605 434898 533647 435134
rect 533883 434898 533925 435134
rect 533605 434866 533925 434898
rect 542046 435454 542366 435486
rect 542046 435218 542088 435454
rect 542324 435218 542366 435454
rect 542046 435134 542366 435218
rect 542046 434898 542088 435134
rect 542324 434898 542366 435134
rect 542046 434866 542366 434898
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 541794 399454 542414 425068
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 538811 319428 538877 319429
rect 538811 319364 538812 319428
rect 538876 319364 538877 319428
rect 538811 319363 538877 319364
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 479568 259174 479888 259206
rect 479568 258938 479610 259174
rect 479846 258938 479888 259174
rect 479568 258854 479888 258938
rect 479568 258618 479610 258854
rect 479846 258618 479888 258854
rect 479568 258586 479888 258618
rect 510288 259174 510608 259206
rect 510288 258938 510330 259174
rect 510566 258938 510608 259174
rect 510288 258854 510608 258938
rect 510288 258618 510330 258854
rect 510566 258618 510608 258854
rect 510288 258586 510608 258618
rect 464208 255454 464528 255486
rect 464208 255218 464250 255454
rect 464486 255218 464528 255454
rect 464208 255134 464528 255218
rect 464208 254898 464250 255134
rect 464486 254898 464528 255134
rect 464208 254866 464528 254898
rect 494928 255454 495248 255486
rect 494928 255218 494970 255454
rect 495206 255218 495248 255454
rect 494928 255134 495248 255218
rect 494928 254898 494970 255134
rect 495206 254898 495248 255134
rect 494928 254866 495248 254898
rect 525648 255454 525968 255486
rect 525648 255218 525690 255454
rect 525926 255218 525968 255454
rect 525648 255134 525968 255218
rect 525648 254898 525690 255134
rect 525926 254898 525968 255134
rect 525648 254866 525968 254898
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 459834 209494 460454 244938
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 479568 223174 479888 223206
rect 479568 222938 479610 223174
rect 479846 222938 479888 223174
rect 479568 222854 479888 222938
rect 479568 222618 479610 222854
rect 479846 222618 479888 222854
rect 479568 222586 479888 222618
rect 510288 223174 510608 223206
rect 510288 222938 510330 223174
rect 510566 222938 510608 223174
rect 510288 222854 510608 222938
rect 510288 222618 510330 222854
rect 510566 222618 510608 222854
rect 510288 222586 510608 222618
rect 464208 219454 464528 219486
rect 464208 219218 464250 219454
rect 464486 219218 464528 219454
rect 464208 219134 464528 219218
rect 464208 218898 464250 219134
rect 464486 218898 464528 219134
rect 464208 218866 464528 218898
rect 494928 219454 495248 219486
rect 494928 219218 494970 219454
rect 495206 219218 495248 219454
rect 494928 219134 495248 219218
rect 494928 218898 494970 219134
rect 495206 218898 495248 219134
rect 494928 218866 495248 218898
rect 525648 219454 525968 219486
rect 525648 219218 525690 219454
rect 525926 219218 525968 219454
rect 525648 219134 525968 219218
rect 525648 218898 525690 219134
rect 525926 218898 525968 219134
rect 525648 218866 525968 218898
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 458955 39268 459021 39269
rect 458955 39204 458956 39268
rect 459020 39204 459021 39268
rect 458955 39203 459021 39204
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 183454 470414 201919
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 187174 474134 201919
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 190894 477854 201919
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 194614 481574 201919
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 484674 198334 485294 201919
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 488394 166054 489014 201919
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 139281 489014 165498
rect 505794 183454 506414 201919
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 139281 506414 146898
rect 509514 187174 510134 201919
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 139281 510134 150618
rect 513234 190894 513854 201919
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 139281 513854 154338
rect 516954 194614 517574 201919
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 139281 517574 158058
rect 520674 198334 521294 201919
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 139281 521294 161778
rect 524394 166054 525014 201919
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 139281 525014 165498
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 139281 532454 172938
rect 538814 137869 538874 319363
rect 541794 291454 542414 326898
rect 545514 403174 546134 438618
rect 546266 439174 546586 439206
rect 546266 438938 546308 439174
rect 546544 438938 546586 439174
rect 546266 438854 546586 438938
rect 546266 438618 546308 438854
rect 546544 438618 546586 438854
rect 546266 438586 546586 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 542675 315348 542741 315349
rect 542675 315284 542676 315348
rect 542740 315284 542741 315348
rect 542675 315283 542741 315284
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 538811 137868 538877 137869
rect 538811 137804 538812 137868
rect 538876 137804 538877 137868
rect 538811 137803 538877 137804
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484208 111454 484528 111486
rect 484208 111218 484250 111454
rect 484486 111218 484528 111454
rect 484208 111134 484528 111218
rect 484208 110898 484250 111134
rect 484486 110898 484528 111134
rect 484208 110866 484528 110898
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 90334 485294 125778
rect 499568 115174 499888 115206
rect 499568 114938 499610 115174
rect 499846 114938 499888 115174
rect 499568 114854 499888 114938
rect 499568 114618 499610 114854
rect 499846 114618 499888 114854
rect 499568 114586 499888 114618
rect 530288 115174 530608 115206
rect 530288 114938 530330 115174
rect 530566 114938 530608 115174
rect 530288 114854 530608 114938
rect 530288 114618 530330 114854
rect 530566 114618 530608 114854
rect 530288 114586 530608 114618
rect 514928 111454 515248 111486
rect 514928 111218 514970 111454
rect 515206 111218 515248 111454
rect 514928 111134 515248 111218
rect 514928 110898 514970 111134
rect 515206 110898 515248 111134
rect 514928 110866 515248 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 58054 489014 82599
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 61774 492734 82599
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 65494 496454 82599
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 82599
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 79174 510134 82599
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 46894 513854 82599
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 50614 517574 82599
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 54334 521294 82599
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 58054 525014 82599
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 61774 528734 82599
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 65494 532454 82599
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 75454 542414 110898
rect 542678 84421 542738 315283
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 542675 84420 542741 84421
rect 542675 84356 542676 84420
rect 542740 84356 542741 84420
rect 542675 84355 542741 84356
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 51692 546134 78618
rect 549234 406894 549854 442338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556291 699820 556357 699821
rect 556291 699756 556292 699820
rect 556356 699756 556357 699820
rect 556291 699755 556357 699756
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 550487 435454 550807 435486
rect 550487 435218 550529 435454
rect 550765 435218 550807 435454
rect 550487 435134 550807 435218
rect 550487 434898 550529 435134
rect 550765 434898 550807 435134
rect 550487 434866 550807 434898
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 552954 410614 553574 446058
rect 554707 439174 555027 439206
rect 554707 438938 554749 439174
rect 554985 438938 555027 439174
rect 554707 438854 555027 438938
rect 554707 438618 554749 438854
rect 554985 438618 555027 438854
rect 554707 438586 555027 438618
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 377884 553574 410058
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 554876 367174 555196 367206
rect 554876 366938 554918 367174
rect 555154 366938 555196 367174
rect 554876 366854 555196 366938
rect 554876 366618 554918 366854
rect 555154 366618 555196 366854
rect 554876 366586 555196 366618
rect 552910 363454 553230 363486
rect 552910 363218 552952 363454
rect 553188 363218 553230 363454
rect 552910 363134 553230 363218
rect 552910 362898 552952 363134
rect 553188 362898 553230 363134
rect 552910 362866 553230 362898
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 552954 338614 553574 360068
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 556294 321469 556354 699755
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378243 557294 413778
rect 556674 378007 556706 378243
rect 556942 378007 557026 378243
rect 557262 378007 557294 378243
rect 556674 377884 557294 378007
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 377884 561014 381498
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 377884 564734 385218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 558809 367174 559129 367206
rect 558809 366938 558851 367174
rect 559087 366938 559129 367174
rect 558809 366854 559129 366938
rect 558809 366618 558851 366854
rect 559087 366618 559129 366854
rect 558809 366586 559129 366618
rect 562742 367174 563062 367206
rect 562742 366938 562784 367174
rect 563020 366938 563062 367174
rect 562742 366854 563062 366938
rect 562742 366618 562784 366854
rect 563020 366618 563062 366854
rect 562742 366586 563062 366618
rect 566675 367174 566995 367206
rect 566675 366938 566717 367174
rect 566953 366938 566995 367174
rect 566675 366854 566995 366938
rect 566675 366618 566717 366854
rect 566953 366618 566995 366854
rect 566675 366586 566995 366618
rect 556843 363454 557163 363486
rect 556843 363218 556885 363454
rect 557121 363218 557163 363454
rect 556843 363134 557163 363218
rect 556843 362898 556885 363134
rect 557121 362898 557163 363134
rect 556843 362866 557163 362898
rect 560776 363454 561096 363486
rect 560776 363218 560818 363454
rect 561054 363218 561096 363454
rect 560776 363134 561096 363218
rect 560776 362898 560818 363134
rect 561054 362898 561096 363134
rect 560776 362866 561096 362898
rect 564709 363454 565029 363486
rect 564709 363218 564751 363454
rect 564987 363218 565029 363454
rect 564709 363134 565029 363218
rect 564709 362898 564751 363134
rect 564987 362898 565029 363134
rect 564709 362866 565029 362898
rect 556674 342334 557294 360068
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556291 321468 556357 321469
rect 556291 321404 556292 321468
rect 556356 321404 556357 321468
rect 556291 321403 556357 321404
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 51692 553574 86058
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 545888 43174 546208 43206
rect 545888 42938 545930 43174
rect 546166 42938 546208 43174
rect 545888 42854 546208 42938
rect 545888 42618 545930 42854
rect 546166 42618 546208 42854
rect 545888 42586 546208 42618
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 543416 39454 543736 39486
rect 543416 39218 543458 39454
rect 543694 39218 543736 39454
rect 543416 39134 543736 39218
rect 543416 38898 543458 39134
rect 543694 38898 543736 39134
rect 543416 38866 543736 38898
rect 548361 39454 548681 39486
rect 548361 39218 548403 39454
rect 548639 39218 548681 39454
rect 548361 39134 548681 39218
rect 548361 38898 548403 39134
rect 548639 38898 548681 39134
rect 548361 38866 548681 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 30068
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 46338
rect 550833 43174 551153 43206
rect 550833 42938 550875 43174
rect 551111 42938 551153 43174
rect 550833 42854 551153 42938
rect 550833 42618 550875 42854
rect 551111 42618 551153 42854
rect 550833 42586 551153 42618
rect 555778 43174 556098 43206
rect 555778 42938 555820 43174
rect 556056 42938 556098 43174
rect 555778 42854 556098 42938
rect 555778 42618 555820 42854
rect 556056 42618 556098 42854
rect 555778 42586 556098 42618
rect 553306 39454 553626 39486
rect 553306 39218 553348 39454
rect 553584 39218 553626 39454
rect 553306 39134 553626 39218
rect 553306 38898 553348 39134
rect 553584 38898 553626 39134
rect 553306 38866 553626 38898
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 30068
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 18334 557294 53778
rect 560394 346054 561014 360068
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 51692 561014 57498
rect 564114 349774 564734 360068
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 560723 43174 561043 43206
rect 560723 42938 560765 43174
rect 561001 42938 561043 43174
rect 560723 42854 561043 42938
rect 560723 42618 560765 42854
rect 561001 42618 561043 42854
rect 560723 42586 561043 42618
rect 558251 39454 558571 39486
rect 558251 39218 558293 39454
rect 558529 39218 558571 39454
rect 558251 39134 558571 39218
rect 558251 38898 558293 39134
rect 558529 38898 558571 39134
rect 558251 38866 558571 38898
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 22054 561014 30068
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 24250 651218 24486 651454
rect 24250 650898 24486 651134
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 39610 654938 39846 655174
rect 39610 654618 39846 654854
rect 70330 654938 70566 655174
rect 70330 654618 70566 654854
rect 101050 654938 101286 655174
rect 101050 654618 101286 654854
rect 131770 654938 132006 655174
rect 131770 654618 132006 654854
rect 162490 654938 162726 655174
rect 162490 654618 162726 654854
rect 193210 654938 193446 655174
rect 193210 654618 193446 654854
rect 223930 654938 224166 655174
rect 223930 654618 224166 654854
rect 254650 654938 254886 655174
rect 254650 654618 254886 654854
rect 285370 654938 285606 655174
rect 285370 654618 285606 654854
rect 316090 654938 316326 655174
rect 316090 654618 316326 654854
rect 346810 654938 347046 655174
rect 346810 654618 347046 654854
rect 54970 651218 55206 651454
rect 54970 650898 55206 651134
rect 85690 651218 85926 651454
rect 85690 650898 85926 651134
rect 116410 651218 116646 651454
rect 116410 650898 116646 651134
rect 147130 651218 147366 651454
rect 147130 650898 147366 651134
rect 177850 651218 178086 651454
rect 177850 650898 178086 651134
rect 208570 651218 208806 651454
rect 208570 650898 208806 651134
rect 239290 651218 239526 651454
rect 239290 650898 239526 651134
rect 270010 651218 270246 651454
rect 270010 650898 270246 651134
rect 300730 651218 300966 651454
rect 300730 650898 300966 651134
rect 331450 651218 331686 651454
rect 331450 650898 331686 651134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24250 615218 24486 615454
rect 24250 614898 24486 615134
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 39610 618938 39846 619174
rect 39610 618618 39846 618854
rect 70330 618938 70566 619174
rect 70330 618618 70566 618854
rect 101050 618938 101286 619174
rect 101050 618618 101286 618854
rect 131770 618938 132006 619174
rect 131770 618618 132006 618854
rect 162490 618938 162726 619174
rect 162490 618618 162726 618854
rect 193210 618938 193446 619174
rect 193210 618618 193446 618854
rect 223930 618938 224166 619174
rect 223930 618618 224166 618854
rect 254650 618938 254886 619174
rect 254650 618618 254886 618854
rect 285370 618938 285606 619174
rect 285370 618618 285606 618854
rect 316090 618938 316326 619174
rect 316090 618618 316326 618854
rect 346810 618938 347046 619174
rect 346810 618618 347046 618854
rect 54970 615218 55206 615454
rect 54970 614898 55206 615134
rect 85690 615218 85926 615454
rect 85690 614898 85926 615134
rect 116410 615218 116646 615454
rect 116410 614898 116646 615134
rect 147130 615218 147366 615454
rect 147130 614898 147366 615134
rect 177850 615218 178086 615454
rect 177850 614898 178086 615134
rect 208570 615218 208806 615454
rect 208570 614898 208806 615134
rect 239290 615218 239526 615454
rect 239290 614898 239526 615134
rect 270010 615218 270246 615454
rect 270010 614898 270246 615134
rect 300730 615218 300966 615454
rect 300730 614898 300966 615134
rect 331450 615218 331686 615454
rect 331450 614898 331686 615134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 24250 579218 24486 579454
rect 24250 578898 24486 579134
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 39610 582938 39846 583174
rect 39610 582618 39846 582854
rect 70330 582938 70566 583174
rect 70330 582618 70566 582854
rect 101050 582938 101286 583174
rect 101050 582618 101286 582854
rect 131770 582938 132006 583174
rect 131770 582618 132006 582854
rect 162490 582938 162726 583174
rect 162490 582618 162726 582854
rect 193210 582938 193446 583174
rect 193210 582618 193446 582854
rect 223930 582938 224166 583174
rect 223930 582618 224166 582854
rect 254650 582938 254886 583174
rect 254650 582618 254886 582854
rect 285370 582938 285606 583174
rect 285370 582618 285606 582854
rect 316090 582938 316326 583174
rect 316090 582618 316326 582854
rect 346810 582938 347046 583174
rect 346810 582618 347046 582854
rect 54970 579218 55206 579454
rect 54970 578898 55206 579134
rect 85690 579218 85926 579454
rect 85690 578898 85926 579134
rect 116410 579218 116646 579454
rect 116410 578898 116646 579134
rect 147130 579218 147366 579454
rect 147130 578898 147366 579134
rect 177850 579218 178086 579454
rect 177850 578898 178086 579134
rect 208570 579218 208806 579454
rect 208570 578898 208806 579134
rect 239290 579218 239526 579454
rect 239290 578898 239526 579134
rect 270010 579218 270246 579454
rect 270010 578898 270246 579134
rect 300730 579218 300966 579454
rect 300730 578898 300966 579134
rect 331450 579218 331686 579454
rect 331450 578898 331686 579134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 24250 543218 24486 543454
rect 24250 542898 24486 543134
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 39610 546938 39846 547174
rect 39610 546618 39846 546854
rect 70330 546938 70566 547174
rect 70330 546618 70566 546854
rect 101050 546938 101286 547174
rect 101050 546618 101286 546854
rect 131770 546938 132006 547174
rect 131770 546618 132006 546854
rect 162490 546938 162726 547174
rect 162490 546618 162726 546854
rect 193210 546938 193446 547174
rect 193210 546618 193446 546854
rect 223930 546938 224166 547174
rect 223930 546618 224166 546854
rect 254650 546938 254886 547174
rect 254650 546618 254886 546854
rect 285370 546938 285606 547174
rect 285370 546618 285606 546854
rect 316090 546938 316326 547174
rect 316090 546618 316326 546854
rect 346810 546938 347046 547174
rect 346810 546618 347046 546854
rect 54970 543218 55206 543454
rect 54970 542898 55206 543134
rect 85690 543218 85926 543454
rect 85690 542898 85926 543134
rect 116410 543218 116646 543454
rect 116410 542898 116646 543134
rect 147130 543218 147366 543454
rect 147130 542898 147366 543134
rect 177850 543218 178086 543454
rect 177850 542898 178086 543134
rect 208570 543218 208806 543454
rect 208570 542898 208806 543134
rect 239290 543218 239526 543454
rect 239290 542898 239526 543134
rect 270010 543218 270246 543454
rect 270010 542898 270246 543134
rect 300730 543218 300966 543454
rect 300730 542898 300966 543134
rect 331450 543218 331686 543454
rect 331450 542898 331686 543134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 24250 507218 24486 507454
rect 24250 506898 24486 507134
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 39610 510938 39846 511174
rect 39610 510618 39846 510854
rect 70330 510938 70566 511174
rect 70330 510618 70566 510854
rect 101050 510938 101286 511174
rect 101050 510618 101286 510854
rect 131770 510938 132006 511174
rect 131770 510618 132006 510854
rect 162490 510938 162726 511174
rect 162490 510618 162726 510854
rect 193210 510938 193446 511174
rect 193210 510618 193446 510854
rect 223930 510938 224166 511174
rect 223930 510618 224166 510854
rect 254650 510938 254886 511174
rect 254650 510618 254886 510854
rect 285370 510938 285606 511174
rect 285370 510618 285606 510854
rect 316090 510938 316326 511174
rect 316090 510618 316326 510854
rect 346810 510938 347046 511174
rect 346810 510618 347046 510854
rect 54970 507218 55206 507454
rect 54970 506898 55206 507134
rect 85690 507218 85926 507454
rect 85690 506898 85926 507134
rect 116410 507218 116646 507454
rect 116410 506898 116646 507134
rect 147130 507218 147366 507454
rect 147130 506898 147366 507134
rect 177850 507218 178086 507454
rect 177850 506898 178086 507134
rect 208570 507218 208806 507454
rect 208570 506898 208806 507134
rect 239290 507218 239526 507454
rect 239290 506898 239526 507134
rect 270010 507218 270246 507454
rect 270010 506898 270246 507134
rect 300730 507218 300966 507454
rect 300730 506898 300966 507134
rect 331450 507218 331686 507454
rect 331450 506898 331686 507134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 24250 471218 24486 471454
rect 24250 470898 24486 471134
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 39610 474938 39846 475174
rect 39610 474618 39846 474854
rect 70330 474938 70566 475174
rect 70330 474618 70566 474854
rect 101050 474938 101286 475174
rect 101050 474618 101286 474854
rect 131770 474938 132006 475174
rect 131770 474618 132006 474854
rect 162490 474938 162726 475174
rect 162490 474618 162726 474854
rect 193210 474938 193446 475174
rect 193210 474618 193446 474854
rect 223930 474938 224166 475174
rect 223930 474618 224166 474854
rect 254650 474938 254886 475174
rect 254650 474618 254886 474854
rect 285370 474938 285606 475174
rect 285370 474618 285606 474854
rect 316090 474938 316326 475174
rect 316090 474618 316326 474854
rect 346810 474938 347046 475174
rect 346810 474618 347046 474854
rect 54970 471218 55206 471454
rect 54970 470898 55206 471134
rect 85690 471218 85926 471454
rect 85690 470898 85926 471134
rect 116410 471218 116646 471454
rect 116410 470898 116646 471134
rect 147130 471218 147366 471454
rect 147130 470898 147366 471134
rect 177850 471218 178086 471454
rect 177850 470898 178086 471134
rect 208570 471218 208806 471454
rect 208570 470898 208806 471134
rect 239290 471218 239526 471454
rect 239290 470898 239526 471134
rect 270010 471218 270246 471454
rect 270010 470898 270246 471134
rect 300730 471218 300966 471454
rect 300730 470898 300966 471134
rect 331450 471218 331686 471454
rect 331450 470898 331686 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 24250 435218 24486 435454
rect 24250 434898 24486 435134
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 39610 438938 39846 439174
rect 39610 438618 39846 438854
rect 70330 438938 70566 439174
rect 70330 438618 70566 438854
rect 101050 438938 101286 439174
rect 101050 438618 101286 438854
rect 131770 438938 132006 439174
rect 131770 438618 132006 438854
rect 162490 438938 162726 439174
rect 162490 438618 162726 438854
rect 193210 438938 193446 439174
rect 193210 438618 193446 438854
rect 223930 438938 224166 439174
rect 223930 438618 224166 438854
rect 254650 438938 254886 439174
rect 254650 438618 254886 438854
rect 285370 438938 285606 439174
rect 285370 438618 285606 438854
rect 316090 438938 316326 439174
rect 316090 438618 316326 438854
rect 346810 438938 347046 439174
rect 346810 438618 347046 438854
rect 54970 435218 55206 435454
rect 54970 434898 55206 435134
rect 85690 435218 85926 435454
rect 85690 434898 85926 435134
rect 116410 435218 116646 435454
rect 116410 434898 116646 435134
rect 147130 435218 147366 435454
rect 147130 434898 147366 435134
rect 177850 435218 178086 435454
rect 177850 434898 178086 435134
rect 208570 435218 208806 435454
rect 208570 434898 208806 435134
rect 239290 435218 239526 435454
rect 239290 434898 239526 435134
rect 270010 435218 270246 435454
rect 270010 434898 270246 435134
rect 300730 435218 300966 435454
rect 300730 434898 300966 435134
rect 331450 435218 331686 435454
rect 331450 434898 331686 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 24250 399218 24486 399454
rect 24250 398898 24486 399134
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 39610 402938 39846 403174
rect 39610 402618 39846 402854
rect 70330 402938 70566 403174
rect 70330 402618 70566 402854
rect 101050 402938 101286 403174
rect 101050 402618 101286 402854
rect 131770 402938 132006 403174
rect 131770 402618 132006 402854
rect 162490 402938 162726 403174
rect 162490 402618 162726 402854
rect 193210 402938 193446 403174
rect 193210 402618 193446 402854
rect 223930 402938 224166 403174
rect 223930 402618 224166 402854
rect 254650 402938 254886 403174
rect 254650 402618 254886 402854
rect 285370 402938 285606 403174
rect 285370 402618 285606 402854
rect 316090 402938 316326 403174
rect 316090 402618 316326 402854
rect 346810 402938 347046 403174
rect 346810 402618 347046 402854
rect 54970 399218 55206 399454
rect 54970 398898 55206 399134
rect 85690 399218 85926 399454
rect 85690 398898 85926 399134
rect 116410 399218 116646 399454
rect 116410 398898 116646 399134
rect 147130 399218 147366 399454
rect 147130 398898 147366 399134
rect 177850 399218 178086 399454
rect 177850 398898 178086 399134
rect 208570 399218 208806 399454
rect 208570 398898 208806 399134
rect 239290 399218 239526 399454
rect 239290 398898 239526 399134
rect 270010 399218 270246 399454
rect 270010 398898 270246 399134
rect 300730 399218 300966 399454
rect 300730 398898 300966 399134
rect 331450 399218 331686 399454
rect 331450 398898 331686 399134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 24250 363218 24486 363454
rect 24250 362898 24486 363134
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 39610 366938 39846 367174
rect 39610 366618 39846 366854
rect 70330 366938 70566 367174
rect 70330 366618 70566 366854
rect 101050 366938 101286 367174
rect 101050 366618 101286 366854
rect 131770 366938 132006 367174
rect 131770 366618 132006 366854
rect 162490 366938 162726 367174
rect 162490 366618 162726 366854
rect 193210 366938 193446 367174
rect 193210 366618 193446 366854
rect 223930 366938 224166 367174
rect 223930 366618 224166 366854
rect 254650 366938 254886 367174
rect 254650 366618 254886 366854
rect 285370 366938 285606 367174
rect 285370 366618 285606 366854
rect 316090 366938 316326 367174
rect 316090 366618 316326 366854
rect 346810 366938 347046 367174
rect 346810 366618 347046 366854
rect 54970 363218 55206 363454
rect 54970 362898 55206 363134
rect 85690 363218 85926 363454
rect 85690 362898 85926 363134
rect 116410 363218 116646 363454
rect 116410 362898 116646 363134
rect 147130 363218 147366 363454
rect 147130 362898 147366 363134
rect 177850 363218 178086 363454
rect 177850 362898 178086 363134
rect 208570 363218 208806 363454
rect 208570 362898 208806 363134
rect 239290 363218 239526 363454
rect 239290 362898 239526 363134
rect 270010 363218 270246 363454
rect 270010 362898 270246 363134
rect 300730 363218 300966 363454
rect 300730 362898 300966 363134
rect 331450 363218 331686 363454
rect 331450 362898 331686 363134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 24250 327218 24486 327454
rect 24250 326898 24486 327134
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 39610 330938 39846 331174
rect 39610 330618 39846 330854
rect 70330 330938 70566 331174
rect 70330 330618 70566 330854
rect 101050 330938 101286 331174
rect 101050 330618 101286 330854
rect 131770 330938 132006 331174
rect 131770 330618 132006 330854
rect 162490 330938 162726 331174
rect 162490 330618 162726 330854
rect 193210 330938 193446 331174
rect 193210 330618 193446 330854
rect 223930 330938 224166 331174
rect 223930 330618 224166 330854
rect 254650 330938 254886 331174
rect 254650 330618 254886 330854
rect 285370 330938 285606 331174
rect 285370 330618 285606 330854
rect 316090 330938 316326 331174
rect 316090 330618 316326 330854
rect 346810 330938 347046 331174
rect 346810 330618 347046 330854
rect 54970 327218 55206 327454
rect 54970 326898 55206 327134
rect 85690 327218 85926 327454
rect 85690 326898 85926 327134
rect 116410 327218 116646 327454
rect 116410 326898 116646 327134
rect 147130 327218 147366 327454
rect 147130 326898 147366 327134
rect 177850 327218 178086 327454
rect 177850 326898 178086 327134
rect 208570 327218 208806 327454
rect 208570 326898 208806 327134
rect 239290 327218 239526 327454
rect 239290 326898 239526 327134
rect 270010 327218 270246 327454
rect 270010 326898 270246 327134
rect 300730 327218 300966 327454
rect 300730 326898 300966 327134
rect 331450 327218 331686 327454
rect 331450 326898 331686 327134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 24250 291218 24486 291454
rect 24250 290898 24486 291134
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 39610 294938 39846 295174
rect 39610 294618 39846 294854
rect 70330 294938 70566 295174
rect 70330 294618 70566 294854
rect 101050 294938 101286 295174
rect 101050 294618 101286 294854
rect 131770 294938 132006 295174
rect 131770 294618 132006 294854
rect 162490 294938 162726 295174
rect 162490 294618 162726 294854
rect 193210 294938 193446 295174
rect 193210 294618 193446 294854
rect 223930 294938 224166 295174
rect 223930 294618 224166 294854
rect 254650 294938 254886 295174
rect 254650 294618 254886 294854
rect 285370 294938 285606 295174
rect 285370 294618 285606 294854
rect 316090 294938 316326 295174
rect 316090 294618 316326 294854
rect 346810 294938 347046 295174
rect 346810 294618 347046 294854
rect 54970 291218 55206 291454
rect 54970 290898 55206 291134
rect 85690 291218 85926 291454
rect 85690 290898 85926 291134
rect 116410 291218 116646 291454
rect 116410 290898 116646 291134
rect 147130 291218 147366 291454
rect 147130 290898 147366 291134
rect 177850 291218 178086 291454
rect 177850 290898 178086 291134
rect 208570 291218 208806 291454
rect 208570 290898 208806 291134
rect 239290 291218 239526 291454
rect 239290 290898 239526 291134
rect 270010 291218 270246 291454
rect 270010 290898 270246 291134
rect 300730 291218 300966 291454
rect 300730 290898 300966 291134
rect 331450 291218 331686 291454
rect 331450 290898 331686 291134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 24250 255218 24486 255454
rect 24250 254898 24486 255134
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 39610 258938 39846 259174
rect 39610 258618 39846 258854
rect 70330 258938 70566 259174
rect 70330 258618 70566 258854
rect 101050 258938 101286 259174
rect 101050 258618 101286 258854
rect 131770 258938 132006 259174
rect 131770 258618 132006 258854
rect 162490 258938 162726 259174
rect 162490 258618 162726 258854
rect 193210 258938 193446 259174
rect 193210 258618 193446 258854
rect 223930 258938 224166 259174
rect 223930 258618 224166 258854
rect 254650 258938 254886 259174
rect 254650 258618 254886 258854
rect 285370 258938 285606 259174
rect 285370 258618 285606 258854
rect 316090 258938 316326 259174
rect 316090 258618 316326 258854
rect 346810 258938 347046 259174
rect 346810 258618 347046 258854
rect 54970 255218 55206 255454
rect 54970 254898 55206 255134
rect 85690 255218 85926 255454
rect 85690 254898 85926 255134
rect 116410 255218 116646 255454
rect 116410 254898 116646 255134
rect 147130 255218 147366 255454
rect 147130 254898 147366 255134
rect 177850 255218 178086 255454
rect 177850 254898 178086 255134
rect 208570 255218 208806 255454
rect 208570 254898 208806 255134
rect 239290 255218 239526 255454
rect 239290 254898 239526 255134
rect 270010 255218 270246 255454
rect 270010 254898 270246 255134
rect 300730 255218 300966 255454
rect 300730 254898 300966 255134
rect 331450 255218 331686 255454
rect 331450 254898 331686 255134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 24250 219218 24486 219454
rect 24250 218898 24486 219134
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 39610 222938 39846 223174
rect 39610 222618 39846 222854
rect 70330 222938 70566 223174
rect 70330 222618 70566 222854
rect 101050 222938 101286 223174
rect 101050 222618 101286 222854
rect 131770 222938 132006 223174
rect 131770 222618 132006 222854
rect 162490 222938 162726 223174
rect 162490 222618 162726 222854
rect 193210 222938 193446 223174
rect 193210 222618 193446 222854
rect 223930 222938 224166 223174
rect 223930 222618 224166 222854
rect 254650 222938 254886 223174
rect 254650 222618 254886 222854
rect 285370 222938 285606 223174
rect 285370 222618 285606 222854
rect 316090 222938 316326 223174
rect 316090 222618 316326 222854
rect 346810 222938 347046 223174
rect 346810 222618 347046 222854
rect 54970 219218 55206 219454
rect 54970 218898 55206 219134
rect 85690 219218 85926 219454
rect 85690 218898 85926 219134
rect 116410 219218 116646 219454
rect 116410 218898 116646 219134
rect 147130 219218 147366 219454
rect 147130 218898 147366 219134
rect 177850 219218 178086 219454
rect 177850 218898 178086 219134
rect 208570 219218 208806 219454
rect 208570 218898 208806 219134
rect 239290 219218 239526 219454
rect 239290 218898 239526 219134
rect 270010 219218 270246 219454
rect 270010 218898 270246 219134
rect 300730 219218 300966 219454
rect 300730 218898 300966 219134
rect 331450 219218 331686 219454
rect 331450 218898 331686 219134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24250 183218 24486 183454
rect 24250 182898 24486 183134
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 39610 186938 39846 187174
rect 39610 186618 39846 186854
rect 70330 186938 70566 187174
rect 70330 186618 70566 186854
rect 101050 186938 101286 187174
rect 101050 186618 101286 186854
rect 131770 186938 132006 187174
rect 131770 186618 132006 186854
rect 162490 186938 162726 187174
rect 162490 186618 162726 186854
rect 193210 186938 193446 187174
rect 193210 186618 193446 186854
rect 223930 186938 224166 187174
rect 223930 186618 224166 186854
rect 254650 186938 254886 187174
rect 254650 186618 254886 186854
rect 285370 186938 285606 187174
rect 285370 186618 285606 186854
rect 316090 186938 316326 187174
rect 316090 186618 316326 186854
rect 346810 186938 347046 187174
rect 346810 186618 347046 186854
rect 54970 183218 55206 183454
rect 54970 182898 55206 183134
rect 85690 183218 85926 183454
rect 85690 182898 85926 183134
rect 116410 183218 116646 183454
rect 116410 182898 116646 183134
rect 147130 183218 147366 183454
rect 147130 182898 147366 183134
rect 177850 183218 178086 183454
rect 177850 182898 178086 183134
rect 208570 183218 208806 183454
rect 208570 182898 208806 183134
rect 239290 183218 239526 183454
rect 239290 182898 239526 183134
rect 270010 183218 270246 183454
rect 270010 182898 270246 183134
rect 300730 183218 300966 183454
rect 300730 182898 300966 183134
rect 331450 183218 331686 183454
rect 331450 182898 331686 183134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 24250 147218 24486 147454
rect 24250 146898 24486 147134
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 39610 150938 39846 151174
rect 39610 150618 39846 150854
rect 70330 150938 70566 151174
rect 70330 150618 70566 150854
rect 101050 150938 101286 151174
rect 101050 150618 101286 150854
rect 131770 150938 132006 151174
rect 131770 150618 132006 150854
rect 162490 150938 162726 151174
rect 162490 150618 162726 150854
rect 193210 150938 193446 151174
rect 193210 150618 193446 150854
rect 223930 150938 224166 151174
rect 223930 150618 224166 150854
rect 254650 150938 254886 151174
rect 254650 150618 254886 150854
rect 285370 150938 285606 151174
rect 285370 150618 285606 150854
rect 316090 150938 316326 151174
rect 316090 150618 316326 150854
rect 346810 150938 347046 151174
rect 346810 150618 347046 150854
rect 54970 147218 55206 147454
rect 54970 146898 55206 147134
rect 85690 147218 85926 147454
rect 85690 146898 85926 147134
rect 116410 147218 116646 147454
rect 116410 146898 116646 147134
rect 147130 147218 147366 147454
rect 147130 146898 147366 147134
rect 177850 147218 178086 147454
rect 177850 146898 178086 147134
rect 208570 147218 208806 147454
rect 208570 146898 208806 147134
rect 239290 147218 239526 147454
rect 239290 146898 239526 147134
rect 270010 147218 270246 147454
rect 270010 146898 270246 147134
rect 300730 147218 300966 147454
rect 300730 146898 300966 147134
rect 331450 147218 331686 147454
rect 331450 146898 331686 147134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 24250 111218 24486 111454
rect 24250 110898 24486 111134
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 39610 114938 39846 115174
rect 39610 114618 39846 114854
rect 70330 114938 70566 115174
rect 70330 114618 70566 114854
rect 101050 114938 101286 115174
rect 101050 114618 101286 114854
rect 131770 114938 132006 115174
rect 131770 114618 132006 114854
rect 162490 114938 162726 115174
rect 162490 114618 162726 114854
rect 193210 114938 193446 115174
rect 193210 114618 193446 114854
rect 223930 114938 224166 115174
rect 223930 114618 224166 114854
rect 254650 114938 254886 115174
rect 254650 114618 254886 114854
rect 285370 114938 285606 115174
rect 285370 114618 285606 114854
rect 316090 114938 316326 115174
rect 316090 114618 316326 114854
rect 346810 114938 347046 115174
rect 346810 114618 347046 114854
rect 54970 111218 55206 111454
rect 54970 110898 55206 111134
rect 85690 111218 85926 111454
rect 85690 110898 85926 111134
rect 116410 111218 116646 111454
rect 116410 110898 116646 111134
rect 147130 111218 147366 111454
rect 147130 110898 147366 111134
rect 177850 111218 178086 111454
rect 177850 110898 178086 111134
rect 208570 111218 208806 111454
rect 208570 110898 208806 111134
rect 239290 111218 239526 111454
rect 239290 110898 239526 111134
rect 270010 111218 270246 111454
rect 270010 110898 270246 111134
rect 300730 111218 300966 111454
rect 300730 110898 300966 111134
rect 331450 111218 331686 111454
rect 331450 110898 331686 111134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 24250 75218 24486 75454
rect 24250 74898 24486 75134
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 39610 78938 39846 79174
rect 39610 78618 39846 78854
rect 70330 78938 70566 79174
rect 70330 78618 70566 78854
rect 101050 78938 101286 79174
rect 101050 78618 101286 78854
rect 131770 78938 132006 79174
rect 131770 78618 132006 78854
rect 162490 78938 162726 79174
rect 162490 78618 162726 78854
rect 193210 78938 193446 79174
rect 193210 78618 193446 78854
rect 223930 78938 224166 79174
rect 223930 78618 224166 78854
rect 254650 78938 254886 79174
rect 254650 78618 254886 78854
rect 285370 78938 285606 79174
rect 285370 78618 285606 78854
rect 316090 78938 316326 79174
rect 316090 78618 316326 78854
rect 346810 78938 347046 79174
rect 346810 78618 347046 78854
rect 54970 75218 55206 75454
rect 54970 74898 55206 75134
rect 85690 75218 85926 75454
rect 85690 74898 85926 75134
rect 116410 75218 116646 75454
rect 116410 74898 116646 75134
rect 147130 75218 147366 75454
rect 147130 74898 147366 75134
rect 177850 75218 178086 75454
rect 177850 74898 178086 75134
rect 208570 75218 208806 75454
rect 208570 74898 208806 75134
rect 239290 75218 239526 75454
rect 239290 74898 239526 75134
rect 270010 75218 270246 75454
rect 270010 74898 270246 75134
rect 300730 75218 300966 75454
rect 300730 74898 300966 75134
rect 331450 75218 331686 75454
rect 331450 74898 331686 75134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 404459 327218 404695 327454
rect 404459 326898 404695 327134
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 407932 330938 408168 331174
rect 407932 330618 408168 330854
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 411405 327218 411641 327454
rect 411405 326898 411641 327134
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 414878 330938 415114 331174
rect 414878 330618 415114 330854
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 426666 438938 426902 439174
rect 426666 438618 426902 438854
rect 432347 438938 432583 439174
rect 432347 438618 432583 438854
rect 438028 438938 438264 439174
rect 438028 438618 438264 438854
rect 443709 438938 443945 439174
rect 443709 438618 443945 438854
rect 423826 435218 424062 435454
rect 423826 434898 424062 435134
rect 429507 435218 429743 435454
rect 429507 434898 429743 435134
rect 435188 435218 435424 435454
rect 435188 434898 435424 435134
rect 440869 435218 441105 435454
rect 440869 434898 441105 435134
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 418351 327218 418587 327454
rect 418351 326898 418587 327134
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 421824 330938 422060 331174
rect 421824 330618 422060 330854
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 425297 327218 425533 327454
rect 425297 326898 425533 327134
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 428770 330938 429006 331174
rect 428770 330618 429006 330854
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 452205 507218 452441 507454
rect 452205 506898 452441 507134
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 453424 510938 453660 511174
rect 453424 510618 453660 510854
rect 454643 507218 454879 507454
rect 454643 506898 454879 507134
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 479610 654938 479846 655174
rect 479610 654618 479846 654854
rect 510330 654938 510566 655174
rect 510330 654618 510566 654854
rect 464250 651218 464486 651454
rect 464250 650898 464486 651134
rect 494970 651218 495206 651454
rect 494970 650898 495206 651134
rect 455862 510938 456098 511174
rect 455862 510618 456098 510854
rect 458300 510938 458536 511174
rect 458300 510618 458536 510854
rect 457081 507218 457317 507454
rect 457081 506898 457317 507134
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 525690 651218 525926 651454
rect 525690 650898 525926 651134
rect 524426 633818 524662 634054
rect 524746 633818 524982 634054
rect 524426 633498 524662 633734
rect 524746 633498 524982 633734
rect 479610 618938 479846 619174
rect 479610 618618 479846 618854
rect 510330 618938 510566 619174
rect 510330 618618 510566 618854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 460738 510938 460974 511174
rect 460738 510618 460974 510854
rect 459519 507218 459755 507454
rect 459519 506898 459755 507134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 454250 363218 454486 363454
rect 454250 362898 454486 363134
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 429610 150938 429846 151174
rect 429610 150618 429846 150854
rect 414250 147218 414486 147454
rect 414250 146898 414486 147134
rect 444970 147218 445206 147454
rect 444970 146898 445206 147134
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 454250 327218 454486 327454
rect 454250 326898 454486 327134
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473458 435218 473694 435454
rect 473458 434898 473694 435134
rect 475930 438938 476166 439174
rect 475930 438618 476166 438854
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 478403 435218 478639 435454
rect 478403 434898 478639 435134
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 483424 510938 483660 511174
rect 483424 510618 483660 510854
rect 485862 510938 486098 511174
rect 485862 510618 486098 510854
rect 488300 510938 488536 511174
rect 488300 510618 488536 510854
rect 490738 510938 490974 511174
rect 490738 510618 490974 510854
rect 482205 507218 482441 507454
rect 482205 506898 482441 507134
rect 484643 507218 484879 507454
rect 484643 506898 484879 507134
rect 487081 507218 487317 507454
rect 487081 506898 487317 507134
rect 489519 507218 489755 507454
rect 489519 506898 489755 507134
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480875 438938 481111 439174
rect 480875 438618 481111 438854
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 483348 435218 483584 435454
rect 483348 434898 483584 435134
rect 485820 438938 486056 439174
rect 485820 438618 486056 438854
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453771 488662 454007
rect 488746 453771 488982 454007
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 490765 438938 491001 439174
rect 490765 438618 491001 438854
rect 488293 435218 488529 435454
rect 488293 434898 488529 435134
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 469610 366938 469846 367174
rect 469610 366618 469846 366854
rect 484970 363218 485206 363454
rect 484970 362898 485206 363134
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 500330 366938 500566 367174
rect 500330 366618 500566 366854
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 469610 330938 469846 331174
rect 469610 330618 469846 330854
rect 484970 327218 485206 327454
rect 484970 326898 485206 327134
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 500330 330938 500566 331174
rect 500330 330618 500566 330854
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 525690 615218 525926 615454
rect 525690 614898 525926 615134
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 528146 637538 528382 637774
rect 528466 637538 528702 637774
rect 528146 637218 528382 637454
rect 528466 637218 528702 637454
rect 528146 601538 528382 601774
rect 528466 601538 528702 601774
rect 528146 601218 528382 601454
rect 528466 601218 528702 601454
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 525206 435218 525442 435454
rect 525206 434898 525442 435134
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 531866 641258 532102 641494
rect 532186 641258 532422 641494
rect 531866 640938 532102 641174
rect 532186 640938 532422 641174
rect 531866 605258 532102 605494
rect 532186 605258 532422 605494
rect 531866 604938 532102 605174
rect 532186 604938 532422 605174
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 529426 438938 529662 439174
rect 529426 438618 529662 438854
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 537867 438938 538103 439174
rect 537867 438618 538103 438854
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 533647 435218 533883 435454
rect 533647 434898 533883 435134
rect 542088 435218 542324 435454
rect 542088 434898 542324 435134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 479610 258938 479846 259174
rect 479610 258618 479846 258854
rect 510330 258938 510566 259174
rect 510330 258618 510566 258854
rect 464250 255218 464486 255454
rect 464250 254898 464486 255134
rect 494970 255218 495206 255454
rect 494970 254898 495206 255134
rect 525690 255218 525926 255454
rect 525690 254898 525926 255134
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 479610 222938 479846 223174
rect 479610 222618 479846 222854
rect 510330 222938 510566 223174
rect 510330 222618 510566 222854
rect 464250 219218 464486 219454
rect 464250 218898 464486 219134
rect 494970 219218 495206 219454
rect 494970 218898 495206 219134
rect 525690 219218 525926 219454
rect 525690 218898 525926 219134
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 546308 438938 546544 439174
rect 546308 438618 546544 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484250 111218 484486 111454
rect 484250 110898 484486 111134
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 499610 114938 499846 115174
rect 499610 114618 499846 114854
rect 530330 114938 530566 115174
rect 530330 114618 530566 114854
rect 514970 111218 515206 111454
rect 514970 110898 515206 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 550529 435218 550765 435454
rect 550529 434898 550765 435134
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 554749 438938 554985 439174
rect 554749 438618 554985 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 554918 366938 555154 367174
rect 554918 366618 555154 366854
rect 552952 363218 553188 363454
rect 552952 362898 553188 363134
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378007 556942 378243
rect 557026 378007 557262 378243
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 558851 366938 559087 367174
rect 558851 366618 559087 366854
rect 562784 366938 563020 367174
rect 562784 366618 563020 366854
rect 566717 366938 566953 367174
rect 566717 366618 566953 366854
rect 556885 363218 557121 363454
rect 556885 362898 557121 363134
rect 560818 363218 561054 363454
rect 560818 362898 561054 363134
rect 564751 363218 564987 363454
rect 564751 362898 564987 363134
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 545930 42938 546166 43174
rect 545930 42618 546166 42854
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 543458 39218 543694 39454
rect 543458 38898 543694 39134
rect 548403 39218 548639 39454
rect 548403 38898 548639 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 550875 42938 551111 43174
rect 550875 42618 551111 42854
rect 555820 42938 556056 43174
rect 555820 42618 556056 42854
rect 553348 39218 553584 39454
rect 553348 38898 553584 39134
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 560765 42938 561001 43174
rect 560765 42618 561001 42854
rect 558293 39218 558529 39454
rect 558293 38898 558529 39134
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 39610 655174
rect 39846 654938 70330 655174
rect 70566 654938 101050 655174
rect 101286 654938 131770 655174
rect 132006 654938 162490 655174
rect 162726 654938 193210 655174
rect 193446 654938 223930 655174
rect 224166 654938 254650 655174
rect 254886 654938 285370 655174
rect 285606 654938 316090 655174
rect 316326 654938 346810 655174
rect 347046 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 479610 655174
rect 479846 654938 510330 655174
rect 510566 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 39610 654854
rect 39846 654618 70330 654854
rect 70566 654618 101050 654854
rect 101286 654618 131770 654854
rect 132006 654618 162490 654854
rect 162726 654618 193210 654854
rect 193446 654618 223930 654854
rect 224166 654618 254650 654854
rect 254886 654618 285370 654854
rect 285606 654618 316090 654854
rect 316326 654618 346810 654854
rect 347046 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 479610 654854
rect 479846 654618 510330 654854
rect 510566 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 24250 651454
rect 24486 651218 54970 651454
rect 55206 651218 85690 651454
rect 85926 651218 116410 651454
rect 116646 651218 147130 651454
rect 147366 651218 177850 651454
rect 178086 651218 208570 651454
rect 208806 651218 239290 651454
rect 239526 651218 270010 651454
rect 270246 651218 300730 651454
rect 300966 651218 331450 651454
rect 331686 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 464250 651454
rect 464486 651218 494970 651454
rect 495206 651218 525690 651454
rect 525926 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 24250 651134
rect 24486 650898 54970 651134
rect 55206 650898 85690 651134
rect 85926 650898 116410 651134
rect 116646 650898 147130 651134
rect 147366 650898 177850 651134
rect 178086 650898 208570 651134
rect 208806 650898 239290 651134
rect 239526 650898 270010 651134
rect 270246 650898 300730 651134
rect 300966 650898 331450 651134
rect 331686 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 464250 651134
rect 464486 650898 494970 651134
rect 495206 650898 525690 651134
rect 525926 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 531866 641494
rect 532102 641258 532186 641494
rect 532422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 531866 641174
rect 532102 640938 532186 641174
rect 532422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 528146 637774
rect 528382 637538 528466 637774
rect 528702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 528146 637454
rect 528382 637218 528466 637454
rect 528702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 524426 634054
rect 524662 633818 524746 634054
rect 524982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 524426 633734
rect 524662 633498 524746 633734
rect 524982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 39610 619174
rect 39846 618938 70330 619174
rect 70566 618938 101050 619174
rect 101286 618938 131770 619174
rect 132006 618938 162490 619174
rect 162726 618938 193210 619174
rect 193446 618938 223930 619174
rect 224166 618938 254650 619174
rect 254886 618938 285370 619174
rect 285606 618938 316090 619174
rect 316326 618938 346810 619174
rect 347046 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 479610 619174
rect 479846 618938 510330 619174
rect 510566 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 39610 618854
rect 39846 618618 70330 618854
rect 70566 618618 101050 618854
rect 101286 618618 131770 618854
rect 132006 618618 162490 618854
rect 162726 618618 193210 618854
rect 193446 618618 223930 618854
rect 224166 618618 254650 618854
rect 254886 618618 285370 618854
rect 285606 618618 316090 618854
rect 316326 618618 346810 618854
rect 347046 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 479610 618854
rect 479846 618618 510330 618854
rect 510566 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 24250 615454
rect 24486 615218 54970 615454
rect 55206 615218 85690 615454
rect 85926 615218 116410 615454
rect 116646 615218 147130 615454
rect 147366 615218 177850 615454
rect 178086 615218 208570 615454
rect 208806 615218 239290 615454
rect 239526 615218 270010 615454
rect 270246 615218 300730 615454
rect 300966 615218 331450 615454
rect 331686 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 525690 615454
rect 525926 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 24250 615134
rect 24486 614898 54970 615134
rect 55206 614898 85690 615134
rect 85926 614898 116410 615134
rect 116646 614898 147130 615134
rect 147366 614898 177850 615134
rect 178086 614898 208570 615134
rect 208806 614898 239290 615134
rect 239526 614898 270010 615134
rect 270246 614898 300730 615134
rect 300966 614898 331450 615134
rect 331686 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 525690 615134
rect 525926 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 531866 605494
rect 532102 605258 532186 605494
rect 532422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 531866 605174
rect 532102 604938 532186 605174
rect 532422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 528146 601774
rect 528382 601538 528466 601774
rect 528702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 528146 601454
rect 528382 601218 528466 601454
rect 528702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 39610 583174
rect 39846 582938 70330 583174
rect 70566 582938 101050 583174
rect 101286 582938 131770 583174
rect 132006 582938 162490 583174
rect 162726 582938 193210 583174
rect 193446 582938 223930 583174
rect 224166 582938 254650 583174
rect 254886 582938 285370 583174
rect 285606 582938 316090 583174
rect 316326 582938 346810 583174
rect 347046 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 39610 582854
rect 39846 582618 70330 582854
rect 70566 582618 101050 582854
rect 101286 582618 131770 582854
rect 132006 582618 162490 582854
rect 162726 582618 193210 582854
rect 193446 582618 223930 582854
rect 224166 582618 254650 582854
rect 254886 582618 285370 582854
rect 285606 582618 316090 582854
rect 316326 582618 346810 582854
rect 347046 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 24250 579454
rect 24486 579218 54970 579454
rect 55206 579218 85690 579454
rect 85926 579218 116410 579454
rect 116646 579218 147130 579454
rect 147366 579218 177850 579454
rect 178086 579218 208570 579454
rect 208806 579218 239290 579454
rect 239526 579218 270010 579454
rect 270246 579218 300730 579454
rect 300966 579218 331450 579454
rect 331686 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 24250 579134
rect 24486 578898 54970 579134
rect 55206 578898 85690 579134
rect 85926 578898 116410 579134
rect 116646 578898 147130 579134
rect 147366 578898 177850 579134
rect 178086 578898 208570 579134
rect 208806 578898 239290 579134
rect 239526 578898 270010 579134
rect 270246 578898 300730 579134
rect 300966 578898 331450 579134
rect 331686 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 39610 547174
rect 39846 546938 70330 547174
rect 70566 546938 101050 547174
rect 101286 546938 131770 547174
rect 132006 546938 162490 547174
rect 162726 546938 193210 547174
rect 193446 546938 223930 547174
rect 224166 546938 254650 547174
rect 254886 546938 285370 547174
rect 285606 546938 316090 547174
rect 316326 546938 346810 547174
rect 347046 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 39610 546854
rect 39846 546618 70330 546854
rect 70566 546618 101050 546854
rect 101286 546618 131770 546854
rect 132006 546618 162490 546854
rect 162726 546618 193210 546854
rect 193446 546618 223930 546854
rect 224166 546618 254650 546854
rect 254886 546618 285370 546854
rect 285606 546618 316090 546854
rect 316326 546618 346810 546854
rect 347046 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 24250 543454
rect 24486 543218 54970 543454
rect 55206 543218 85690 543454
rect 85926 543218 116410 543454
rect 116646 543218 147130 543454
rect 147366 543218 177850 543454
rect 178086 543218 208570 543454
rect 208806 543218 239290 543454
rect 239526 543218 270010 543454
rect 270246 543218 300730 543454
rect 300966 543218 331450 543454
rect 331686 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 24250 543134
rect 24486 542898 54970 543134
rect 55206 542898 85690 543134
rect 85926 542898 116410 543134
rect 116646 542898 147130 543134
rect 147366 542898 177850 543134
rect 178086 542898 208570 543134
rect 208806 542898 239290 543134
rect 239526 542898 270010 543134
rect 270246 542898 300730 543134
rect 300966 542898 331450 543134
rect 331686 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 39610 511174
rect 39846 510938 70330 511174
rect 70566 510938 101050 511174
rect 101286 510938 131770 511174
rect 132006 510938 162490 511174
rect 162726 510938 193210 511174
rect 193446 510938 223930 511174
rect 224166 510938 254650 511174
rect 254886 510938 285370 511174
rect 285606 510938 316090 511174
rect 316326 510938 346810 511174
rect 347046 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 453424 511174
rect 453660 510938 455862 511174
rect 456098 510938 458300 511174
rect 458536 510938 460738 511174
rect 460974 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 483424 511174
rect 483660 510938 485862 511174
rect 486098 510938 488300 511174
rect 488536 510938 490738 511174
rect 490974 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 39610 510854
rect 39846 510618 70330 510854
rect 70566 510618 101050 510854
rect 101286 510618 131770 510854
rect 132006 510618 162490 510854
rect 162726 510618 193210 510854
rect 193446 510618 223930 510854
rect 224166 510618 254650 510854
rect 254886 510618 285370 510854
rect 285606 510618 316090 510854
rect 316326 510618 346810 510854
rect 347046 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 453424 510854
rect 453660 510618 455862 510854
rect 456098 510618 458300 510854
rect 458536 510618 460738 510854
rect 460974 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 483424 510854
rect 483660 510618 485862 510854
rect 486098 510618 488300 510854
rect 488536 510618 490738 510854
rect 490974 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 24250 507454
rect 24486 507218 54970 507454
rect 55206 507218 85690 507454
rect 85926 507218 116410 507454
rect 116646 507218 147130 507454
rect 147366 507218 177850 507454
rect 178086 507218 208570 507454
rect 208806 507218 239290 507454
rect 239526 507218 270010 507454
rect 270246 507218 300730 507454
rect 300966 507218 331450 507454
rect 331686 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 452205 507454
rect 452441 507218 454643 507454
rect 454879 507218 457081 507454
rect 457317 507218 459519 507454
rect 459755 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 482205 507454
rect 482441 507218 484643 507454
rect 484879 507218 487081 507454
rect 487317 507218 489519 507454
rect 489755 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 24250 507134
rect 24486 506898 54970 507134
rect 55206 506898 85690 507134
rect 85926 506898 116410 507134
rect 116646 506898 147130 507134
rect 147366 506898 177850 507134
rect 178086 506898 208570 507134
rect 208806 506898 239290 507134
rect 239526 506898 270010 507134
rect 270246 506898 300730 507134
rect 300966 506898 331450 507134
rect 331686 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 452205 507134
rect 452441 506898 454643 507134
rect 454879 506898 457081 507134
rect 457317 506898 459519 507134
rect 459755 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 482205 507134
rect 482441 506898 484643 507134
rect 484879 506898 487081 507134
rect 487317 506898 489519 507134
rect 489755 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 39610 475174
rect 39846 474938 70330 475174
rect 70566 474938 101050 475174
rect 101286 474938 131770 475174
rect 132006 474938 162490 475174
rect 162726 474938 193210 475174
rect 193446 474938 223930 475174
rect 224166 474938 254650 475174
rect 254886 474938 285370 475174
rect 285606 474938 316090 475174
rect 316326 474938 346810 475174
rect 347046 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 39610 474854
rect 39846 474618 70330 474854
rect 70566 474618 101050 474854
rect 101286 474618 131770 474854
rect 132006 474618 162490 474854
rect 162726 474618 193210 474854
rect 193446 474618 223930 474854
rect 224166 474618 254650 474854
rect 254886 474618 285370 474854
rect 285606 474618 316090 474854
rect 316326 474618 346810 474854
rect 347046 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 24250 471454
rect 24486 471218 54970 471454
rect 55206 471218 85690 471454
rect 85926 471218 116410 471454
rect 116646 471218 147130 471454
rect 147366 471218 177850 471454
rect 178086 471218 208570 471454
rect 208806 471218 239290 471454
rect 239526 471218 270010 471454
rect 270246 471218 300730 471454
rect 300966 471218 331450 471454
rect 331686 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 24250 471134
rect 24486 470898 54970 471134
rect 55206 470898 85690 471134
rect 85926 470898 116410 471134
rect 116646 470898 147130 471134
rect 147366 470898 177850 471134
rect 178086 470898 208570 471134
rect 208806 470898 239290 471134
rect 239526 470898 270010 471134
rect 270246 470898 300730 471134
rect 300966 470898 331450 471134
rect 331686 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 454007 524426 454054
rect 452982 453818 488426 454007
rect -8726 453771 488426 453818
rect 488662 453771 488746 454007
rect 488982 453818 524426 454007
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect 488982 453771 592650 453818
rect -8726 453734 592650 453771
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 39610 439174
rect 39846 438938 70330 439174
rect 70566 438938 101050 439174
rect 101286 438938 131770 439174
rect 132006 438938 162490 439174
rect 162726 438938 193210 439174
rect 193446 438938 223930 439174
rect 224166 438938 254650 439174
rect 254886 438938 285370 439174
rect 285606 438938 316090 439174
rect 316326 438938 346810 439174
rect 347046 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 426666 439174
rect 426902 438938 432347 439174
rect 432583 438938 438028 439174
rect 438264 438938 443709 439174
rect 443945 438938 475930 439174
rect 476166 438938 480875 439174
rect 481111 438938 485820 439174
rect 486056 438938 490765 439174
rect 491001 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 529426 439174
rect 529662 438938 537867 439174
rect 538103 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546308 439174
rect 546544 438938 554749 439174
rect 554985 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 39610 438854
rect 39846 438618 70330 438854
rect 70566 438618 101050 438854
rect 101286 438618 131770 438854
rect 132006 438618 162490 438854
rect 162726 438618 193210 438854
rect 193446 438618 223930 438854
rect 224166 438618 254650 438854
rect 254886 438618 285370 438854
rect 285606 438618 316090 438854
rect 316326 438618 346810 438854
rect 347046 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 426666 438854
rect 426902 438618 432347 438854
rect 432583 438618 438028 438854
rect 438264 438618 443709 438854
rect 443945 438618 475930 438854
rect 476166 438618 480875 438854
rect 481111 438618 485820 438854
rect 486056 438618 490765 438854
rect 491001 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 529426 438854
rect 529662 438618 537867 438854
rect 538103 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546308 438854
rect 546544 438618 554749 438854
rect 554985 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 24250 435454
rect 24486 435218 54970 435454
rect 55206 435218 85690 435454
rect 85926 435218 116410 435454
rect 116646 435218 147130 435454
rect 147366 435218 177850 435454
rect 178086 435218 208570 435454
rect 208806 435218 239290 435454
rect 239526 435218 270010 435454
rect 270246 435218 300730 435454
rect 300966 435218 331450 435454
rect 331686 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 423826 435454
rect 424062 435218 429507 435454
rect 429743 435218 435188 435454
rect 435424 435218 440869 435454
rect 441105 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 473458 435454
rect 473694 435218 478403 435454
rect 478639 435218 483348 435454
rect 483584 435218 488293 435454
rect 488529 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 525206 435454
rect 525442 435218 533647 435454
rect 533883 435218 542088 435454
rect 542324 435218 550529 435454
rect 550765 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 24250 435134
rect 24486 434898 54970 435134
rect 55206 434898 85690 435134
rect 85926 434898 116410 435134
rect 116646 434898 147130 435134
rect 147366 434898 177850 435134
rect 178086 434898 208570 435134
rect 208806 434898 239290 435134
rect 239526 434898 270010 435134
rect 270246 434898 300730 435134
rect 300966 434898 331450 435134
rect 331686 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 423826 435134
rect 424062 434898 429507 435134
rect 429743 434898 435188 435134
rect 435424 434898 440869 435134
rect 441105 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 473458 435134
rect 473694 434898 478403 435134
rect 478639 434898 483348 435134
rect 483584 434898 488293 435134
rect 488529 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 525206 435134
rect 525442 434898 533647 435134
rect 533883 434898 542088 435134
rect 542324 434898 550529 435134
rect 550765 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 39610 403174
rect 39846 402938 70330 403174
rect 70566 402938 101050 403174
rect 101286 402938 131770 403174
rect 132006 402938 162490 403174
rect 162726 402938 193210 403174
rect 193446 402938 223930 403174
rect 224166 402938 254650 403174
rect 254886 402938 285370 403174
rect 285606 402938 316090 403174
rect 316326 402938 346810 403174
rect 347046 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 39610 402854
rect 39846 402618 70330 402854
rect 70566 402618 101050 402854
rect 101286 402618 131770 402854
rect 132006 402618 162490 402854
rect 162726 402618 193210 402854
rect 193446 402618 223930 402854
rect 224166 402618 254650 402854
rect 254886 402618 285370 402854
rect 285606 402618 316090 402854
rect 316326 402618 346810 402854
rect 347046 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 24250 399454
rect 24486 399218 54970 399454
rect 55206 399218 85690 399454
rect 85926 399218 116410 399454
rect 116646 399218 147130 399454
rect 147366 399218 177850 399454
rect 178086 399218 208570 399454
rect 208806 399218 239290 399454
rect 239526 399218 270010 399454
rect 270246 399218 300730 399454
rect 300966 399218 331450 399454
rect 331686 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 24250 399134
rect 24486 398898 54970 399134
rect 55206 398898 85690 399134
rect 85926 398898 116410 399134
rect 116646 398898 147130 399134
rect 147366 398898 177850 399134
rect 178086 398898 208570 399134
rect 208806 398898 239290 399134
rect 239526 398898 270010 399134
rect 270246 398898 300730 399134
rect 300966 398898 331450 399134
rect 331686 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378243 589182 378334
rect 521262 378098 556706 378243
rect -8726 378014 556706 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 378007 556706 378014
rect 556942 378007 557026 378243
rect 557262 378098 589182 378243
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect 557262 378014 592650 378098
rect 557262 378007 589182 378014
rect 521262 377778 589182 378007
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 39610 367174
rect 39846 366938 70330 367174
rect 70566 366938 101050 367174
rect 101286 366938 131770 367174
rect 132006 366938 162490 367174
rect 162726 366938 193210 367174
rect 193446 366938 223930 367174
rect 224166 366938 254650 367174
rect 254886 366938 285370 367174
rect 285606 366938 316090 367174
rect 316326 366938 346810 367174
rect 347046 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 469610 367174
rect 469846 366938 500330 367174
rect 500566 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 554918 367174
rect 555154 366938 558851 367174
rect 559087 366938 562784 367174
rect 563020 366938 566717 367174
rect 566953 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 39610 366854
rect 39846 366618 70330 366854
rect 70566 366618 101050 366854
rect 101286 366618 131770 366854
rect 132006 366618 162490 366854
rect 162726 366618 193210 366854
rect 193446 366618 223930 366854
rect 224166 366618 254650 366854
rect 254886 366618 285370 366854
rect 285606 366618 316090 366854
rect 316326 366618 346810 366854
rect 347046 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 469610 366854
rect 469846 366618 500330 366854
rect 500566 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 554918 366854
rect 555154 366618 558851 366854
rect 559087 366618 562784 366854
rect 563020 366618 566717 366854
rect 566953 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 24250 363454
rect 24486 363218 54970 363454
rect 55206 363218 85690 363454
rect 85926 363218 116410 363454
rect 116646 363218 147130 363454
rect 147366 363218 177850 363454
rect 178086 363218 208570 363454
rect 208806 363218 239290 363454
rect 239526 363218 270010 363454
rect 270246 363218 300730 363454
rect 300966 363218 331450 363454
rect 331686 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 454250 363454
rect 454486 363218 484970 363454
rect 485206 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 552952 363454
rect 553188 363218 556885 363454
rect 557121 363218 560818 363454
rect 561054 363218 564751 363454
rect 564987 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 24250 363134
rect 24486 362898 54970 363134
rect 55206 362898 85690 363134
rect 85926 362898 116410 363134
rect 116646 362898 147130 363134
rect 147366 362898 177850 363134
rect 178086 362898 208570 363134
rect 208806 362898 239290 363134
rect 239526 362898 270010 363134
rect 270246 362898 300730 363134
rect 300966 362898 331450 363134
rect 331686 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 454250 363134
rect 454486 362898 484970 363134
rect 485206 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 552952 363134
rect 553188 362898 556885 363134
rect 557121 362898 560818 363134
rect 561054 362898 564751 363134
rect 564987 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 39610 331174
rect 39846 330938 70330 331174
rect 70566 330938 101050 331174
rect 101286 330938 131770 331174
rect 132006 330938 162490 331174
rect 162726 330938 193210 331174
rect 193446 330938 223930 331174
rect 224166 330938 254650 331174
rect 254886 330938 285370 331174
rect 285606 330938 316090 331174
rect 316326 330938 346810 331174
rect 347046 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 407932 331174
rect 408168 330938 414878 331174
rect 415114 330938 421824 331174
rect 422060 330938 428770 331174
rect 429006 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 469610 331174
rect 469846 330938 500330 331174
rect 500566 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 39610 330854
rect 39846 330618 70330 330854
rect 70566 330618 101050 330854
rect 101286 330618 131770 330854
rect 132006 330618 162490 330854
rect 162726 330618 193210 330854
rect 193446 330618 223930 330854
rect 224166 330618 254650 330854
rect 254886 330618 285370 330854
rect 285606 330618 316090 330854
rect 316326 330618 346810 330854
rect 347046 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 407932 330854
rect 408168 330618 414878 330854
rect 415114 330618 421824 330854
rect 422060 330618 428770 330854
rect 429006 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 469610 330854
rect 469846 330618 500330 330854
rect 500566 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 24250 327454
rect 24486 327218 54970 327454
rect 55206 327218 85690 327454
rect 85926 327218 116410 327454
rect 116646 327218 147130 327454
rect 147366 327218 177850 327454
rect 178086 327218 208570 327454
rect 208806 327218 239290 327454
rect 239526 327218 270010 327454
rect 270246 327218 300730 327454
rect 300966 327218 331450 327454
rect 331686 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 404459 327454
rect 404695 327218 411405 327454
rect 411641 327218 418351 327454
rect 418587 327218 425297 327454
rect 425533 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 454250 327454
rect 454486 327218 484970 327454
rect 485206 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 24250 327134
rect 24486 326898 54970 327134
rect 55206 326898 85690 327134
rect 85926 326898 116410 327134
rect 116646 326898 147130 327134
rect 147366 326898 177850 327134
rect 178086 326898 208570 327134
rect 208806 326898 239290 327134
rect 239526 326898 270010 327134
rect 270246 326898 300730 327134
rect 300966 326898 331450 327134
rect 331686 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 404459 327134
rect 404695 326898 411405 327134
rect 411641 326898 418351 327134
rect 418587 326898 425297 327134
rect 425533 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 454250 327134
rect 454486 326898 484970 327134
rect 485206 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 39610 295174
rect 39846 294938 70330 295174
rect 70566 294938 101050 295174
rect 101286 294938 131770 295174
rect 132006 294938 162490 295174
rect 162726 294938 193210 295174
rect 193446 294938 223930 295174
rect 224166 294938 254650 295174
rect 254886 294938 285370 295174
rect 285606 294938 316090 295174
rect 316326 294938 346810 295174
rect 347046 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 39610 294854
rect 39846 294618 70330 294854
rect 70566 294618 101050 294854
rect 101286 294618 131770 294854
rect 132006 294618 162490 294854
rect 162726 294618 193210 294854
rect 193446 294618 223930 294854
rect 224166 294618 254650 294854
rect 254886 294618 285370 294854
rect 285606 294618 316090 294854
rect 316326 294618 346810 294854
rect 347046 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 24250 291454
rect 24486 291218 54970 291454
rect 55206 291218 85690 291454
rect 85926 291218 116410 291454
rect 116646 291218 147130 291454
rect 147366 291218 177850 291454
rect 178086 291218 208570 291454
rect 208806 291218 239290 291454
rect 239526 291218 270010 291454
rect 270246 291218 300730 291454
rect 300966 291218 331450 291454
rect 331686 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 24250 291134
rect 24486 290898 54970 291134
rect 55206 290898 85690 291134
rect 85926 290898 116410 291134
rect 116646 290898 147130 291134
rect 147366 290898 177850 291134
rect 178086 290898 208570 291134
rect 208806 290898 239290 291134
rect 239526 290898 270010 291134
rect 270246 290898 300730 291134
rect 300966 290898 331450 291134
rect 331686 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 39610 259174
rect 39846 258938 70330 259174
rect 70566 258938 101050 259174
rect 101286 258938 131770 259174
rect 132006 258938 162490 259174
rect 162726 258938 193210 259174
rect 193446 258938 223930 259174
rect 224166 258938 254650 259174
rect 254886 258938 285370 259174
rect 285606 258938 316090 259174
rect 316326 258938 346810 259174
rect 347046 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 479610 259174
rect 479846 258938 510330 259174
rect 510566 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 39610 258854
rect 39846 258618 70330 258854
rect 70566 258618 101050 258854
rect 101286 258618 131770 258854
rect 132006 258618 162490 258854
rect 162726 258618 193210 258854
rect 193446 258618 223930 258854
rect 224166 258618 254650 258854
rect 254886 258618 285370 258854
rect 285606 258618 316090 258854
rect 316326 258618 346810 258854
rect 347046 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 479610 258854
rect 479846 258618 510330 258854
rect 510566 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 24250 255454
rect 24486 255218 54970 255454
rect 55206 255218 85690 255454
rect 85926 255218 116410 255454
rect 116646 255218 147130 255454
rect 147366 255218 177850 255454
rect 178086 255218 208570 255454
rect 208806 255218 239290 255454
rect 239526 255218 270010 255454
rect 270246 255218 300730 255454
rect 300966 255218 331450 255454
rect 331686 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 464250 255454
rect 464486 255218 494970 255454
rect 495206 255218 525690 255454
rect 525926 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 24250 255134
rect 24486 254898 54970 255134
rect 55206 254898 85690 255134
rect 85926 254898 116410 255134
rect 116646 254898 147130 255134
rect 147366 254898 177850 255134
rect 178086 254898 208570 255134
rect 208806 254898 239290 255134
rect 239526 254898 270010 255134
rect 270246 254898 300730 255134
rect 300966 254898 331450 255134
rect 331686 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 464250 255134
rect 464486 254898 494970 255134
rect 495206 254898 525690 255134
rect 525926 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 39610 223174
rect 39846 222938 70330 223174
rect 70566 222938 101050 223174
rect 101286 222938 131770 223174
rect 132006 222938 162490 223174
rect 162726 222938 193210 223174
rect 193446 222938 223930 223174
rect 224166 222938 254650 223174
rect 254886 222938 285370 223174
rect 285606 222938 316090 223174
rect 316326 222938 346810 223174
rect 347046 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 479610 223174
rect 479846 222938 510330 223174
rect 510566 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 39610 222854
rect 39846 222618 70330 222854
rect 70566 222618 101050 222854
rect 101286 222618 131770 222854
rect 132006 222618 162490 222854
rect 162726 222618 193210 222854
rect 193446 222618 223930 222854
rect 224166 222618 254650 222854
rect 254886 222618 285370 222854
rect 285606 222618 316090 222854
rect 316326 222618 346810 222854
rect 347046 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 479610 222854
rect 479846 222618 510330 222854
rect 510566 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 24250 219454
rect 24486 219218 54970 219454
rect 55206 219218 85690 219454
rect 85926 219218 116410 219454
rect 116646 219218 147130 219454
rect 147366 219218 177850 219454
rect 178086 219218 208570 219454
rect 208806 219218 239290 219454
rect 239526 219218 270010 219454
rect 270246 219218 300730 219454
rect 300966 219218 331450 219454
rect 331686 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 464250 219454
rect 464486 219218 494970 219454
rect 495206 219218 525690 219454
rect 525926 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 24250 219134
rect 24486 218898 54970 219134
rect 55206 218898 85690 219134
rect 85926 218898 116410 219134
rect 116646 218898 147130 219134
rect 147366 218898 177850 219134
rect 178086 218898 208570 219134
rect 208806 218898 239290 219134
rect 239526 218898 270010 219134
rect 270246 218898 300730 219134
rect 300966 218898 331450 219134
rect 331686 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 464250 219134
rect 464486 218898 494970 219134
rect 495206 218898 525690 219134
rect 525926 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 39610 187174
rect 39846 186938 70330 187174
rect 70566 186938 101050 187174
rect 101286 186938 131770 187174
rect 132006 186938 162490 187174
rect 162726 186938 193210 187174
rect 193446 186938 223930 187174
rect 224166 186938 254650 187174
rect 254886 186938 285370 187174
rect 285606 186938 316090 187174
rect 316326 186938 346810 187174
rect 347046 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 39610 186854
rect 39846 186618 70330 186854
rect 70566 186618 101050 186854
rect 101286 186618 131770 186854
rect 132006 186618 162490 186854
rect 162726 186618 193210 186854
rect 193446 186618 223930 186854
rect 224166 186618 254650 186854
rect 254886 186618 285370 186854
rect 285606 186618 316090 186854
rect 316326 186618 346810 186854
rect 347046 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 24250 183454
rect 24486 183218 54970 183454
rect 55206 183218 85690 183454
rect 85926 183218 116410 183454
rect 116646 183218 147130 183454
rect 147366 183218 177850 183454
rect 178086 183218 208570 183454
rect 208806 183218 239290 183454
rect 239526 183218 270010 183454
rect 270246 183218 300730 183454
rect 300966 183218 331450 183454
rect 331686 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 24250 183134
rect 24486 182898 54970 183134
rect 55206 182898 85690 183134
rect 85926 182898 116410 183134
rect 116646 182898 147130 183134
rect 147366 182898 177850 183134
rect 178086 182898 208570 183134
rect 208806 182898 239290 183134
rect 239526 182898 270010 183134
rect 270246 182898 300730 183134
rect 300966 182898 331450 183134
rect 331686 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 39610 151174
rect 39846 150938 70330 151174
rect 70566 150938 101050 151174
rect 101286 150938 131770 151174
rect 132006 150938 162490 151174
rect 162726 150938 193210 151174
rect 193446 150938 223930 151174
rect 224166 150938 254650 151174
rect 254886 150938 285370 151174
rect 285606 150938 316090 151174
rect 316326 150938 346810 151174
rect 347046 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 429610 151174
rect 429846 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 39610 150854
rect 39846 150618 70330 150854
rect 70566 150618 101050 150854
rect 101286 150618 131770 150854
rect 132006 150618 162490 150854
rect 162726 150618 193210 150854
rect 193446 150618 223930 150854
rect 224166 150618 254650 150854
rect 254886 150618 285370 150854
rect 285606 150618 316090 150854
rect 316326 150618 346810 150854
rect 347046 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 429610 150854
rect 429846 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 24250 147454
rect 24486 147218 54970 147454
rect 55206 147218 85690 147454
rect 85926 147218 116410 147454
rect 116646 147218 147130 147454
rect 147366 147218 177850 147454
rect 178086 147218 208570 147454
rect 208806 147218 239290 147454
rect 239526 147218 270010 147454
rect 270246 147218 300730 147454
rect 300966 147218 331450 147454
rect 331686 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 414250 147454
rect 414486 147218 444970 147454
rect 445206 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 24250 147134
rect 24486 146898 54970 147134
rect 55206 146898 85690 147134
rect 85926 146898 116410 147134
rect 116646 146898 147130 147134
rect 147366 146898 177850 147134
rect 178086 146898 208570 147134
rect 208806 146898 239290 147134
rect 239526 146898 270010 147134
rect 270246 146898 300730 147134
rect 300966 146898 331450 147134
rect 331686 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 414250 147134
rect 414486 146898 444970 147134
rect 445206 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 39610 115174
rect 39846 114938 70330 115174
rect 70566 114938 101050 115174
rect 101286 114938 131770 115174
rect 132006 114938 162490 115174
rect 162726 114938 193210 115174
rect 193446 114938 223930 115174
rect 224166 114938 254650 115174
rect 254886 114938 285370 115174
rect 285606 114938 316090 115174
rect 316326 114938 346810 115174
rect 347046 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 499610 115174
rect 499846 114938 530330 115174
rect 530566 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 39610 114854
rect 39846 114618 70330 114854
rect 70566 114618 101050 114854
rect 101286 114618 131770 114854
rect 132006 114618 162490 114854
rect 162726 114618 193210 114854
rect 193446 114618 223930 114854
rect 224166 114618 254650 114854
rect 254886 114618 285370 114854
rect 285606 114618 316090 114854
rect 316326 114618 346810 114854
rect 347046 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 499610 114854
rect 499846 114618 530330 114854
rect 530566 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 24250 111454
rect 24486 111218 54970 111454
rect 55206 111218 85690 111454
rect 85926 111218 116410 111454
rect 116646 111218 147130 111454
rect 147366 111218 177850 111454
rect 178086 111218 208570 111454
rect 208806 111218 239290 111454
rect 239526 111218 270010 111454
rect 270246 111218 300730 111454
rect 300966 111218 331450 111454
rect 331686 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 484250 111454
rect 484486 111218 514970 111454
rect 515206 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 24250 111134
rect 24486 110898 54970 111134
rect 55206 110898 85690 111134
rect 85926 110898 116410 111134
rect 116646 110898 147130 111134
rect 147366 110898 177850 111134
rect 178086 110898 208570 111134
rect 208806 110898 239290 111134
rect 239526 110898 270010 111134
rect 270246 110898 300730 111134
rect 300966 110898 331450 111134
rect 331686 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 484250 111134
rect 484486 110898 514970 111134
rect 515206 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 39610 79174
rect 39846 78938 70330 79174
rect 70566 78938 101050 79174
rect 101286 78938 131770 79174
rect 132006 78938 162490 79174
rect 162726 78938 193210 79174
rect 193446 78938 223930 79174
rect 224166 78938 254650 79174
rect 254886 78938 285370 79174
rect 285606 78938 316090 79174
rect 316326 78938 346810 79174
rect 347046 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 39610 78854
rect 39846 78618 70330 78854
rect 70566 78618 101050 78854
rect 101286 78618 131770 78854
rect 132006 78618 162490 78854
rect 162726 78618 193210 78854
rect 193446 78618 223930 78854
rect 224166 78618 254650 78854
rect 254886 78618 285370 78854
rect 285606 78618 316090 78854
rect 316326 78618 346810 78854
rect 347046 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 24250 75454
rect 24486 75218 54970 75454
rect 55206 75218 85690 75454
rect 85926 75218 116410 75454
rect 116646 75218 147130 75454
rect 147366 75218 177850 75454
rect 178086 75218 208570 75454
rect 208806 75218 239290 75454
rect 239526 75218 270010 75454
rect 270246 75218 300730 75454
rect 300966 75218 331450 75454
rect 331686 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 24250 75134
rect 24486 74898 54970 75134
rect 55206 74898 85690 75134
rect 85926 74898 116410 75134
rect 116646 74898 147130 75134
rect 147366 74898 177850 75134
rect 178086 74898 208570 75134
rect 208806 74898 239290 75134
rect 239526 74898 270010 75134
rect 270246 74898 300730 75134
rect 300966 74898 331450 75134
rect 331686 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545930 43174
rect 546166 42938 550875 43174
rect 551111 42938 555820 43174
rect 556056 42938 560765 43174
rect 561001 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545930 42854
rect 546166 42618 550875 42854
rect 551111 42618 555820 42854
rect 556056 42618 560765 42854
rect 561001 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 543458 39454
rect 543694 39218 548403 39454
rect 548639 39218 553348 39454
rect 553584 39218 558293 39454
rect 558529 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 543458 39134
rect 543694 38898 548403 39134
rect 548639 38898 553348 39134
rect 553584 38898 558293 39134
rect 558529 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use posit_unit  posit_unit
timestamp 0
transform 1 0 460000 0 1 200000
box 0 2128 70000 67504
use multiplexer  proj_multiplexer
timestamp 0
transform 1 0 450000 0 1 322000
box 0 0 60000 64000
use tholin_avalonsemi_5401  tholin_avalonsemi_5401
timestamp 0
transform 1 0 520000 0 1 425000
box 1066 0 36000 36000
use tholin_avalonsemi_tbb1143  tholin_avalonsemi_tbb1143
timestamp 0
transform 1 0 400000 0 1 305000
box 1066 2048 30000 30000
use tt2_tholin_diceroll  tt2_tholin_diceroll
timestamp 0
transform 1 0 470000 0 1 432000
box 1066 0 21043 22000
use tt2_tholin_multiplexed_counter  tt2_tholin_multiplexed_counter
timestamp 0
transform 1 0 550000 0 1 360000
box 842 0 17098 18000
use tt2_tholin_multiplier  tt2_tholin_multiplier
timestamp 0
transform 1 0 450000 0 1 500000
box 0 0 11118 16584
use tt2_tholin_namebadge  tt2_tholin_namebadge
timestamp 0
transform 1 0 420000 0 1 420000
box 1066 0 23987 25000
use tune_player  tune_player
timestamp 0
transform 1 0 540000 0 1 30000
box 0 2128 21043 19632
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 410000 0 1 120000
box 1066 1504 40000 40000
use wrapped_MC14500  wrapped_MC14500
timestamp 0
transform 1 0 480000 0 1 500000
box 566 0 12000 18000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 480000 0 1 80000
box 1066 2128 60000 60000
use wrapped_as2650  wrapped_as2650
timestamp 0
transform 1 0 460000 0 1 600000
box 0 0 68816 67992
use wrapped_as512512512  wrapped_as512512512
timestamp 0
transform 1 0 20000 0 1 45000
box 1066 2128 340000 637616
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 674393 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 674393 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 674393 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 674393 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 674393 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 674393 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 674393 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 674393 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 49367 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 674393 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 127767 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 157249 434414 422599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 442833 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 385580 470414 598927 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 668393 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 82599 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 139281 506414 201919 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 259417 506414 598927 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 668393 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 425068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 460836 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 674393 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 674393 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 674393 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 674393 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 674393 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 674393 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 674393 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 674393 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 49367 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 674393 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 127767 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 157249 441854 422599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 442833 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 259417 477854 322287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 385225 477854 598927 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 668393 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 82599 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 139281 513854 201919 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 259417 513854 598927 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 668393 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 49367 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 259417 485294 322068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 385580 485294 500068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 517884 485294 598927 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 82599 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 139281 521294 201919 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 259417 521294 598927 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 360068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 377884 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 45068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 49367 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 127767 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 157249 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 500068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 517884 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 259417 492734 322287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 385225 492734 598927 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 668393 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 82599 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 259417 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 360068 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 377884 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 49367 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 127767 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 157249 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 517884 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 139281 489014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 259417 489014 322287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 453692 489014 500068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 517884 489014 598927 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 668393 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 82599 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 139281 525014 201919 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 259417 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 30068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 51692 561014 360068 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 377884 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 674393 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 674393 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 674393 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 674393 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 674393 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 674393 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 674393 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 45068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 49367 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 674393 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 127767 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 157249 424454 420068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 444412 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 500068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 517884 460454 598927 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 668393 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 259417 496454 598927 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 668393 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 82599 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 139281 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 674393 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 674393 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 674393 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 674393 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 674393 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 674393 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 674393 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 674393 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 49367 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 674393 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 127767 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 157249 438134 420068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 444412 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 453692 474134 598927 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 668393 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 82599 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 139281 510134 201919 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 259417 510134 598927 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 668393 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 30068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 51692 546134 446095 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 457897 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 674393 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 674393 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 674393 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 674393 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 684676 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 674393 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 674393 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 45068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 684676 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 49367 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 674393 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 120068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 159644 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 259417 481574 322287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 453692 481574 598927 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 668393 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 82599 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 139281 517574 201919 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 259417 517574 598927 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 668393 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 30068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 51692 553574 360068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 377884 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 331568 651336 331568 651336 0 vccd1
rlabel via4 333704 46776 333704 46776 0 vccd2
rlabel via4 485144 126216 485144 126216 0 vdda1
rlabel via4 528584 637656 528584 637656 0 vdda2
rlabel via4 20864 669936 20864 669936 0 vssa1
rlabel via4 352304 677376 352304 677376 0 vssa2
rlabel via4 346928 655056 346928 655056 0 vssd1
rlabel via4 481424 122496 481424 122496 0 vssd2
rlabel metal1 423062 447542 423062 447542 0 design_clk
rlabel metal2 411624 159868 411624 159868 0 dsi_all\[0\]
rlabel metal1 444222 331330 444222 331330 0 dsi_all\[10\]
rlabel metal2 447166 331585 447166 331585 0 dsi_all\[11\]
rlabel metal3 448784 332588 448784 332588 0 dsi_all\[12\]
rlabel metal1 445464 332622 445464 332622 0 dsi_all\[13\]
rlabel metal2 447166 333387 447166 333387 0 dsi_all\[14\]
rlabel metal2 447258 334305 447258 334305 0 dsi_all\[15\]
rlabel metal1 444912 334050 444912 334050 0 dsi_all\[16\]
rlabel metal2 447166 335699 447166 335699 0 dsi_all\[17\]
rlabel metal2 447258 336005 447258 336005 0 dsi_all\[18\]
rlabel metal2 447166 337059 447166 337059 0 dsi_all\[19\]
rlabel metal3 450156 503423 450156 503423 0 dsi_all\[1\]
rlabel metal2 431250 304334 431250 304334 0 dsi_all\[20\]
rlabel metal2 447166 338453 447166 338453 0 dsi_all\[21\]
rlabel metal2 385710 316030 385710 316030 0 dsi_all\[22\]
rlabel metal1 445510 339558 445510 339558 0 dsi_all\[23\]
rlabel metal2 447166 340119 447166 340119 0 dsi_all\[24\]
rlabel metal2 447166 341207 447166 341207 0 dsi_all\[25\]
rlabel metal2 447258 341513 447258 341513 0 dsi_all\[26\]
rlabel metal3 449060 325788 449060 325788 0 dsi_all\[2\]
rlabel metal1 407928 160514 407928 160514 0 dsi_all\[3\]
rlabel metal2 425116 159732 425116 159732 0 dsi_all\[4\]
rlabel metal1 409722 160310 409722 160310 0 dsi_all\[5\]
rlabel metal2 431496 159868 431496 159868 0 dsi_all\[6\]
rlabel metal3 448646 329188 448646 329188 0 dsi_all\[7\]
rlabel metal3 448876 329868 448876 329868 0 dsi_all\[8\]
rlabel metal1 443670 330582 443670 330582 0 dsi_all\[9\]
rlabel metal2 488697 322116 488697 322116 0 dso_6502\[0\]
rlabel via2 452594 135133 452594 135133 0 dso_6502\[10\]
rlabel via2 452594 136493 452594 136493 0 dso_6502\[11\]
rlabel via2 452594 137853 452594 137853 0 dso_6502\[12\]
rlabel metal2 452594 139281 452594 139281 0 dso_6502\[13\]
rlabel metal2 452134 140607 452134 140607 0 dso_6502\[14\]
rlabel via2 452594 141933 452594 141933 0 dso_6502\[15\]
rlabel metal1 476284 271286 476284 271286 0 dso_6502\[16\]
rlabel via2 452594 144653 452594 144653 0 dso_6502\[17\]
rlabel metal2 452594 146081 452594 146081 0 dso_6502\[18\]
rlabel metal1 476146 275366 476146 275366 0 dso_6502\[19\]
rlabel metal2 489026 299380 489026 299380 0 dso_6502\[1\]
rlabel metal1 473110 315350 473110 315350 0 dso_6502\[20\]
rlabel metal3 451160 150076 451160 150076 0 dso_6502\[21\]
rlabel metal1 476146 272510 476146 272510 0 dso_6502\[22\]
rlabel metal2 452134 152881 452134 152881 0 dso_6502\[23\]
rlabel metal3 451022 154156 451022 154156 0 dso_6502\[24\]
rlabel metal3 450976 155516 450976 155516 0 dso_6502\[25\]
rlabel via2 452594 156893 452594 156893 0 dso_6502\[26\]
rlabel metal2 489249 322116 489249 322116 0 dso_6502\[2\]
rlabel metal2 489525 322116 489525 322116 0 dso_6502\[3\]
rlabel metal1 489348 319090 489348 319090 0 dso_6502\[4\]
rlabel metal1 471178 275298 471178 275298 0 dso_6502\[5\]
rlabel metal1 471362 268430 471362 268430 0 dso_6502\[6\]
rlabel via2 452594 131053 452594 131053 0 dso_6502\[7\]
rlabel metal1 472282 309774 472282 309774 0 dso_6502\[8\]
rlabel via2 452502 133773 452502 133773 0 dso_6502\[9\]
rlabel metal2 503785 385900 503785 385900 0 dso_LCD\[0\]
rlabel metal2 504337 385900 504337 385900 0 dso_LCD\[1\]
rlabel metal2 505310 388576 505310 388576 0 dso_LCD\[2\]
rlabel metal2 506046 389256 506046 389256 0 dso_LCD\[3\]
rlabel metal2 506637 385900 506637 385900 0 dso_LCD\[4\]
rlabel metal2 507281 385900 507281 385900 0 dso_LCD\[5\]
rlabel metal2 508063 385900 508063 385900 0 dso_LCD\[6\]
rlabel metal2 508753 385900 508753 385900 0 dso_LCD\[7\]
rlabel metal3 540492 82348 540492 82348 0 dso_as1802\[0\]
rlabel metal3 540630 102748 540630 102748 0 dso_as1802\[10\]
rlabel metal3 539948 104705 539948 104705 0 dso_as1802\[11\]
rlabel metal3 540676 106828 540676 106828 0 dso_as1802\[12\]
rlabel metal3 539948 108785 539948 108785 0 dso_as1802\[13\]
rlabel metal3 540722 110908 540722 110908 0 dso_as1802\[14\]
rlabel via2 539741 113220 539741 113220 0 dso_as1802\[15\]
rlabel metal3 540078 114988 540078 114988 0 dso_as1802\[16\]
rlabel metal3 540768 117028 540768 117028 0 dso_as1802\[17\]
rlabel metal3 540538 119068 540538 119068 0 dso_as1802\[18\]
rlabel metal3 540124 121108 540124 121108 0 dso_as1802\[19\]
rlabel metal3 541343 84388 541343 84388 0 dso_as1802\[1\]
rlabel metal3 540170 123148 540170 123148 0 dso_as1802\[20\]
rlabel metal2 501354 315039 501354 315039 0 dso_as1802\[21\]
rlabel metal3 541075 137836 541075 137836 0 dso_as1802\[22\]
rlabel metal3 541550 129268 541550 129268 0 dso_as1802\[23\]
rlabel metal1 541052 139230 541052 139230 0 dso_as1802\[24\]
rlabel metal3 541366 133348 541366 133348 0 dso_as1802\[25\]
rlabel metal1 539258 136578 539258 136578 0 dso_as1802\[26\]
rlabel via2 539603 86836 539603 86836 0 dso_as1802\[2\]
rlabel metal3 541458 88468 541458 88468 0 dso_as1802\[3\]
rlabel metal3 541320 90508 541320 90508 0 dso_as1802\[4\]
rlabel metal3 540584 92548 540584 92548 0 dso_as1802\[5\]
rlabel metal3 541412 94588 541412 94588 0 dso_as1802\[6\]
rlabel metal3 541274 96628 541274 96628 0 dso_as1802\[7\]
rlabel via2 539925 99212 539925 99212 0 dso_as1802\[8\]
rlabel metal3 541228 100708 541228 100708 0 dso_as1802\[9\]
rlabel metal2 463121 385900 463121 385900 0 dso_as2650\[0\]
rlabel metal3 459732 626348 459732 626348 0 dso_as2650\[10\]
rlabel metal2 471217 385900 471217 385900 0 dso_as2650\[11\]
rlabel metal2 472190 387471 472190 387471 0 dso_as2650\[12\]
rlabel metal2 472926 389239 472926 389239 0 dso_as2650\[13\]
rlabel metal3 459525 636140 459525 636140 0 dso_as2650\[14\]
rlabel metal3 459502 638588 459502 638588 0 dso_as2650\[15\]
rlabel metal2 468510 494258 468510 494258 0 dso_as2650\[16\]
rlabel metal3 459548 643484 459548 643484 0 dso_as2650\[17\]
rlabel metal2 461610 494394 461610 494394 0 dso_as2650\[18\]
rlabel metal1 458942 602786 458942 602786 0 dso_as2650\[19\]
rlabel metal2 463903 385900 463903 385900 0 dso_as2650\[1\]
rlabel metal2 468602 493544 468602 493544 0 dso_as2650\[20\]
rlabel metal2 461794 492558 461794 492558 0 dso_as2650\[21\]
rlabel metal2 459172 602684 459172 602684 0 dso_as2650\[22\]
rlabel metal2 480286 387318 480286 387318 0 dso_as2650\[23\]
rlabel metal2 481022 387386 481022 387386 0 dso_as2650\[24\]
rlabel metal2 481758 387284 481758 387284 0 dso_as2650\[25\]
rlabel metal2 482494 387182 482494 387182 0 dso_as2650\[26\]
rlabel metal2 464593 385900 464593 385900 0 dso_as2650\[2\]
rlabel metal2 465375 385900 465375 385900 0 dso_as2650\[3\]
rlabel metal2 466111 385900 466111 385900 0 dso_as2650\[4\]
rlabel metal2 466755 385900 466755 385900 0 dso_as2650\[5\]
rlabel metal2 467537 385900 467537 385900 0 dso_as2650\[6\]
rlabel metal2 468273 385900 468273 385900 0 dso_as2650\[7\]
rlabel metal2 469246 387522 469246 387522 0 dso_as2650\[8\]
rlabel metal2 469745 385900 469745 385900 0 dso_as2650\[9\]
rlabel metal2 429226 367778 429226 367778 0 dso_as512512512\[0\]
rlabel metal2 447350 371943 447350 371943 0 dso_as512512512\[10\]
rlabel metal2 447166 372249 447166 372249 0 dso_as512512512\[11\]
rlabel metal2 447350 373303 447350 373303 0 dso_as512512512\[12\]
rlabel metal2 447166 373677 447166 373677 0 dso_as512512512\[13\]
rlabel metal2 411930 449854 411930 449854 0 dso_as512512512\[14\]
rlabel metal2 410550 455396 410550 455396 0 dso_as512512512\[15\]
rlabel metal2 407790 461550 407790 461550 0 dso_as512512512\[16\]
rlabel metal2 447166 376397 447166 376397 0 dso_as512512512\[17\]
rlabel metal2 447350 377451 447350 377451 0 dso_as512512512\[18\]
rlabel metal2 367770 478856 367770 478856 0 dso_as512512512\[19\]
rlabel metal1 444866 365602 444866 365602 0 dso_as512512512\[1\]
rlabel metal2 370714 485078 370714 485078 0 dso_as512512512\[20\]
rlabel metal2 371910 490586 371910 490586 0 dso_as512512512\[21\]
rlabel metal2 406410 496740 406410 496740 0 dso_as512512512\[22\]
rlabel metal2 447534 380511 447534 380511 0 dso_as512512512\[23\]
rlabel metal2 403650 507790 403650 507790 0 dso_as512512512\[24\]
rlabel metal2 447350 381871 447350 381871 0 dso_as512512512\[25\]
rlabel metal2 447166 382177 447166 382177 0 dso_as512512512\[26\]
rlabel metal2 447350 383265 447350 383265 0 dso_as512512512\[27\]
rlabel metal2 447166 366469 447166 366469 0 dso_as512512512\[2\]
rlabel metal1 444820 366962 444820 366962 0 dso_as512512512\[3\]
rlabel metal2 447350 367863 447350 367863 0 dso_as512512512\[4\]
rlabel metal2 447166 368169 447166 368169 0 dso_as512512512\[5\]
rlabel metal2 447350 369189 447350 369189 0 dso_as512512512\[6\]
rlabel metal2 447166 369563 447166 369563 0 dso_as512512512\[7\]
rlabel metal2 447350 370583 447350 370583 0 dso_as512512512\[8\]
rlabel metal2 447166 370889 447166 370889 0 dso_as512512512\[9\]
rlabel metal2 483131 385900 483131 385900 0 dso_as5401\[0\]
rlabel metal2 490590 387862 490590 387862 0 dso_as5401\[10\]
rlabel metal2 535203 425068 535203 425068 0 dso_as5401\[11\]
rlabel metal2 491825 385900 491825 385900 0 dso_as5401\[12\]
rlabel metal2 537779 425068 537779 425068 0 dso_as5401\[13\]
rlabel metal2 539067 425068 539067 425068 0 dso_as5401\[14\]
rlabel metal2 540355 425068 540355 425068 0 dso_as5401\[15\]
rlabel metal2 541834 422630 541834 422630 0 dso_as5401\[16\]
rlabel metal2 542931 425068 542931 425068 0 dso_as5401\[17\]
rlabel metal2 544219 425068 544219 425068 0 dso_as5401\[18\]
rlabel metal2 545698 424092 545698 424092 0 dso_as5401\[19\]
rlabel metal2 483966 387454 483966 387454 0 dso_as5401\[1\]
rlabel metal2 546795 425068 546795 425068 0 dso_as5401\[20\]
rlabel metal2 498449 385900 498449 385900 0 dso_as5401\[21\]
rlabel metal2 522330 406198 522330 406198 0 dso_as5401\[22\]
rlabel metal2 499921 385900 499921 385900 0 dso_as5401\[23\]
rlabel metal2 500894 387386 500894 387386 0 dso_as5401\[24\]
rlabel metal2 501393 385900 501393 385900 0 dso_as5401\[25\]
rlabel metal2 502366 387352 502366 387352 0 dso_as5401\[26\]
rlabel metal2 484702 387318 484702 387318 0 dso_as5401\[2\]
rlabel metal2 485438 387284 485438 387284 0 dso_as5401\[3\]
rlabel metal2 485983 385900 485983 385900 0 dso_as5401\[4\]
rlabel metal2 486910 387250 486910 387250 0 dso_as5401\[5\]
rlabel metal2 487409 385900 487409 385900 0 dso_as5401\[6\]
rlabel metal2 488382 387216 488382 387216 0 dso_as5401\[7\]
rlabel metal2 488881 385900 488881 385900 0 dso_as5401\[8\]
rlabel metal2 489854 387182 489854 387182 0 dso_as5401\[9\]
rlabel metal2 522330 369580 522330 369580 0 dso_counter\[0\]
rlabel metal2 547170 371314 547170 371314 0 dso_counter\[10\]
rlabel metal2 567042 359458 567042 359458 0 dso_counter\[11\]
rlabel metal3 511650 379236 511650 379236 0 dso_counter\[1\]
rlabel metal2 544410 369274 544410 369274 0 dso_counter\[2\]
rlabel metal3 511006 380324 511006 380324 0 dso_counter\[3\]
rlabel metal3 511420 380868 511420 380868 0 dso_counter\[4\]
rlabel metal2 558210 359560 558210 359560 0 dso_counter\[5\]
rlabel metal2 547262 367268 547262 367268 0 dso_counter\[6\]
rlabel metal2 561154 359254 561154 359254 0 dso_counter\[7\]
rlabel metal2 562626 359322 562626 359322 0 dso_counter\[8\]
rlabel metal2 519662 370566 519662 370566 0 dso_counter\[9\]
rlabel metal2 456734 387386 456734 387386 0 dso_diceroll\[0\]
rlabel metal2 457233 385900 457233 385900 0 dso_diceroll\[1\]
rlabel metal2 458206 390616 458206 390616 0 dso_diceroll\[2\]
rlabel metal2 458705 385900 458705 385900 0 dso_diceroll\[3\]
rlabel metal1 481620 429182 481620 429182 0 dso_diceroll\[4\]
rlabel metal1 484334 429182 484334 429182 0 dso_diceroll\[5\]
rlabel metal2 461150 387862 461150 387862 0 dso_diceroll\[6\]
rlabel metal2 461886 387488 461886 387488 0 dso_diceroll\[7\]
rlabel metal3 448968 352308 448968 352308 0 dso_mc14500\[0\]
rlabel via2 450317 353260 450317 353260 0 dso_mc14500\[1\]
rlabel metal3 449014 353668 449014 353668 0 dso_mc14500\[2\]
rlabel metal3 449796 354348 449796 354348 0 dso_mc14500\[3\]
rlabel metal2 484902 500140 484902 500140 0 dso_mc14500\[4\]
rlabel metal2 486512 500140 486512 500140 0 dso_mc14500\[5\]
rlabel metal2 487478 500140 487478 500140 0 dso_mc14500\[6\]
rlabel metal2 488766 500140 488766 500140 0 dso_mc14500\[7\]
rlabel metal3 449566 357748 449566 357748 0 dso_mc14500\[8\]
rlabel metal2 450793 385900 450793 385900 0 dso_multiplier\[0\]
rlabel metal2 451437 385900 451437 385900 0 dso_multiplier\[1\]
rlabel metal2 452081 385900 452081 385900 0 dso_multiplier\[2\]
rlabel metal2 452955 385900 452955 385900 0 dso_multiplier\[3\]
rlabel metal2 453790 387522 453790 387522 0 dso_multiplier\[4\]
rlabel metal2 454289 385900 454289 385900 0 dso_multiplier\[5\]
rlabel metal2 455025 385900 455025 385900 0 dso_multiplier\[6\]
rlabel metal2 461058 498518 461058 498518 0 dso_multiplier\[7\]
rlabel metal2 487370 319610 487370 319610 0 dso_posit\[0\]
rlabel metal2 487593 322116 487593 322116 0 dso_posit\[1\]
rlabel metal1 487554 319294 487554 319294 0 dso_posit\[2\]
rlabel metal2 487968 319124 487968 319124 0 dso_posit\[3\]
rlabel metal2 447166 358955 447166 358955 0 dso_tbb1143\[0\]
rlabel metal2 447350 359329 447350 359329 0 dso_tbb1143\[1\]
rlabel metal1 444866 360298 444866 360298 0 dso_tbb1143\[2\]
rlabel metal2 447166 360689 447166 360689 0 dso_tbb1143\[3\]
rlabel metal2 447166 361709 447166 361709 0 dso_tbb1143\[4\]
rlabel metal1 444820 361658 444820 361658 0 dso_tbb1143\[5\]
rlabel metal2 447166 363103 447166 363103 0 dso_tbb1143\[6\]
rlabel metal2 447350 363409 447350 363409 0 dso_tbb1143\[7\]
rlabel metal3 540684 48635 540684 48635 0 dso_tune
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 461886 320484 461886 320484 0 io_in[10]
rlabel metal3 582046 511292 582046 511292 0 io_in[11]
rlabel metal2 579922 563703 579922 563703 0 io_in[12]
rlabel metal3 581908 617508 581908 617508 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal2 559682 701685 559682 701685 0 io_in[15]
rlabel metal2 444222 371433 444222 371433 0 io_in[16]
rlabel metal2 429870 702178 429870 702178 0 io_in[17]
rlabel metal2 365010 702144 365010 702144 0 io_in[18]
rlabel metal2 449374 503982 449374 503982 0 io_in[19]
rlabel metal2 563730 175644 563730 175644 0 io_in[1]
rlabel metal2 235198 702076 235198 702076 0 io_in[20]
rlabel metal3 444199 421940 444199 421940 0 io_in[21]
rlabel metal2 445142 510476 445142 510476 0 io_in[22]
rlabel metal2 40526 701957 40526 701957 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 2016 632060 2016 632060 0 io_in[25]
rlabel metal3 1786 579972 1786 579972 0 io_in[26]
rlabel metal3 2154 527884 2154 527884 0 io_in[27]
rlabel metal2 3542 678436 3542 678436 0 io_in[28]
rlabel metal3 2016 423572 2016 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal3 2154 371348 2154 371348 0 io_in[30]
rlabel metal1 389804 215322 389804 215322 0 io_in[31]
rlabel metal2 20930 59959 20930 59959 0 io_in[32]
rlabel metal3 2108 214948 2108 214948 0 io_in[33]
rlabel metal3 2200 162860 2200 162860 0 io_in[34]
rlabel metal3 1855 110636 1855 110636 0 io_in[35]
rlabel metal3 1878 71604 1878 71604 0 io_in[36]
rlabel metal3 1924 32436 1924 32436 0 io_in[37]
rlabel metal2 580198 126463 580198 126463 0 io_in[3]
rlabel metal2 580198 166413 580198 166413 0 io_in[4]
rlabel metal3 581218 205700 581218 205700 0 io_in[5]
rlabel via2 580198 245565 580198 245565 0 io_in[6]
rlabel metal2 461610 308890 461610 308890 0 io_in[7]
rlabel metal2 580198 352019 580198 352019 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel metal2 565110 169592 565110 169592 0 io_oeb[0]
rlabel metal2 580198 484517 580198 484517 0 io_oeb[10]
rlabel metal2 580198 537319 580198 537319 0 io_oeb[11]
rlabel metal2 580198 590835 580198 590835 0 io_oeb[12]
rlabel metal3 581954 644028 581954 644028 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal3 523411 465732 523411 465732 0 io_oeb[15]
rlabel metal2 445694 354841 445694 354841 0 io_oeb[16]
rlabel metal2 397486 519802 397486 519802 0 io_oeb[17]
rlabel metal1 331890 703018 331890 703018 0 io_oeb[18]
rlabel metal2 446522 502758 446522 502758 0 io_oeb[19]
rlabel metal2 580198 73049 580198 73049 0 io_oeb[1]
rlabel metal4 449604 510884 449604 510884 0 io_oeb[20]
rlabel metal2 137172 703596 137172 703596 0 io_oeb[21]
rlabel metal2 445234 511003 445234 511003 0 io_oeb[22]
rlabel metal2 446798 502605 446798 502605 0 io_oeb[23]
rlabel metal3 2039 658172 2039 658172 0 io_oeb[24]
rlabel metal3 1855 606084 1855 606084 0 io_oeb[25]
rlabel metal3 2200 553860 2200 553860 0 io_oeb[26]
rlabel metal3 2062 501772 2062 501772 0 io_oeb[27]
rlabel metal3 1924 449548 1924 449548 0 io_oeb[28]
rlabel metal1 5336 61302 5336 61302 0 io_oeb[29]
rlabel metal2 579830 112965 579830 112965 0 io_oeb[2]
rlabel metal1 5520 57902 5520 57902 0 io_oeb[30]
rlabel metal3 1970 293148 1970 293148 0 io_oeb[31]
rlabel metal3 2016 241060 2016 241060 0 io_oeb[32]
rlabel metal3 2154 188836 2154 188836 0 io_oeb[33]
rlabel metal3 1786 136748 1786 136748 0 io_oeb[34]
rlabel metal3 2039 84660 2039 84660 0 io_oeb[35]
rlabel metal3 1878 45492 1878 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580198 152915 580198 152915 0 io_oeb[3]
rlabel metal2 580198 192831 580198 192831 0 io_oeb[4]
rlabel metal2 580014 232781 580014 232781 0 io_oeb[5]
rlabel metal2 580198 272697 580198 272697 0 io_oeb[6]
rlabel metal2 580198 322609 580198 322609 0 io_oeb[7]
rlabel metal2 580198 378301 580198 378301 0 io_oeb[8]
rlabel metal3 582138 431596 582138 431596 0 io_oeb[9]
rlabel metal2 580014 20213 580014 20213 0 io_out[0]
rlabel metal2 469154 321956 469154 321956 0 io_out[10]
rlabel metal3 582000 524484 582000 524484 0 io_out[11]
rlabel metal3 581954 577660 581954 577660 0 io_out[12]
rlabel metal2 469982 321752 469982 321752 0 io_out[13]
rlabel metal2 470258 321786 470258 321786 0 io_out[14]
rlabel metal2 470534 321004 470534 321004 0 io_out[15]
rlabel metal2 442842 365685 442842 365685 0 io_out[16]
rlabel metal2 449466 327964 449466 327964 0 io_out[17]
rlabel metal2 348818 702110 348818 702110 0 io_out[18]
rlabel metal4 444268 505240 444268 505240 0 io_out[19]
rlabel metal2 580198 60163 580198 60163 0 io_out[1]
rlabel metal2 219006 702042 219006 702042 0 io_out[20]
rlabel metal2 153226 697228 153226 697228 0 io_out[21]
rlabel metal2 88366 693845 88366 693845 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal1 3542 678436 3542 678436 0 io_out[24]
rlabel metal3 1947 619140 1947 619140 0 io_out[25]
rlabel metal3 1832 566916 1832 566916 0 io_out[26]
rlabel metal3 2108 514828 2108 514828 0 io_out[27]
rlabel metal3 1878 462604 1878 462604 0 io_out[28]
rlabel metal3 2154 410516 2154 410516 0 io_out[29]
rlabel metal2 580198 100079 580198 100079 0 io_out[2]
rlabel metal1 370484 56338 370484 56338 0 io_out[30]
rlabel metal2 21344 55284 21344 55284 0 io_out[31]
rlabel metal3 1924 254116 1924 254116 0 io_out[32]
rlabel metal3 2062 201892 2062 201892 0 io_out[33]
rlabel metal3 1832 149804 1832 149804 0 io_out[34]
rlabel metal3 1947 97580 1947 97580 0 io_out[35]
rlabel metal3 1970 58548 1970 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel via2 580198 139349 580198 139349 0 io_out[3]
rlabel metal2 580198 179265 580198 179265 0 io_out[4]
rlabel metal2 580198 219215 580198 219215 0 io_out[5]
rlabel metal2 467997 322116 467997 322116 0 io_out[6]
rlabel metal2 580198 312647 580198 312647 0 io_out[7]
rlabel metal2 580198 364735 580198 364735 0 io_out[8]
rlabel metal2 468878 320664 468878 320664 0 io_out[9]
rlabel metal2 488106 292973 488106 292973 0 oeb_6502
rlabel via2 539373 137700 539373 137700 0 oeb_as1802
rlabel metal2 462622 387522 462622 387522 0 oeb_as2650
rlabel via2 447166 383571 447166 383571 0 oeb_as512512512
rlabel metal2 502865 385900 502865 385900 0 oeb_as5401
rlabel metal3 449290 358428 449290 358428 0 oeb_mc14500
rlabel metal2 448010 159868 448010 159868 0 rst_6502
rlabel via1 427754 444533 427754 444533 0 rst_LCD
rlabel metal3 449888 345508 449888 345508 0 rst_as1802
rlabel via2 450133 346324 450133 346324 0 rst_as2650
rlabel metal2 447166 347633 447166 347633 0 rst_as512512512
rlabel via2 450179 347276 450179 347276 0 rst_as5401
rlabel via2 450363 348636 450363 348636 0 rst_counter
rlabel via2 450685 349044 450685 349044 0 rst_diceroll
rlabel metal3 450087 349996 450087 349996 0 rst_mc14500
rlabel metal3 449934 350268 449934 350268 0 rst_posit
rlabel metal2 447166 350761 447166 350761 0 rst_tbb1143
rlabel metal3 450041 351084 450041 351084 0 rst_tune
rlabel metal2 598 1843 598 1843 0 wb_clk_i
rlabel metal2 1702 1911 1702 1911 0 wb_rst_i
rlabel metal2 2898 1214 2898 1214 0 wbs_ack_o
rlabel metal2 409262 175559 409262 175559 0 wbs_adr_i[0]
rlabel metal2 409170 175576 409170 175576 0 wbs_adr_i[10]
rlabel metal2 406778 175576 406778 175576 0 wbs_adr_i[11]
rlabel metal1 255070 44846 255070 44846 0 wbs_adr_i[12]
rlabel metal2 58236 16560 58236 16560 0 wbs_adr_i[13]
rlabel metal2 61863 340 61863 340 0 wbs_adr_i[14]
rlabel metal2 406410 175440 406410 175440 0 wbs_adr_i[15]
rlabel metal2 406686 175508 406686 175508 0 wbs_adr_i[16]
rlabel metal2 404018 175372 404018 175372 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 403926 172431 403926 172431 0 wbs_adr_i[1]
rlabel metal2 83076 16560 83076 16560 0 wbs_adr_i[20]
rlabel metal2 86703 340 86703 340 0 wbs_adr_i[21]
rlabel metal2 90153 340 90153 340 0 wbs_adr_i[22]
rlabel metal2 93978 3627 93978 3627 0 wbs_adr_i[23]
rlabel metal2 97060 16560 97060 16560 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 104321 340 104321 340 0 wbs_adr_i[26]
rlabel metal1 253046 44642 253046 44642 0 wbs_adr_i[27]
rlabel metal2 111642 1792 111642 1792 0 wbs_adr_i[28]
rlabel metal2 114993 340 114993 340 0 wbs_adr_i[29]
rlabel metal2 17066 1962 17066 1962 0 wbs_adr_i[2]
rlabel metal2 118818 3627 118818 3627 0 wbs_adr_i[30]
rlabel metal2 121900 16560 121900 16560 0 wbs_adr_i[31]
rlabel metal2 21298 16560 21298 16560 0 wbs_adr_i[3]
rlabel metal2 26397 340 26397 340 0 wbs_adr_i[4]
rlabel metal2 450570 159426 450570 159426 0 wbs_adr_i[5]
rlabel metal2 450846 176664 450846 176664 0 wbs_adr_i[6]
rlabel metal2 36977 340 36977 340 0 wbs_adr_i[7]
rlabel metal2 40473 340 40473 340 0 wbs_adr_i[8]
rlabel metal2 44298 3627 44298 3627 0 wbs_adr_i[9]
rlabel metal2 3857 340 3857 340 0 wbs_cyc_i
rlabel metal2 392610 151844 392610 151844 0 wbs_dat_i[0]
rlabel metal2 392702 152048 392702 152048 0 wbs_dat_i[10]
rlabel metal2 52578 2234 52578 2234 0 wbs_dat_i[11]
rlabel metal2 55660 16560 55660 16560 0 wbs_dat_i[12]
rlabel metal2 59517 340 59517 340 0 wbs_dat_i[13]
rlabel metal2 62698 16560 62698 16560 0 wbs_dat_i[14]
rlabel metal2 392886 167314 392886 167314 0 wbs_dat_i[15]
rlabel metal2 390218 167246 390218 167246 0 wbs_dat_i[16]
rlabel metal2 390034 167042 390034 167042 0 wbs_dat_i[17]
rlabel metal2 77418 3627 77418 3627 0 wbs_dat_i[18]
rlabel metal2 80500 16560 80500 16560 0 wbs_dat_i[19]
rlabel metal2 389850 150501 389850 150501 0 wbs_dat_i[1]
rlabel metal2 390126 167348 390126 167348 0 wbs_dat_i[20]
rlabel metal2 387550 171190 387550 171190 0 wbs_dat_i[21]
rlabel metal2 387366 168776 387366 168776 0 wbs_dat_i[22]
rlabel metal2 94937 340 94937 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102212 16560 102212 16560 0 wbs_dat_i[25]
rlabel metal2 387458 166124 387458 166124 0 wbs_dat_i[26]
rlabel metal2 384514 165716 384514 165716 0 wbs_dat_i[27]
rlabel metal2 384606 168538 384606 168538 0 wbs_dat_i[28]
rlabel metal2 116196 16560 116196 16560 0 wbs_dat_i[29]
rlabel metal2 18117 340 18117 340 0 wbs_dat_i[2]
rlabel metal2 119370 16560 119370 16560 0 wbs_dat_i[30]
rlabel metal2 123273 340 123273 340 0 wbs_dat_i[31]
rlabel metal2 22809 340 22809 340 0 wbs_dat_i[3]
rlabel metal2 27738 2064 27738 2064 0 wbs_dat_i[4]
rlabel metal2 31089 340 31089 340 0 wbs_dat_i[5]
rlabel metal2 519754 315894 519754 315894 0 wbs_dat_i[6]
rlabel metal2 37858 16560 37858 16560 0 wbs_dat_i[7]
rlabel metal2 41676 16560 41676 16560 0 wbs_dat_i[8]
rlabel metal2 45257 340 45257 340 0 wbs_dat_i[9]
rlabel metal2 9837 340 9837 340 0 wbs_dat_o[0]
rlabel metal2 520766 318002 520766 318002 0 wbs_dat_o[10]
rlabel metal2 450662 160106 450662 160106 0 wbs_dat_o[11]
rlabel metal2 57033 340 57033 340 0 wbs_dat_o[12]
rlabel metal2 60858 17398 60858 17398 0 wbs_dat_o[13]
rlabel metal2 63940 16560 63940 16560 0 wbs_dat_o[14]
rlabel metal2 519386 322116 519386 322116 0 wbs_dat_o[15]
rlabel metal1 445648 291754 445648 291754 0 wbs_dat_o[16]
rlabel metal2 74796 16560 74796 16560 0 wbs_dat_o[17]
rlabel metal2 78377 340 78377 340 0 wbs_dat_o[18]
rlabel metal2 82110 2030 82110 2030 0 wbs_dat_o[19]
rlabel metal2 14766 2098 14766 2098 0 wbs_dat_o[1]
rlabel metal2 373290 161602 373290 161602 0 wbs_dat_o[20]
rlabel metal2 373566 161704 373566 161704 0 wbs_dat_o[21]
rlabel metal2 92782 1860 92782 1860 0 wbs_dat_o[22]
rlabel metal2 96041 340 96041 340 0 wbs_dat_o[23]
rlabel metal2 99636 16560 99636 16560 0 wbs_dat_o[24]
rlabel metal2 103362 1826 103362 1826 0 wbs_dat_o[25]
rlabel metal2 370714 161874 370714 161874 0 wbs_dat_o[26]
rlabel metal2 110538 1758 110538 1758 0 wbs_dat_o[27]
rlabel metal2 113620 16560 113620 16560 0 wbs_dat_o[28]
rlabel metal2 117477 340 117477 340 0 wbs_dat_o[29]
rlabel metal2 19412 16560 19412 16560 0 wbs_dat_o[2]
rlabel metal2 120881 340 120881 340 0 wbs_dat_o[30]
rlabel metal2 124706 2166 124706 2166 0 wbs_dat_o[31]
rlabel metal2 24242 1928 24242 1928 0 wbs_dat_o[3]
rlabel metal2 368230 167195 368230 167195 0 wbs_dat_o[4]
rlabel metal2 368138 158882 368138 158882 0 wbs_dat_o[5]
rlabel metal2 36018 2200 36018 2200 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 42957 340 42957 340 0 wbs_dat_o[8]
rlabel metal2 368046 158848 368046 158848 0 wbs_dat_o[9]
rlabel metal2 5290 2115 5290 2115 0 wbs_stb_i
rlabel metal2 6486 2047 6486 2047 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
