VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_MC14500
  CLASS BLOCK ;
  FOREIGN wrapped_MC14500 ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 90.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 86.000 15.230 90.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.580 4.000 9.780 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.260 4.000 27.460 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.620 4.000 62.820 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.300 4.000 80.500 ;
    END
  END io_in[4]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.530 0.000 57.090 4.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 0.000 3.270 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.690 0.000 9.250 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.670 0.000 15.230 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 0.000 21.210 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.630 0.000 27.190 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.610 0.000 33.170 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.590 0.000 39.150 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.570 0.000 45.130 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 0.000 51.110 4.000 ;
    END
  END io_out[8]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.570 86.000 45.130 90.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.815 10.640 12.415 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.005 10.640 24.605 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.195 10.640 36.795 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.385 10.640 48.985 79.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.910 10.640 18.510 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.100 10.640 30.700 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.290 10.640 42.890 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.480 10.640 55.080 79.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 78.965 ;
      LAYER met1 ;
        RECT 2.830 10.640 56.970 79.120 ;
      LAYER met2 ;
        RECT 2.860 85.720 14.390 86.770 ;
        RECT 15.510 85.720 44.290 86.770 ;
        RECT 45.410 85.720 56.940 86.770 ;
        RECT 2.860 4.280 56.940 85.720 ;
        RECT 3.550 4.000 8.410 4.280 ;
        RECT 9.530 4.000 14.390 4.280 ;
        RECT 15.510 4.000 20.370 4.280 ;
        RECT 21.490 4.000 26.350 4.280 ;
        RECT 27.470 4.000 32.330 4.280 ;
        RECT 33.450 4.000 38.310 4.280 ;
        RECT 39.430 4.000 44.290 4.280 ;
        RECT 45.410 4.000 50.270 4.280 ;
        RECT 51.390 4.000 56.250 4.280 ;
      LAYER met3 ;
        RECT 4.400 78.900 55.070 80.065 ;
        RECT 4.000 63.220 55.070 78.900 ;
        RECT 4.400 61.220 55.070 63.220 ;
        RECT 4.000 45.540 55.070 61.220 ;
        RECT 4.400 43.540 55.070 45.540 ;
        RECT 4.000 27.860 55.070 43.540 ;
        RECT 4.400 25.860 55.070 27.860 ;
        RECT 4.000 10.180 55.070 25.860 ;
        RECT 4.400 9.015 55.070 10.180 ;
  END
END wrapped_MC14500
END LIBRARY

