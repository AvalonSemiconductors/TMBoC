// This is the unpowered netlist.
module tholin_avalonsemi_tbb1143 (clk,
    rst,
    io_in,
    io_out);
 input clk;
 input rst;
 input [5:0] io_in;
 output [7:0] io_out;

 wire \CIRCUIT_2223.CLK ;
 wire \CIRCUIT_2223.GATES_1.input1[0] ;
 wire \CIRCUIT_2223.GATES_1.input1[1] ;
 wire \CIRCUIT_2223.GATES_1.input1[2] ;
 wire \CIRCUIT_2223.GATES_1.input1[3] ;
 wire \CIRCUIT_2223.GATES_11.input2 ;
 wire clknet_0_clk;
 wire \CIRCUIT_2223.GATES_2.input2 ;
 wire \CIRCUIT_2223.GATES_3.input2 ;
 wire \CIRCUIT_2223.GATES_4.input1[0] ;
 wire \CIRCUIT_2223.GATES_4.input1[1] ;
 wire \CIRCUIT_2223.GATES_4.input1[2] ;
 wire \CIRCUIT_2223.GATES_4.input1[3] ;
 wire \CIRCUIT_2223.GATES_5.input2 ;
 wire \CIRCUIT_2223.MEMORY_18.clock ;
 wire \CIRCUIT_2223.MEMORY_18.d ;
 wire \CIRCUIT_2223.MEMORY_18.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_19.d ;
 wire \CIRCUIT_2223.MEMORY_19.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_20.d ;
 wire \CIRCUIT_2223.MEMORY_20.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_21.d ;
 wire \CIRCUIT_2223.MEMORY_21.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_22.d ;
 wire \CIRCUIT_2223.MEMORY_22.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_23.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_24.d ;
 wire \CIRCUIT_2223.MEMORY_24.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_25.d ;
 wire \CIRCUIT_2223.MEMORY_25.s_currentState ;
 wire \CIRCUIT_2223.MEMORY_26.s_currentState ;
 wire \CIRCUIT_2223.s_logisimNet48 ;
 wire \CIRCUIT_2223.tone_generator_1.GATES_1.result ;
 wire \CIRCUIT_2223.tone_generator_1.GATES_2.result ;
 wire \CIRCUIT_2223.tone_generator_1.GATES_3.result ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d ;
 wire \CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_27.result ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d ;
 wire \CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_27.result ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d ;
 wire \CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ;
 wire \CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire \slow_clock[0] ;
 wire \slow_clock[1] ;
 wire \slow_clock[2] ;
 wire \slow_clock[3] ;
 wire \slow_clock[4] ;
 wire \slow_clock[5] ;
 wire \slow_clock[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_0__195_;
 wire clknet_1_0__leaf__195_;
 wire clknet_1_1__leaf__195_;
 wire clknet_0__262_;
 wire clknet_1_0__leaf__262_;
 wire clknet_1_1__leaf__262_;
 wire clknet_0__263_;
 wire clknet_1_0__leaf__263_;
 wire clknet_1_1__leaf__263_;
 wire clknet_0__281_;
 wire clknet_1_0__leaf__281_;
 wire clknet_1_1__leaf__281_;
 wire clknet_0__282_;
 wire clknet_1_0__leaf__282_;
 wire clknet_1_1__leaf__282_;
 wire clknet_0__235_;
 wire clknet_1_0__leaf__235_;
 wire clknet_1_1__leaf__235_;
 wire clknet_0__236_;
 wire clknet_1_0__leaf__236_;
 wire clknet_1_1__leaf__236_;
 wire clknet_0__212_;
 wire clknet_1_0__leaf__212_;
 wire clknet_1_1__leaf__212_;
 wire clknet_0__213_;
 wire clknet_1_0__leaf__213_;
 wire clknet_1_1__leaf__213_;
 wire net28;

 sky130_fd_sc_hd__inv_2 _380_ (.A(net18),
    .Y(_117_));
 sky130_fd_sc_hd__clkbuf_4 _381_ (.A(net20),
    .X(_179_));
 sky130_fd_sc_hd__inv_2 _382_ (.A(_179_),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _383_ (.A(_179_),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(_179_),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _385_ (.A(_179_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _386_ (.A(_179_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(_179_),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(_179_),
    .Y(_102_));
 sky130_fd_sc_hd__and4_2 _389_ (.A(net2),
    .B(net1),
    .C(\CIRCUIT_2223.GATES_1.input1[0] ),
    .D(\CIRCUIT_2223.GATES_1.input1[1] ),
    .X(_180_));
 sky130_fd_sc_hd__and4_1 _390_ (.A(net2),
    .B(net1),
    .C(\CIRCUIT_2223.GATES_1.input1[2] ),
    .D(\CIRCUIT_2223.GATES_1.input1[3] ),
    .X(_181_));
 sky130_fd_sc_hd__nand2_2 _391_ (.A(_180_),
    .B(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__mux2_1 _392_ (.A0(net6),
    .A1(\CIRCUIT_2223.s_logisimNet48 ),
    .S(_182_),
    .X(_183_));
 sky130_fd_sc_hd__clkbuf_1 _393_ (.A(_183_),
    .X(_178_));
 sky130_fd_sc_hd__clkbuf_4 _394_ (.A(net5),
    .X(_184_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(_184_),
    .A1(\CIRCUIT_2223.GATES_5.input2 ),
    .S(_182_),
    .X(_185_));
 sky130_fd_sc_hd__clkbuf_1 _396_ (.A(_185_),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_4 _397_ (.A(net4),
    .X(_186_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(_186_),
    .A1(\CIRCUIT_2223.GATES_3.input2 ),
    .S(_182_),
    .X(_187_));
 sky130_fd_sc_hd__clkbuf_1 _399_ (.A(_187_),
    .X(_176_));
 sky130_fd_sc_hd__buf_2 _400_ (.A(net3),
    .X(_188_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(_188_),
    .A1(\CIRCUIT_2223.GATES_2.input2 ),
    .S(_182_),
    .X(_189_));
 sky130_fd_sc_hd__clkbuf_1 _402_ (.A(_189_),
    .X(_175_));
 sky130_fd_sc_hd__nand2_2 _403_ (.A(net18),
    .B(net7),
    .Y(_190_));
 sky130_fd_sc_hd__buf_8 _404_ (.A(_190_),
    .X(_191_));
 sky130_fd_sc_hd__buf_6 _405_ (.A(_191_),
    .X(_000_));
 sky130_fd_sc_hd__o211ai_4 _406_ (.A1(\CIRCUIT_2223.GATES_1.input1[2] ),
    .A2(\CIRCUIT_2223.GATES_1.input1[3] ),
    .B1(net2),
    .C1(net1),
    .Y(_192_));
 sky130_fd_sc_hd__o211ai_4 _407_ (.A1(\CIRCUIT_2223.GATES_1.input1[0] ),
    .A2(\CIRCUIT_2223.GATES_1.input1[1] ),
    .B1(net2),
    .C1(net1),
    .Y(_193_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(\CIRCUIT_2223.MEMORY_23.s_currentState ),
    .Y(\CIRCUIT_2223.GATES_11.input2 ));
 sky130_fd_sc_hd__nand2_2 _410_ (.A(clknet_1_1__leaf_clk),
    .B(\CIRCUIT_2223.GATES_11.input2 ),
    .Y(_195_));
 sky130_fd_sc_hd__xor2_1 _411_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ),
    .X(_196_));
 sky130_fd_sc_hd__xor2_1 _412_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ),
    .X(_197_));
 sky130_fd_sc_hd__xor2_1 _413_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ),
    .X(_198_));
 sky130_fd_sc_hd__xor2_1 _414_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ),
    .X(_199_));
 sky130_fd_sc_hd__or4_1 _415_ (.A(_196_),
    .B(_197_),
    .C(_198_),
    .D(_199_),
    .X(_200_));
 sky130_fd_sc_hd__or2_1 _416_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ),
    .X(_201_));
 sky130_fd_sc_hd__nand2_1 _417_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ),
    .Y(_202_));
 sky130_fd_sc_hd__or2_1 _418_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ),
    .X(_203_));
 sky130_fd_sc_hd__nand2_1 _419_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ),
    .Y(_204_));
 sky130_fd_sc_hd__xor2_1 _420_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ),
    .X(_205_));
 sky130_fd_sc_hd__a221o_1 _421_ (.A1(_201_),
    .A2(_202_),
    .B1(_203_),
    .B2(_204_),
    .C1(_205_),
    .X(_206_));
 sky130_fd_sc_hd__xor2_1 _422_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ),
    .X(_207_));
 sky130_fd_sc_hd__xor2_1 _423_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ),
    .X(_208_));
 sky130_fd_sc_hd__xor2_1 _424_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ),
    .X(_209_));
 sky130_fd_sc_hd__xor2_1 _425_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ),
    .X(_210_));
 sky130_fd_sc_hd__or4_1 _426_ (.A(_207_),
    .B(_208_),
    .C(_209_),
    .D(_210_),
    .X(_211_));
 sky130_fd_sc_hd__nor3_1 _427_ (.A(_200_),
    .B(_206_),
    .C(_211_),
    .Y(\CIRCUIT_2223.tone_generator_2_2.GATES_27.result ));
 sky130_fd_sc_hd__a32o_2 _428_ (.A1(net24),
    .A2(_192_),
    .A3(_194_),
    .B1(clknet_1_1__leaf__195_),
    .B2(\CIRCUIT_2223.tone_generator_2_2.GATES_27.result ),
    .X(_212_));
 sky130_fd_sc_hd__buf_1 _429_ (.A(clknet_1_1__leaf__212_),
    .X(_213_));
 sky130_fd_sc_hd__xor2_2 _430_ (.A(_000_),
    .B(clknet_1_0__leaf__213_),
    .X(_094_));
 sky130_fd_sc_hd__xor2_2 _431_ (.A(_000_),
    .B(clknet_1_0__leaf__213_),
    .X(_092_));
 sky130_fd_sc_hd__xor2_2 _432_ (.A(_000_),
    .B(clknet_1_0__leaf__213_),
    .X(_090_));
 sky130_fd_sc_hd__xor2_2 _433_ (.A(_000_),
    .B(clknet_1_0__leaf__213_),
    .X(_088_));
 sky130_fd_sc_hd__xor2_2 _434_ (.A(_000_),
    .B(clknet_1_0__leaf__213_),
    .X(_086_));
 sky130_fd_sc_hd__buf_8 _435_ (.A(_191_),
    .X(_214_));
 sky130_fd_sc_hd__xor2_2 _436_ (.A(_214_),
    .B(clknet_1_1__leaf__213_),
    .X(_084_));
 sky130_fd_sc_hd__xor2_2 _437_ (.A(_214_),
    .B(clknet_1_1__leaf__213_),
    .X(_081_));
 sky130_fd_sc_hd__xor2_2 _438_ (.A(_214_),
    .B(clknet_1_1__leaf__213_),
    .X(_079_));
 sky130_fd_sc_hd__xor2_2 _439_ (.A(_214_),
    .B(clknet_1_1__leaf__213_),
    .X(_077_));
 sky130_fd_sc_hd__xor2_2 _440_ (.A(_214_),
    .B(clknet_1_1__leaf__213_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_16 _441_ (.A(_190_),
    .X(_215_));
 sky130_fd_sc_hd__xor2_1 _442_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ),
    .X(_216_));
 sky130_fd_sc_hd__xor2_1 _443_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ),
    .X(_217_));
 sky130_fd_sc_hd__xor2_1 _444_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ),
    .X(_218_));
 sky130_fd_sc_hd__xor2_1 _445_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ),
    .X(_219_));
 sky130_fd_sc_hd__or4_1 _446_ (.A(_216_),
    .B(_217_),
    .C(_218_),
    .D(_219_),
    .X(_220_));
 sky130_fd_sc_hd__or2_1 _447_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ),
    .X(_221_));
 sky130_fd_sc_hd__nand2_1 _448_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ),
    .Y(_222_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ),
    .Y(_223_));
 sky130_fd_sc_hd__or2_1 _450_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ),
    .X(_224_));
 sky130_fd_sc_hd__xor2_1 _451_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ),
    .X(_225_));
 sky130_fd_sc_hd__a221o_1 _452_ (.A1(_221_),
    .A2(_222_),
    .B1(_223_),
    .B2(_224_),
    .C1(_225_),
    .X(_226_));
 sky130_fd_sc_hd__xor2_1 _453_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ),
    .X(_227_));
 sky130_fd_sc_hd__xor2_1 _454_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ),
    .X(_228_));
 sky130_fd_sc_hd__xor2_1 _455_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ),
    .X(_229_));
 sky130_fd_sc_hd__xor2_1 _456_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ),
    .X(_230_));
 sky130_fd_sc_hd__or4_1 _457_ (.A(_227_),
    .B(_228_),
    .C(_229_),
    .D(_230_),
    .X(_231_));
 sky130_fd_sc_hd__nor3_1 _458_ (.A(_220_),
    .B(_226_),
    .C(_231_),
    .Y(\CIRCUIT_2223.tone_generator_2_1.GATES_27.result ));
 sky130_fd_sc_hd__and4b_1 _459_ (.A_N(\CIRCUIT_2223.GATES_1.input1[3] ),
    .B(\CIRCUIT_2223.GATES_1.input1[2] ),
    .C(net1),
    .D(net2),
    .X(_232_));
 sky130_fd_sc_hd__clkbuf_2 _460_ (.A(_232_),
    .X(_233_));
 sky130_fd_sc_hd__and3b_1 _461_ (.A_N(_180_),
    .B(_233_),
    .C(net19),
    .X(_234_));
 sky130_fd_sc_hd__a21oi_2 _462_ (.A1(clknet_1_0__leaf__195_),
    .A2(\CIRCUIT_2223.tone_generator_2_1.GATES_27.result ),
    .B1(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__buf_1 _463_ (.A(clknet_1_0__leaf__235_),
    .X(_236_));
 sky130_fd_sc_hd__xnor2_2 _464_ (.A(_215_),
    .B(clknet_1_0__leaf__236_),
    .Y(_073_));
 sky130_fd_sc_hd__xnor2_2 _465_ (.A(_215_),
    .B(clknet_1_0__leaf__236_),
    .Y(_071_));
 sky130_fd_sc_hd__xnor2_2 _466_ (.A(_215_),
    .B(clknet_1_1__leaf__236_),
    .Y(_069_));
 sky130_fd_sc_hd__buf_8 _467_ (.A(_190_),
    .X(_237_));
 sky130_fd_sc_hd__xnor2_2 _468_ (.A(_237_),
    .B(clknet_1_1__leaf__236_),
    .Y(_067_));
 sky130_fd_sc_hd__xnor2_2 _469_ (.A(_237_),
    .B(clknet_1_1__leaf__236_),
    .Y(_065_));
 sky130_fd_sc_hd__xnor2_2 _470_ (.A(_237_),
    .B(clknet_1_1__leaf__236_),
    .Y(_063_));
 sky130_fd_sc_hd__xnor2_2 _471_ (.A(_237_),
    .B(clknet_1_1__leaf__236_),
    .Y(_060_));
 sky130_fd_sc_hd__xnor2_2 _472_ (.A(_237_),
    .B(clknet_1_0__leaf__236_),
    .Y(_058_));
 sky130_fd_sc_hd__xnor2_2 _473_ (.A(_237_),
    .B(clknet_1_0__leaf__236_),
    .Y(_056_));
 sky130_fd_sc_hd__xnor2_2 _474_ (.A(_237_),
    .B(clknet_1_0__leaf__236_),
    .Y(_054_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__nand2_1 _476_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ),
    .Y(_238_));
 sky130_fd_sc_hd__or2_1 _477_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ),
    .X(_239_));
 sky130_fd_sc_hd__or2_1 _478_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ),
    .X(_240_));
 sky130_fd_sc_hd__nand2_1 _479_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ),
    .Y(_241_));
 sky130_fd_sc_hd__xor2_1 _480_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ),
    .X(_242_));
 sky130_fd_sc_hd__a221o_1 _481_ (.A1(_238_),
    .A2(_239_),
    .B1(_240_),
    .B2(_241_),
    .C1(_242_),
    .X(_243_));
 sky130_fd_sc_hd__nand2_1 _482_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ),
    .Y(_244_));
 sky130_fd_sc_hd__or2_1 _483_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ),
    .X(_245_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ),
    .Y(_246_));
 sky130_fd_sc_hd__or2_1 _485_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ),
    .X(_247_));
 sky130_fd_sc_hd__a22o_1 _486_ (.A1(_244_),
    .A2(_245_),
    .B1(_246_),
    .B2(_247_),
    .X(_248_));
 sky130_fd_sc_hd__xor2_1 _487_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ),
    .X(_249_));
 sky130_fd_sc_hd__xor2_1 _488_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ),
    .X(_250_));
 sky130_fd_sc_hd__xor2_1 _489_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ),
    .X(_251_));
 sky130_fd_sc_hd__xor2_1 _490_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ),
    .X(_252_));
 sky130_fd_sc_hd__xor2_1 _491_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ),
    .X(_253_));
 sky130_fd_sc_hd__xor2_1 _492_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ),
    .X(_254_));
 sky130_fd_sc_hd__or4_1 _493_ (.A(_251_),
    .B(_252_),
    .C(_253_),
    .D(_254_),
    .X(_255_));
 sky130_fd_sc_hd__or4_1 _494_ (.A(_248_),
    .B(_249_),
    .C(_250_),
    .D(_255_),
    .X(_256_));
 sky130_fd_sc_hd__inv_2 _495_ (.A(\CIRCUIT_2223.GATES_1.input1[1] ),
    .Y(_257_));
 sky130_fd_sc_hd__and4b_1 _496_ (.A_N(\CIRCUIT_2223.GATES_1.input1[2] ),
    .B(\CIRCUIT_2223.GATES_1.input1[3] ),
    .C(net2),
    .D(net1),
    .X(_258_));
 sky130_fd_sc_hd__clkbuf_2 _497_ (.A(_258_),
    .X(_259_));
 sky130_fd_sc_hd__nand2_2 _498_ (.A(_180_),
    .B(_233_),
    .Y(_260_));
 sky130_fd_sc_hd__a21boi_1 _499_ (.A1(_257_),
    .A2(_259_),
    .B1_N(_260_),
    .Y(_261_));
 sky130_fd_sc_hd__o32a_2 _500_ (.A1(net27),
    .A2(_243_),
    .A3(_256_),
    .B1(_261_),
    .B2(_117_),
    .X(_262_));
 sky130_fd_sc_hd__buf_1 _501_ (.A(clknet_1_0__leaf__262_),
    .X(_263_));
 sky130_fd_sc_hd__xnor2_2 _502_ (.A(_215_),
    .B(clknet_1_1__leaf__263_),
    .Y(_049_));
 sky130_fd_sc_hd__xnor2_2 _503_ (.A(_237_),
    .B(clknet_1_0__leaf__263_),
    .Y(_047_));
 sky130_fd_sc_hd__xnor2_2 _504_ (.A(_237_),
    .B(clknet_1_0__leaf__263_),
    .Y(_045_));
 sky130_fd_sc_hd__xnor2_2 _505_ (.A(_237_),
    .B(clknet_1_0__leaf__263_),
    .Y(_043_));
 sky130_fd_sc_hd__xnor2_2 _506_ (.A(_191_),
    .B(clknet_1_0__leaf__263_),
    .Y(_041_));
 sky130_fd_sc_hd__xnor2_2 _507_ (.A(_191_),
    .B(clknet_1_0__leaf__263_),
    .Y(_039_));
 sky130_fd_sc_hd__xnor2_2 _508_ (.A(_191_),
    .B(clknet_1_1__leaf__263_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_2 _509_ (.A(_191_),
    .B(clknet_1_1__leaf__263_),
    .Y(_034_));
 sky130_fd_sc_hd__xnor2_2 _510_ (.A(_191_),
    .B(clknet_1_1__leaf__263_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_2 _511_ (.A(_191_),
    .B(clknet_1_1__leaf__263_),
    .Y(_030_));
 sky130_fd_sc_hd__xor2_1 _512_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ),
    .X(_264_));
 sky130_fd_sc_hd__xor2_1 _513_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ),
    .X(_265_));
 sky130_fd_sc_hd__xor2_1 _514_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ),
    .X(_266_));
 sky130_fd_sc_hd__xor2_1 _515_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ),
    .X(_267_));
 sky130_fd_sc_hd__or4_1 _516_ (.A(_264_),
    .B(_265_),
    .C(_266_),
    .D(_267_),
    .X(_268_));
 sky130_fd_sc_hd__or2_1 _517_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ),
    .X(_269_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ),
    .Y(_270_));
 sky130_fd_sc_hd__nand2_1 _519_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ),
    .Y(_271_));
 sky130_fd_sc_hd__or2_1 _520_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ),
    .X(_272_));
 sky130_fd_sc_hd__xor2_1 _521_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ),
    .X(_273_));
 sky130_fd_sc_hd__a221o_1 _522_ (.A1(_269_),
    .A2(_270_),
    .B1(_271_),
    .B2(_272_),
    .C1(_273_),
    .X(_274_));
 sky130_fd_sc_hd__xor2_1 _523_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ),
    .X(_275_));
 sky130_fd_sc_hd__xor2_1 _524_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ),
    .X(_276_));
 sky130_fd_sc_hd__xor2_1 _525_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ),
    .X(_277_));
 sky130_fd_sc_hd__xor2_1 _526_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ),
    .X(_278_));
 sky130_fd_sc_hd__or4_1 _527_ (.A(_275_),
    .B(_276_),
    .C(_277_),
    .D(_278_),
    .X(_279_));
 sky130_fd_sc_hd__nor3_1 _528_ (.A(_268_),
    .B(_274_),
    .C(_279_),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ));
 sky130_fd_sc_hd__a22o_1 _529_ (.A1(_181_),
    .A2(_193_),
    .B1(_259_),
    .B2(\CIRCUIT_2223.GATES_1.input1[1] ),
    .X(_280_));
 sky130_fd_sc_hd__a22o_2 _530_ (.A1(clknet_1_1__leaf__195_),
    .A2(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ),
    .B1(_280_),
    .B2(net24),
    .X(_281_));
 sky130_fd_sc_hd__buf_1 _531_ (.A(clknet_1_1__leaf__281_),
    .X(_282_));
 sky130_fd_sc_hd__xor2_2 _532_ (.A(_000_),
    .B(clknet_1_0__leaf__282_),
    .X(_028_));
 sky130_fd_sc_hd__xor2_2 _533_ (.A(_214_),
    .B(clknet_1_0__leaf__282_),
    .X(_026_));
 sky130_fd_sc_hd__xor2_2 _534_ (.A(_214_),
    .B(clknet_1_0__leaf__282_),
    .X(_024_));
 sky130_fd_sc_hd__xor2_2 _535_ (.A(_214_),
    .B(clknet_1_1__leaf__282_),
    .X(_022_));
 sky130_fd_sc_hd__xor2_2 _536_ (.A(_214_),
    .B(clknet_1_0__leaf__282_),
    .X(_019_));
 sky130_fd_sc_hd__xor2_2 _537_ (.A(_214_),
    .B(clknet_1_1__leaf__282_),
    .X(_017_));
 sky130_fd_sc_hd__xor2_2 _538_ (.A(_215_),
    .B(clknet_1_1__leaf__282_),
    .X(_015_));
 sky130_fd_sc_hd__xor2_2 _539_ (.A(_215_),
    .B(clknet_1_1__leaf__282_),
    .X(_013_));
 sky130_fd_sc_hd__xor2_2 _540_ (.A(_215_),
    .B(clknet_1_1__leaf__282_),
    .X(_011_));
 sky130_fd_sc_hd__xor2_2 _541_ (.A(_215_),
    .B(clknet_1_1__leaf__282_),
    .X(_009_));
 sky130_fd_sc_hd__clkinv_2 _542_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock ));
 sky130_fd_sc_hd__clkinv_2 _543_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d ));
 sky130_fd_sc_hd__clkinv_2 _544_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d ));
 sky130_fd_sc_hd__clkinv_2 _545_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d ));
 sky130_fd_sc_hd__clkinv_2 _546_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d ));
 sky130_fd_sc_hd__inv_2 _547_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d ));
 sky130_fd_sc_hd__clkinv_2 _548_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d ));
 sky130_fd_sc_hd__clkinv_2 _549_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d ));
 sky130_fd_sc_hd__clkinv_2 _550_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d ));
 sky130_fd_sc_hd__clkinv_2 _551_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d ));
 sky130_fd_sc_hd__clkinv_2 _552_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d ));
 sky130_fd_sc_hd__clkinv_2 _553_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d ));
 sky130_fd_sc_hd__clkinv_2 _554_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d ));
 sky130_fd_sc_hd__clkinv_2 _555_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d ));
 sky130_fd_sc_hd__clkinv_2 _556_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock ));
 sky130_fd_sc_hd__clkinv_2 _557_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock ));
 sky130_fd_sc_hd__clkinv_2 _558_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d ));
 sky130_fd_sc_hd__clkinv_2 _559_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d ));
 sky130_fd_sc_hd__clkinv_2 _560_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d ));
 sky130_fd_sc_hd__clkinv_2 _561_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d ));
 sky130_fd_sc_hd__clkinv_2 _562_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d ));
 sky130_fd_sc_hd__clkinv_2 _563_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d ));
 sky130_fd_sc_hd__clkinv_2 _564_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d ));
 sky130_fd_sc_hd__clkinv_2 _565_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d ));
 sky130_fd_sc_hd__clkinv_2 _566_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d ));
 sky130_fd_sc_hd__clkinv_2 _567_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d ));
 sky130_fd_sc_hd__clkinv_2 _568_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock ));
 sky130_fd_sc_hd__clkinv_2 _569_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d ));
 sky130_fd_sc_hd__clkinv_2 _570_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d ));
 sky130_fd_sc_hd__clkinv_2 _571_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d ));
 sky130_fd_sc_hd__clkinv_2 _572_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d ));
 sky130_fd_sc_hd__inv_2 _573_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d ));
 sky130_fd_sc_hd__clkinv_2 _574_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d ));
 sky130_fd_sc_hd__clkinv_2 _575_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d ));
 sky130_fd_sc_hd__clkinv_2 _576_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d ));
 sky130_fd_sc_hd__clkinv_2 _577_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d ));
 sky130_fd_sc_hd__clkinv_2 _578_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d ));
 sky130_fd_sc_hd__clkinv_2 _579_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d ));
 sky130_fd_sc_hd__clkinv_2 _580_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock ));
 sky130_fd_sc_hd__clkinv_2 _581_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d ));
 sky130_fd_sc_hd__clkinv_2 _582_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d ));
 sky130_fd_sc_hd__clkinv_2 _583_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d ));
 sky130_fd_sc_hd__clkinv_2 _584_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d ));
 sky130_fd_sc_hd__clkinv_2 _585_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d ));
 sky130_fd_sc_hd__inv_2 _586_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d ));
 sky130_fd_sc_hd__clkinv_2 _587_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d ));
 sky130_fd_sc_hd__clkinv_2 _588_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d ));
 sky130_fd_sc_hd__clkinv_2 _589_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d ));
 sky130_fd_sc_hd__clkinv_2 _590_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d ));
 sky130_fd_sc_hd__clkinv_2 _591_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d ));
 sky130_fd_sc_hd__clkinv_2 _592_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .Y(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock ));
 sky130_fd_sc_hd__inv_2 _593_ (.A(\CIRCUIT_2223.MEMORY_26.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_18.clock ));
 sky130_fd_sc_hd__clkinv_2 _594_ (.A(\CIRCUIT_2223.MEMORY_25.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_25.d ));
 sky130_fd_sc_hd__clkinv_2 _595_ (.A(net17),
    .Y(\CIRCUIT_2223.MEMORY_24.d ));
 sky130_fd_sc_hd__clkinv_2 _596_ (.A(\CIRCUIT_2223.MEMORY_22.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_22.d ));
 sky130_fd_sc_hd__clkinv_2 _597_ (.A(\CIRCUIT_2223.MEMORY_21.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_21.d ));
 sky130_fd_sc_hd__clkinv_2 _598_ (.A(\CIRCUIT_2223.MEMORY_20.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_20.d ));
 sky130_fd_sc_hd__clkinv_2 _599_ (.A(\CIRCUIT_2223.MEMORY_19.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_19.d ));
 sky130_fd_sc_hd__clkinv_2 _600_ (.A(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .Y(\CIRCUIT_2223.MEMORY_18.d ));
 sky130_fd_sc_hd__and4_1 _601_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[0] ),
    .X(_283_));
 sky130_fd_sc_hd__a22o_1 _602_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[1] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .X(_284_));
 sky130_fd_sc_hd__nand4_1 _603_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[1] ),
    .Y(_285_));
 sky130_fd_sc_hd__nand2_1 _604_ (.A(_284_),
    .B(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__xnor2_1 _605_ (.A(_283_),
    .B(_286_),
    .Y(net9));
 sky130_fd_sc_hd__and4_1 _606_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[2] ),
    .X(_287_));
 sky130_fd_sc_hd__a22oi_1 _607_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[2] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .Y(_288_));
 sky130_fd_sc_hd__or2_1 _608_ (.A(_287_),
    .B(_288_),
    .X(_289_));
 sky130_fd_sc_hd__a21bo_1 _609_ (.A1(_283_),
    .A2(_284_),
    .B1_N(_285_),
    .X(_290_));
 sky130_fd_sc_hd__xnor2_1 _610_ (.A(_289_),
    .B(_290_),
    .Y(net10));
 sky130_fd_sc_hd__and4_1 _611_ (.A(\CIRCUIT_2223.s_logisimNet48 ),
    .B(\CIRCUIT_2223.GATES_5.input2 ),
    .C(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ),
    .D(\CIRCUIT_2223.GATES_4.input1[3] ),
    .X(_291_));
 sky130_fd_sc_hd__a22o_1 _612_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[3] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .X(_292_));
 sky130_fd_sc_hd__and2b_1 _613_ (.A_N(_291_),
    .B(_292_),
    .X(_293_));
 sky130_fd_sc_hd__and2b_1 _614_ (.A_N(_289_),
    .B(_290_),
    .X(_294_));
 sky130_fd_sc_hd__nor2_1 _615_ (.A(_287_),
    .B(_294_),
    .Y(_295_));
 sky130_fd_sc_hd__xnor2_1 _616_ (.A(_293_),
    .B(_295_),
    .Y(net11));
 sky130_fd_sc_hd__a22oi_1 _617_ (.A1(\CIRCUIT_2223.GATES_3.input2 ),
    .A2(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ),
    .B1(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ),
    .B2(\CIRCUIT_2223.GATES_2.input2 ),
    .Y(_296_));
 sky130_fd_sc_hd__and4_1 _618_ (.A(\CIRCUIT_2223.GATES_3.input2 ),
    .B(\CIRCUIT_2223.GATES_2.input2 ),
    .C(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ),
    .X(_297_));
 sky130_fd_sc_hd__nor2_1 _619_ (.A(_296_),
    .B(_297_),
    .Y(_298_));
 sky130_fd_sc_hd__o31a_1 _620_ (.A1(_287_),
    .A2(_294_),
    .A3(_291_),
    .B1(_292_),
    .X(_299_));
 sky130_fd_sc_hd__xor2_1 _621_ (.A(_298_),
    .B(_299_),
    .X(net12));
 sky130_fd_sc_hd__a21o_1 _622_ (.A1(_298_),
    .A2(_299_),
    .B1(_297_),
    .X(net13));
 sky130_fd_sc_hd__a22oi_1 _623_ (.A1(\CIRCUIT_2223.GATES_5.input2 ),
    .A2(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .B1(\CIRCUIT_2223.GATES_4.input1[0] ),
    .B2(\CIRCUIT_2223.s_logisimNet48 ),
    .Y(_300_));
 sky130_fd_sc_hd__nor2_1 _624_ (.A(_283_),
    .B(_300_),
    .Y(net8));
 sky130_fd_sc_hd__xor2_1 _625_ (.A(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState ),
    .X(\CIRCUIT_2223.tone_generator_1.GATES_1.result ));
 sky130_fd_sc_hd__xor2_1 _626_ (.A(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState ),
    .X(\CIRCUIT_2223.tone_generator_1.GATES_2.result ));
 sky130_fd_sc_hd__xor2_1 _627_ (.A(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .B(\CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState ),
    .X(\CIRCUIT_2223.tone_generator_1.GATES_3.result ));
 sky130_fd_sc_hd__nor2_1 _628_ (.A(_243_),
    .B(_256_),
    .Y(\CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result ));
 sky130_fd_sc_hd__and4_2 _629_ (.A(net2),
    .B(net1),
    .C(\CIRCUIT_2223.GATES_1.input1[0] ),
    .D(_257_),
    .X(_301_));
 sky130_fd_sc_hd__nand2_1 _630_ (.A(_259_),
    .B(_301_),
    .Y(_302_));
 sky130_fd_sc_hd__mux2_1 _631_ (.A0(_188_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ),
    .S(_302_),
    .X(_303_));
 sky130_fd_sc_hd__clkbuf_1 _632_ (.A(_303_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _633_ (.A0(_186_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ),
    .S(_302_),
    .X(_304_));
 sky130_fd_sc_hd__clkbuf_1 _634_ (.A(_304_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _635_ (.A0(_184_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ),
    .S(_302_),
    .X(_305_));
 sky130_fd_sc_hd__clkbuf_1 _636_ (.A(_305_),
    .X(_121_));
 sky130_fd_sc_hd__buf_2 _637_ (.A(net7),
    .X(_306_));
 sky130_fd_sc_hd__nor2_1 _638_ (.A(\slow_clock[0] ),
    .B(_306_),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _639_ (.A1(\slow_clock[0] ),
    .A2(\slow_clock[1] ),
    .B1(_306_),
    .Y(_307_));
 sky130_fd_sc_hd__o21a_1 _640_ (.A1(\slow_clock[0] ),
    .A2(\slow_clock[1] ),
    .B1(_307_),
    .X(_123_));
 sky130_fd_sc_hd__a21oi_1 _641_ (.A1(\slow_clock[0] ),
    .A2(\slow_clock[1] ),
    .B1(\slow_clock[2] ),
    .Y(_308_));
 sky130_fd_sc_hd__and3_1 _642_ (.A(\slow_clock[0] ),
    .B(\slow_clock[1] ),
    .C(\slow_clock[2] ),
    .X(_309_));
 sky130_fd_sc_hd__nor3_1 _643_ (.A(_306_),
    .B(_308_),
    .C(_309_),
    .Y(_124_));
 sky130_fd_sc_hd__and4_1 _644_ (.A(\slow_clock[0] ),
    .B(\slow_clock[1] ),
    .C(\slow_clock[2] ),
    .D(\slow_clock[3] ),
    .X(_310_));
 sky130_fd_sc_hd__nor2_1 _645_ (.A(_306_),
    .B(_310_),
    .Y(_311_));
 sky130_fd_sc_hd__o21a_1 _646_ (.A1(\slow_clock[3] ),
    .A2(_309_),
    .B1(_311_),
    .X(_125_));
 sky130_fd_sc_hd__and2_1 _647_ (.A(\slow_clock[4] ),
    .B(_310_),
    .X(_312_));
 sky130_fd_sc_hd__nor2_1 _648_ (.A(_306_),
    .B(_312_),
    .Y(_313_));
 sky130_fd_sc_hd__o21a_1 _649_ (.A1(\slow_clock[4] ),
    .A2(_310_),
    .B1(_313_),
    .X(_126_));
 sky130_fd_sc_hd__and3_1 _650_ (.A(\slow_clock[4] ),
    .B(\slow_clock[5] ),
    .C(_310_),
    .X(_314_));
 sky130_fd_sc_hd__nor2_1 _651_ (.A(_306_),
    .B(_314_),
    .Y(_315_));
 sky130_fd_sc_hd__o21a_1 _652_ (.A1(\slow_clock[5] ),
    .A2(_312_),
    .B1(_315_),
    .X(_127_));
 sky130_fd_sc_hd__and2_1 _653_ (.A(\slow_clock[6] ),
    .B(_314_),
    .X(_316_));
 sky130_fd_sc_hd__nor2_1 _654_ (.A(_306_),
    .B(_316_),
    .Y(_317_));
 sky130_fd_sc_hd__o21a_1 _655_ (.A1(\slow_clock[6] ),
    .A2(_314_),
    .B1(_317_),
    .X(_128_));
 sky130_fd_sc_hd__a21oi_1 _656_ (.A1(net18),
    .A2(_316_),
    .B1(_306_),
    .Y(_318_));
 sky130_fd_sc_hd__o21a_1 _657_ (.A1(net18),
    .A2(_316_),
    .B1(_318_),
    .X(_129_));
 sky130_fd_sc_hd__buf_2 _658_ (.A(net7),
    .X(_319_));
 sky130_fd_sc_hd__nand2_1 _659_ (.A(_179_),
    .B(_319_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _660_ (.A(_179_),
    .B(_319_),
    .Y(_002_));
 sky130_fd_sc_hd__buf_2 _661_ (.A(net20),
    .X(_320_));
 sky130_fd_sc_hd__nand2_1 _662_ (.A(_320_),
    .B(_319_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _663_ (.A(_320_),
    .B(_319_),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_1 _664_ (.A(_320_),
    .B(_319_),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _665_ (.A(_320_),
    .B(_319_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _666_ (.A(_320_),
    .B(_319_),
    .Y(_007_));
 sky130_fd_sc_hd__nand2_1 _667_ (.A(_320_),
    .B(_319_),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_2 _668_ (.A(_180_),
    .B(_259_),
    .Y(_321_));
 sky130_fd_sc_hd__mux2_1 _669_ (.A0(_188_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ),
    .S(_321_),
    .X(_322_));
 sky130_fd_sc_hd__clkbuf_1 _670_ (.A(_322_),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _671_ (.A0(_186_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ),
    .S(_321_),
    .X(_323_));
 sky130_fd_sc_hd__clkbuf_1 _672_ (.A(_323_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _673_ (.A0(_184_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ),
    .S(_321_),
    .X(_324_));
 sky130_fd_sc_hd__clkbuf_1 _674_ (.A(_324_),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _675_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ),
    .S(_321_),
    .X(_325_));
 sky130_fd_sc_hd__clkbuf_1 _676_ (.A(_325_),
    .X(_133_));
 sky130_fd_sc_hd__and4b_2 _677_ (.A_N(\CIRCUIT_2223.GATES_1.input1[0] ),
    .B(\CIRCUIT_2223.GATES_1.input1[1] ),
    .C(net2),
    .D(net1),
    .X(_326_));
 sky130_fd_sc_hd__nand2_1 _678_ (.A(_259_),
    .B(_326_),
    .Y(_327_));
 sky130_fd_sc_hd__mux2_1 _679_ (.A0(_188_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ),
    .S(_327_),
    .X(_328_));
 sky130_fd_sc_hd__clkbuf_1 _680_ (.A(_328_),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _681_ (.A0(_186_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ),
    .S(_327_),
    .X(_329_));
 sky130_fd_sc_hd__clkbuf_1 _682_ (.A(_329_),
    .X(_135_));
 sky130_fd_sc_hd__mux2_1 _683_ (.A0(_184_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ),
    .S(_327_),
    .X(_330_));
 sky130_fd_sc_hd__clkbuf_1 _684_ (.A(_330_),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _685_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ),
    .S(_327_),
    .X(_331_));
 sky130_fd_sc_hd__clkbuf_1 _686_ (.A(_331_),
    .X(_137_));
 sky130_fd_sc_hd__or2b_1 _687_ (.A(net1),
    .B_N(net2),
    .X(_332_));
 sky130_fd_sc_hd__mux2_1 _688_ (.A0(_188_),
    .A1(\CIRCUIT_2223.GATES_1.input1[0] ),
    .S(_332_),
    .X(_333_));
 sky130_fd_sc_hd__clkbuf_1 _689_ (.A(_333_),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _690_ (.A0(_186_),
    .A1(\CIRCUIT_2223.GATES_1.input1[1] ),
    .S(_332_),
    .X(_334_));
 sky130_fd_sc_hd__clkbuf_1 _691_ (.A(_334_),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _692_ (.A0(_184_),
    .A1(\CIRCUIT_2223.GATES_1.input1[2] ),
    .S(_332_),
    .X(_335_));
 sky130_fd_sc_hd__clkbuf_1 _693_ (.A(_335_),
    .X(_140_));
 sky130_fd_sc_hd__mux2_1 _694_ (.A0(net6),
    .A1(\CIRCUIT_2223.GATES_1.input1[3] ),
    .S(_332_),
    .X(_336_));
 sky130_fd_sc_hd__clkbuf_1 _695_ (.A(_336_),
    .X(_141_));
 sky130_fd_sc_hd__clkinv_2 _696_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(_010_));
 sky130_fd_sc_hd__clkinv_2 _697_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(_012_));
 sky130_fd_sc_hd__clkinv_2 _698_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(_014_));
 sky130_fd_sc_hd__clkinv_2 _699_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(_016_));
 sky130_fd_sc_hd__clkinv_2 _700_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _701_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(_020_));
 sky130_fd_sc_hd__xor2_2 _702_ (.A(_215_),
    .B(clknet_1_0__leaf__281_),
    .X(_021_));
 sky130_fd_sc_hd__clkinv_2 _703_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(_023_));
 sky130_fd_sc_hd__clkinv_2 _704_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(_025_));
 sky130_fd_sc_hd__clkinv_2 _705_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(_027_));
 sky130_fd_sc_hd__clkinv_2 _706_ (.A(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(_029_));
 sky130_fd_sc_hd__clkinv_2 _707_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ),
    .Y(_031_));
 sky130_fd_sc_hd__clkinv_2 _708_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ),
    .Y(_033_));
 sky130_fd_sc_hd__clkinv_2 _709_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ),
    .Y(_035_));
 sky130_fd_sc_hd__clkinv_2 _710_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_2 _711_ (.A(_191_),
    .B(clknet_1_1__leaf__262_),
    .Y(_038_));
 sky130_fd_sc_hd__clkinv_2 _712_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ),
    .Y(_040_));
 sky130_fd_sc_hd__clkinv_2 _713_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ),
    .Y(_042_));
 sky130_fd_sc_hd__clkinv_2 _714_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ),
    .Y(_044_));
 sky130_fd_sc_hd__clkinv_2 _715_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ),
    .Y(_046_));
 sky130_fd_sc_hd__clkinv_2 _716_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ),
    .Y(_048_));
 sky130_fd_sc_hd__clkinv_2 _717_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ),
    .Y(_050_));
 sky130_fd_sc_hd__clkinv_2 _718_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ),
    .Y(_051_));
 sky130_fd_sc_hd__clkinv_2 _719_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ),
    .Y(_052_));
 sky130_fd_sc_hd__clkinv_2 _720_ (.A(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ),
    .Y(_053_));
 sky130_fd_sc_hd__nand2_1 _721_ (.A(_180_),
    .B(_192_),
    .Y(_337_));
 sky130_fd_sc_hd__mux2_1 _722_ (.A0(_188_),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ),
    .S(_337_),
    .X(_338_));
 sky130_fd_sc_hd__clkbuf_1 _723_ (.A(_338_),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _724_ (.A0(_186_),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ),
    .S(_337_),
    .X(_339_));
 sky130_fd_sc_hd__clkbuf_1 _725_ (.A(_339_),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _726_ (.A0(_184_),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ),
    .S(_337_),
    .X(_340_));
 sky130_fd_sc_hd__clkbuf_1 _727_ (.A(_340_),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _728_ (.A0(_188_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ),
    .S(_260_),
    .X(_341_));
 sky130_fd_sc_hd__clkbuf_1 _729_ (.A(_341_),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _730_ (.A0(_186_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ),
    .S(_260_),
    .X(_342_));
 sky130_fd_sc_hd__clkbuf_1 _731_ (.A(_342_),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _732_ (.A0(_184_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ),
    .S(_260_),
    .X(_343_));
 sky130_fd_sc_hd__clkbuf_1 _733_ (.A(_343_),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _734_ (.A0(net6),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ),
    .S(_260_),
    .X(_344_));
 sky130_fd_sc_hd__clkbuf_1 _735_ (.A(_344_),
    .X(_148_));
 sky130_fd_sc_hd__nand2_1 _736_ (.A(_193_),
    .B(_259_),
    .Y(_345_));
 sky130_fd_sc_hd__mux2_1 _737_ (.A0(_188_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ),
    .S(_345_),
    .X(_346_));
 sky130_fd_sc_hd__clkbuf_1 _738_ (.A(_346_),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _739_ (.A0(_186_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ),
    .S(_345_),
    .X(_347_));
 sky130_fd_sc_hd__clkbuf_1 _740_ (.A(_347_),
    .X(_150_));
 sky130_fd_sc_hd__mux2_1 _741_ (.A0(_184_),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ),
    .S(_345_),
    .X(_348_));
 sky130_fd_sc_hd__clkbuf_1 _742_ (.A(_348_),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _743_ (.A0(net6),
    .A1(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ),
    .S(_345_),
    .X(_349_));
 sky130_fd_sc_hd__clkbuf_1 _744_ (.A(_349_),
    .X(_152_));
 sky130_fd_sc_hd__inv_2 _745_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ),
    .Y(_055_));
 sky130_fd_sc_hd__clkinv_2 _746_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ),
    .Y(_057_));
 sky130_fd_sc_hd__clkinv_2 _747_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ),
    .Y(_059_));
 sky130_fd_sc_hd__clkinv_2 _748_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ),
    .Y(_061_));
 sky130_fd_sc_hd__xnor2_2 _749_ (.A(_191_),
    .B(clknet_1_1__leaf__235_),
    .Y(_062_));
 sky130_fd_sc_hd__clkinv_2 _750_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ),
    .Y(_064_));
 sky130_fd_sc_hd__clkinv_2 _751_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ),
    .Y(_066_));
 sky130_fd_sc_hd__clkinv_2 _752_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ),
    .Y(_068_));
 sky130_fd_sc_hd__clkinv_2 _753_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ),
    .Y(_070_));
 sky130_fd_sc_hd__clkinv_2 _754_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ),
    .Y(_072_));
 sky130_fd_sc_hd__clkinv_2 _755_ (.A(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_1 _756_ (.A(_181_),
    .B(_193_),
    .Y(_350_));
 sky130_fd_sc_hd__mux2_1 _757_ (.A0(_188_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ),
    .S(_350_),
    .X(_351_));
 sky130_fd_sc_hd__clkbuf_1 _758_ (.A(_351_),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _759_ (.A0(_186_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ),
    .S(_350_),
    .X(_352_));
 sky130_fd_sc_hd__clkbuf_1 _760_ (.A(_352_),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _761_ (.A0(_184_),
    .A1(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ),
    .S(_350_),
    .X(_353_));
 sky130_fd_sc_hd__clkbuf_1 _762_ (.A(_353_),
    .X(_155_));
 sky130_fd_sc_hd__nand2_2 _763_ (.A(_193_),
    .B(_233_),
    .Y(_354_));
 sky130_fd_sc_hd__mux2_1 _764_ (.A0(_188_),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ),
    .S(_354_),
    .X(_355_));
 sky130_fd_sc_hd__clkbuf_1 _765_ (.A(_355_),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _766_ (.A0(_186_),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ),
    .S(_354_),
    .X(_356_));
 sky130_fd_sc_hd__clkbuf_1 _767_ (.A(_356_),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _768_ (.A0(_184_),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ),
    .S(_354_),
    .X(_357_));
 sky130_fd_sc_hd__clkbuf_1 _769_ (.A(_357_),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _770_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ),
    .S(_354_),
    .X(_358_));
 sky130_fd_sc_hd__clkbuf_1 _771_ (.A(_358_),
    .X(_159_));
 sky130_fd_sc_hd__nand2_2 _772_ (.A(_233_),
    .B(_301_),
    .Y(_359_));
 sky130_fd_sc_hd__mux2_1 _773_ (.A0(net3),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ),
    .S(_359_),
    .X(_360_));
 sky130_fd_sc_hd__clkbuf_1 _774_ (.A(_360_),
    .X(_160_));
 sky130_fd_sc_hd__mux2_1 _775_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ),
    .S(_359_),
    .X(_361_));
 sky130_fd_sc_hd__clkbuf_1 _776_ (.A(_361_),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _777_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ),
    .S(_359_),
    .X(_362_));
 sky130_fd_sc_hd__clkbuf_1 _778_ (.A(_362_),
    .X(_162_));
 sky130_fd_sc_hd__mux2_1 _779_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ),
    .S(_359_),
    .X(_363_));
 sky130_fd_sc_hd__clkbuf_1 _780_ (.A(_363_),
    .X(_163_));
 sky130_fd_sc_hd__clkinv_2 _781_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ),
    .Y(_076_));
 sky130_fd_sc_hd__clkinv_2 _782_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ),
    .Y(_078_));
 sky130_fd_sc_hd__clkinv_2 _783_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ),
    .Y(_080_));
 sky130_fd_sc_hd__clkinv_2 _784_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ),
    .Y(_082_));
 sky130_fd_sc_hd__xor2_2 _785_ (.A(_215_),
    .B(clknet_1_0__leaf__212_),
    .X(_083_));
 sky130_fd_sc_hd__inv_2 _786_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _787_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ),
    .Y(_087_));
 sky130_fd_sc_hd__clkinv_2 _788_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ),
    .Y(_089_));
 sky130_fd_sc_hd__clkinv_2 _789_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ),
    .Y(_091_));
 sky130_fd_sc_hd__clkinv_2 _790_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ),
    .Y(_093_));
 sky130_fd_sc_hd__clkinv_2 _791_ (.A(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ),
    .Y(_095_));
 sky130_fd_sc_hd__nand2_1 _792_ (.A(_233_),
    .B(_326_),
    .Y(_364_));
 sky130_fd_sc_hd__mux2_1 _793_ (.A0(net3),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ),
    .S(_364_),
    .X(_365_));
 sky130_fd_sc_hd__clkbuf_1 _794_ (.A(_365_),
    .X(_164_));
 sky130_fd_sc_hd__mux2_1 _795_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ),
    .S(_364_),
    .X(_366_));
 sky130_fd_sc_hd__clkbuf_1 _796_ (.A(_366_),
    .X(_165_));
 sky130_fd_sc_hd__mux2_1 _797_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ),
    .S(_364_),
    .X(_367_));
 sky130_fd_sc_hd__clkbuf_1 _798_ (.A(_367_),
    .X(_166_));
 sky130_fd_sc_hd__nand2_1 _799_ (.A(_192_),
    .B(_301_),
    .Y(_368_));
 sky130_fd_sc_hd__mux2_1 _800_ (.A0(net3),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ),
    .S(_368_),
    .X(_369_));
 sky130_fd_sc_hd__clkbuf_1 _801_ (.A(_369_),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _802_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ),
    .S(_368_),
    .X(_370_));
 sky130_fd_sc_hd__clkbuf_1 _803_ (.A(_370_),
    .X(_168_));
 sky130_fd_sc_hd__mux2_1 _804_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ),
    .S(_368_),
    .X(_371_));
 sky130_fd_sc_hd__clkbuf_1 _805_ (.A(_371_),
    .X(_169_));
 sky130_fd_sc_hd__mux2_1 _806_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ),
    .S(_368_),
    .X(_372_));
 sky130_fd_sc_hd__clkbuf_1 _807_ (.A(_372_),
    .X(_170_));
 sky130_fd_sc_hd__nand2_2 _808_ (.A(_192_),
    .B(_326_),
    .Y(_373_));
 sky130_fd_sc_hd__mux2_1 _809_ (.A0(net3),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ),
    .S(_373_),
    .X(_374_));
 sky130_fd_sc_hd__clkbuf_1 _810_ (.A(_374_),
    .X(_171_));
 sky130_fd_sc_hd__mux2_1 _811_ (.A0(net4),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ),
    .S(_373_),
    .X(_375_));
 sky130_fd_sc_hd__clkbuf_1 _812_ (.A(_375_),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _813_ (.A0(net5),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ),
    .S(_373_),
    .X(_376_));
 sky130_fd_sc_hd__clkbuf_1 _814_ (.A(_376_),
    .X(_173_));
 sky130_fd_sc_hd__mux2_1 _815_ (.A0(net6),
    .A1(\CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ),
    .S(_373_),
    .X(_377_));
 sky130_fd_sc_hd__clkbuf_1 _816_ (.A(_377_),
    .X(_174_));
 sky130_fd_sc_hd__and2_1 _817_ (.A(_181_),
    .B(_326_),
    .X(_378_));
 sky130_fd_sc_hd__clkbuf_1 _818_ (.A(_378_),
    .X(_096_));
 sky130_fd_sc_hd__and2_1 _819_ (.A(_181_),
    .B(_301_),
    .X(_379_));
 sky130_fd_sc_hd__clkbuf_1 _820_ (.A(_379_),
    .X(_097_));
 sky130_fd_sc_hd__nand2_1 _821_ (.A(_320_),
    .B(_319_),
    .Y(_098_));
 sky130_fd_sc_hd__nand2_1 _822_ (.A(_320_),
    .B(_319_),
    .Y(_099_));
 sky130_fd_sc_hd__nand2_1 _823_ (.A(_320_),
    .B(_306_),
    .Y(_100_));
 sky130_fd_sc_hd__nand2_1 _824_ (.A(_320_),
    .B(_306_),
    .Y(_101_));
 sky130_fd_sc_hd__clkinv_2 _825_ (.A(\CIRCUIT_2223.MEMORY_25.s_currentState ),
    .Y(_103_));
 sky130_fd_sc_hd__clkinv_2 _826_ (.A(net17),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _827_ (.A(_179_),
    .Y(_106_));
 sky130_fd_sc_hd__clkinv_2 _828_ (.A(\CIRCUIT_2223.MEMORY_22.s_currentState ),
    .Y(_108_));
 sky130_fd_sc_hd__clkinv_2 _829_ (.A(\CIRCUIT_2223.MEMORY_21.s_currentState ),
    .Y(_110_));
 sky130_fd_sc_hd__clkinv_2 _830_ (.A(\CIRCUIT_2223.MEMORY_20.s_currentState ),
    .Y(_112_));
 sky130_fd_sc_hd__clkinv_2 _831_ (.A(\CIRCUIT_2223.MEMORY_19.s_currentState ),
    .Y(_114_));
 sky130_fd_sc_hd__clkinv_2 _832_ (.A(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .Y(_116_));
 sky130_fd_sc_hd__clkinv_2 _833_ (.A(\CIRCUIT_2223.MEMORY_26.s_currentState ),
    .Y(_118_));
 sky130_fd_sc_hd__dfxtp_1 _834_ (.CLK(net22),
    .D(_119_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _835_ (.CLK(net22),
    .D(_120_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _836_ (.CLK(net23),
    .D(_121_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _837_ (.CLK(clknet_1_0__leaf_clk),
    .D(_122_),
    .Q(\slow_clock[0] ));
 sky130_fd_sc_hd__dfxtp_1 _838_ (.CLK(clknet_1_0__leaf_clk),
    .D(_123_),
    .Q(\slow_clock[1] ));
 sky130_fd_sc_hd__dfxtp_1 _839_ (.CLK(clknet_1_0__leaf_clk),
    .D(_124_),
    .Q(\slow_clock[2] ));
 sky130_fd_sc_hd__dfxtp_1 _840_ (.CLK(clknet_1_0__leaf_clk),
    .D(_125_),
    .Q(\slow_clock[3] ));
 sky130_fd_sc_hd__dfxtp_1 _841_ (.CLK(clknet_1_0__leaf_clk),
    .D(_126_),
    .Q(\slow_clock[4] ));
 sky130_fd_sc_hd__dfxtp_1 _842_ (.CLK(clknet_1_0__leaf_clk),
    .D(_127_),
    .Q(\slow_clock[5] ));
 sky130_fd_sc_hd__dfxtp_1 _843_ (.CLK(clknet_1_1__leaf_clk),
    .D(_128_),
    .Q(\slow_clock[6] ));
 sky130_fd_sc_hd__dfxtp_1 _844_ (.CLK(clknet_1_1__leaf_clk),
    .D(_129_),
    .Q(\CIRCUIT_2223.CLK ));
 sky130_fd_sc_hd__dfxtp_1 _845_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _846_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _847_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _848_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _849_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ),
    .Q(\CIRCUIT_2223.GATES_4.input1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _850_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _851_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.GATES_1.result ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _852_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.GATES_2.result ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _853_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _854_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.GATES_3.result ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _855_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState ),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _856_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState ),
    .SET_B(_000_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _857_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState ),
    .RESET_B(_001_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _858_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState ),
    .SET_B(_002_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _859_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState ),
    .RESET_B(_003_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _860_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState ),
    .SET_B(_004_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _861_ (.CLK(net17),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState ),
    .RESET_B(_005_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _862_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState ),
    .SET_B(_006_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState ));
 sky130_fd_sc_hd__dfstp_1 _863_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState ),
    .SET_B(_007_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _864_ (.CLK(net16),
    .D(\CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState ),
    .RESET_B(_008_),
    .Q(\CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _865_ (.CLK(net22),
    .D(_130_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _866_ (.CLK(net25),
    .D(_131_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _867_ (.CLK(net24),
    .D(_132_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _868_ (.CLK(net24),
    .D(_133_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _869_ (.CLK(net23),
    .D(_134_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _870_ (.CLK(net22),
    .D(_135_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _871_ (.CLK(net22),
    .D(_136_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _872_ (.CLK(net22),
    .D(_137_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _873_ (.CLK(net19),
    .D(_138_),
    .Q(\CIRCUIT_2223.GATES_1.input1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _874_ (.CLK(net20),
    .D(_139_),
    .Q(\CIRCUIT_2223.GATES_1.input1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _875_ (.CLK(net20),
    .D(_140_),
    .Q(\CIRCUIT_2223.GATES_1.input1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _876_ (.CLK(net20),
    .D(_141_),
    .Q(\CIRCUIT_2223.GATES_1.input1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _877_ (.CLK(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result ),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _878_ (.CLK(_010_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock ),
    .RESET_B(_009_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _879_ (.CLK(_012_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d ),
    .RESET_B(_011_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _880_ (.CLK(_014_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d ),
    .RESET_B(_013_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _881_ (.CLK(_016_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d ),
    .RESET_B(_015_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _882_ (.CLK(_018_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d ),
    .RESET_B(_017_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _883_ (.CLK(_020_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d ),
    .RESET_B(_019_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _884_ (.CLK(\CIRCUIT_2223.MEMORY_24.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d ),
    .RESET_B(_021_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _885_ (.CLK(_023_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d ),
    .RESET_B(_022_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _886_ (.CLK(_025_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d ),
    .RESET_B(_024_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _887_ (.CLK(_027_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d ),
    .RESET_B(_026_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _888_ (.CLK(_029_),
    .D(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d ),
    .RESET_B(_028_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _889_ (.CLK(_031_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d ),
    .RESET_B(_030_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _890_ (.CLK(_033_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d ),
    .RESET_B(_032_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _891_ (.CLK(_035_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d ),
    .RESET_B(_034_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _892_ (.CLK(_037_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d ),
    .RESET_B(_036_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _893_ (.CLK(\CIRCUIT_2223.MEMORY_24.s_currentState ),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d ),
    .RESET_B(_038_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _894_ (.CLK(_040_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d ),
    .RESET_B(_039_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _895_ (.CLK(_042_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d ),
    .RESET_B(_041_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _896_ (.CLK(_044_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d ),
    .RESET_B(_043_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _897_ (.CLK(_046_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d ),
    .RESET_B(_045_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _898_ (.CLK(_048_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d ),
    .RESET_B(_047_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _899_ (.CLK(_050_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock ),
    .RESET_B(_049_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _900_ (.CLK(\CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result ),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _901_ (.CLK(_051_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _902_ (.CLK(_052_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _903_ (.CLK(_053_),
    .D(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock ),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _904_ (.CLK(net24),
    .D(_142_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _905_ (.CLK(net25),
    .D(_143_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _906_ (.CLK(net25),
    .D(_144_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _907_ (.CLK(net23),
    .D(_145_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _908_ (.CLK(net23),
    .D(_146_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _909_ (.CLK(net23),
    .D(_147_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _910_ (.CLK(net23),
    .D(_148_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _911_ (.CLK(net22),
    .D(_149_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _912_ (.CLK(net22),
    .D(_150_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _913_ (.CLK(net22),
    .D(_151_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _914_ (.CLK(net22),
    .D(_152_),
    .Q(\CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 ));
 sky130_fd_sc_hd__dfrtp_1 _915_ (.CLK(_055_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d ),
    .RESET_B(_054_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _916_ (.CLK(_057_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d ),
    .RESET_B(_056_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _917_ (.CLK(_059_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d ),
    .RESET_B(_058_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _918_ (.CLK(_061_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d ),
    .RESET_B(_060_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _919_ (.CLK(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d ),
    .RESET_B(_062_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _920_ (.CLK(_064_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d ),
    .RESET_B(_063_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _921_ (.CLK(_066_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d ),
    .RESET_B(_065_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _922_ (.CLK(_068_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d ),
    .RESET_B(_067_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _923_ (.CLK(_070_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d ),
    .RESET_B(_069_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _924_ (.CLK(_072_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d ),
    .RESET_B(_071_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _925_ (.CLK(_074_),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock ),
    .RESET_B(_073_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _926_ (.CLK(\CIRCUIT_2223.tone_generator_2_1.GATES_27.result ),
    .D(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _927_ (.CLK(net24),
    .D(_153_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _928_ (.CLK(net25),
    .D(_154_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _929_ (.CLK(net25),
    .D(_155_),
    .Q(\CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _930_ (.CLK(net19),
    .D(_156_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _931_ (.CLK(net19),
    .D(_157_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _932_ (.CLK(net19),
    .D(_158_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _933_ (.CLK(net19),
    .D(_159_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _934_ (.CLK(net18),
    .D(_160_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _935_ (.CLK(net18),
    .D(_161_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _936_ (.CLK(net18),
    .D(_162_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _937_ (.CLK(net18),
    .D(_163_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 ));
 sky130_fd_sc_hd__dfrtp_1 _938_ (.CLK(_076_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d ),
    .RESET_B(_075_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _939_ (.CLK(_078_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d ),
    .RESET_B(_077_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _940_ (.CLK(_080_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d ),
    .RESET_B(_079_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _941_ (.CLK(_082_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d ),
    .RESET_B(_081_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _942_ (.CLK(\CIRCUIT_2223.MEMORY_18.s_currentState ),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d ),
    .RESET_B(_083_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _943_ (.CLK(_085_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d ),
    .RESET_B(_084_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _944_ (.CLK(_087_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d ),
    .RESET_B(_086_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _945_ (.CLK(_089_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d ),
    .RESET_B(_088_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _946_ (.CLK(_091_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d ),
    .RESET_B(_090_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _947_ (.CLK(_093_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d ),
    .RESET_B(_092_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _948_ (.CLK(_095_),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock ),
    .RESET_B(_094_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _949_ (.CLK(\CIRCUIT_2223.tone_generator_2_2.GATES_27.result ),
    .D(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d ),
    .Q(\CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _950_ (.CLK(net18),
    .D(_164_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _951_ (.CLK(net18),
    .D(_165_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _952_ (.CLK(net19),
    .D(_166_),
    .Q(\CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _953_ (.CLK(net21),
    .D(_167_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _954_ (.CLK(net20),
    .D(_168_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _955_ (.CLK(net21),
    .D(_169_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _956_ (.CLK(net21),
    .D(_170_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _957_ (.CLK(net24),
    .D(_171_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _958_ (.CLK(net24),
    .D(_172_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _959_ (.CLK(net24),
    .D(_173_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _960_ (.CLK(net24),
    .D(_174_),
    .Q(\CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 ));
 sky130_fd_sc_hd__dfxtp_1 _961_ (.CLK(_096_),
    .D(net3),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _962_ (.CLK(_097_),
    .D(net3),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _963_ (.CLK(net20),
    .D(_175_),
    .RESET_B(_098_),
    .Q(\CIRCUIT_2223.GATES_2.input2 ));
 sky130_fd_sc_hd__dfrtp_1 _964_ (.CLK(net20),
    .D(_176_),
    .RESET_B(_099_),
    .Q(\CIRCUIT_2223.GATES_3.input2 ));
 sky130_fd_sc_hd__dfrtp_2 _965_ (.CLK(net20),
    .D(_177_),
    .RESET_B(_100_),
    .Q(\CIRCUIT_2223.GATES_5.input2 ));
 sky130_fd_sc_hd__dfrtp_2 _966_ (.CLK(net20),
    .D(_178_),
    .RESET_B(_101_),
    .Q(\CIRCUIT_2223.s_logisimNet48 ));
 sky130_fd_sc_hd__dfrtp_1 _967_ (.CLK(_103_),
    .D(\CIRCUIT_2223.MEMORY_18.clock ),
    .RESET_B(_102_),
    .Q(\CIRCUIT_2223.MEMORY_26.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _968_ (.CLK(_105_),
    .D(\CIRCUIT_2223.MEMORY_25.d ),
    .RESET_B(_104_),
    .Q(\CIRCUIT_2223.MEMORY_25.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _969_ (.CLK(net26),
    .D(\CIRCUIT_2223.MEMORY_24.d ),
    .RESET_B(_106_),
    .Q(\CIRCUIT_2223.MEMORY_24.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _970_ (.CLK(_108_),
    .D(\CIRCUIT_2223.GATES_11.input2 ),
    .RESET_B(_107_),
    .Q(\CIRCUIT_2223.MEMORY_23.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _971_ (.CLK(_110_),
    .D(\CIRCUIT_2223.MEMORY_22.d ),
    .RESET_B(_109_),
    .Q(\CIRCUIT_2223.MEMORY_22.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _972_ (.CLK(_112_),
    .D(\CIRCUIT_2223.MEMORY_21.d ),
    .RESET_B(_111_),
    .Q(\CIRCUIT_2223.MEMORY_21.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _973_ (.CLK(_114_),
    .D(\CIRCUIT_2223.MEMORY_20.d ),
    .RESET_B(_113_),
    .Q(\CIRCUIT_2223.MEMORY_20.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _974_ (.CLK(_116_),
    .D(\CIRCUIT_2223.MEMORY_19.d ),
    .RESET_B(_115_),
    .Q(\CIRCUIT_2223.MEMORY_19.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _975_ (.CLK(_118_),
    .D(\CIRCUIT_2223.MEMORY_18.d ),
    .RESET_B(_117_),
    .Q(\CIRCUIT_2223.MEMORY_18.s_currentState ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(rst),
    .X(net7));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(io_out[7]));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(\CIRCUIT_2223.MEMORY_24.s_currentState ),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(net21),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(net21),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(net28),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 fanout23 (.A(\CIRCUIT_2223.CLK ),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(\CIRCUIT_2223.CLK ),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout25 (.A(\CIRCUIT_2223.CLK ),
    .X(net25));
 sky130_fd_sc_hd__inv_2 _475__1 (.A(clknet_1_0__leaf__195_),
    .Y(net26));
 sky130_fd_sc_hd__inv_2 _475__2 (.A(clknet_1_1__leaf__195_),
    .Y(net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__195_ (.A(_195_),
    .X(clknet_0__195_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__195_ (.A(clknet_0__195_),
    .X(clknet_1_0__leaf__195_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__195_ (.A(clknet_0__195_),
    .X(clknet_1_1__leaf__195_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__262_ (.A(_262_),
    .X(clknet_0__262_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__262_ (.A(clknet_0__262_),
    .X(clknet_1_0__leaf__262_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__262_ (.A(clknet_0__262_),
    .X(clknet_1_1__leaf__262_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__263_ (.A(_263_),
    .X(clknet_0__263_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__263_ (.A(clknet_0__263_),
    .X(clknet_1_0__leaf__263_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__263_ (.A(clknet_0__263_),
    .X(clknet_1_1__leaf__263_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__281_ (.A(_281_),
    .X(clknet_0__281_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__281_ (.A(clknet_0__281_),
    .X(clknet_1_0__leaf__281_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__281_ (.A(clknet_0__281_),
    .X(clknet_1_1__leaf__281_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__282_ (.A(_282_),
    .X(clknet_0__282_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__282_ (.A(clknet_0__282_),
    .X(clknet_1_0__leaf__282_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__282_ (.A(clknet_0__282_),
    .X(clknet_1_1__leaf__282_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__235_ (.A(_235_),
    .X(clknet_0__235_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__235_ (.A(clknet_0__235_),
    .X(clknet_1_0__leaf__235_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__235_ (.A(clknet_0__235_),
    .X(clknet_1_1__leaf__235_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__236_ (.A(_236_),
    .X(clknet_0__236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__236_ (.A(clknet_0__236_),
    .X(clknet_1_0__leaf__236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__236_ (.A(clknet_0__236_),
    .X(clknet_1_1__leaf__236_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__212_ (.A(_212_),
    .X(clknet_0__212_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__212_ (.A(clknet_0__212_),
    .X(clknet_1_0__leaf__212_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__212_ (.A(clknet_0__212_),
    .X(clknet_1_1__leaf__212_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__213_ (.A(_213_),
    .X(clknet_0__213_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__213_ (.A(clknet_0__213_),
    .X(clknet_1_0__leaf__213_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__213_ (.A(clknet_0__213_),
    .X(clknet_1_1__leaf__213_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\CIRCUIT_2223.CLK ),
    .X(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1_A (.DIODE(\CIRCUIT_2223.CLK ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(\CIRCUIT_2223.CLK ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(\CIRCUIT_2223.CLK ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(\CIRCUIT_2223.CLK ));
 sky130_fd_sc_hd__diode_2 ANTENNA__856__SET_B (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__532__A (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__434__A (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__433__A (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__432__A (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__430__A (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__768__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__761__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__741__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__732__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__726__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__692__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__683__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__673__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__635__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__395__A0 (.DIODE(_184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__766__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__759__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__739__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__730__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__724__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__690__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__681__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__671__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__633__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__398__A0 (.DIODE(_186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__764__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__757__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__737__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__728__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__722__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__688__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__679__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__669__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__631__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__401__A0 (.DIODE(_188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__749__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__711__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__511__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__509__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__508__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__507__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__506__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__435__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__405__A (.DIODE(_191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__785__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__702__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__541__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__540__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__539__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__538__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__502__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__465__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__464__A (.DIODE(_215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__824__B (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__823__B (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__656__B1 (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__654__A (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__651__A (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__648__A (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__645__A (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__643__A (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__639__B1 (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__638__B (.DIODE(_306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__822__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__821__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__667__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__666__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__665__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__664__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__663__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__662__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__660__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__659__B (.DIODE(_319_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__687__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__677__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__629__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__459__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__407__C1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__406__C1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__389__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__962__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__961__D (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__809__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__800__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__793__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__773__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__400__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__811__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__802__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__795__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__775__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__397__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__813__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__804__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__797__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__777__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__394__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__815__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__806__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__779__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__770__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__743__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__734__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__694__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__685__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__675__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__392__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__956__CLK (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__953__CLK (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__955__CLK (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net21));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_287 ();
endmodule

