VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt2_tholin_diceroll
  CLASS BLOCK ;
  FOREIGN tt2_tholin_diceroll ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 106.000 18.770 110.000 ;
    END
  END clk
  PIN io_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 106.000 91.450 110.000 ;
    END
  END io_in
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_out[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 106.000 55.110 110.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.080 10.640 18.680 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.805 10.640 43.405 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.530 10.640 68.130 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.255 10.640 92.855 98.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 29.440 10.640 31.040 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.165 10.640 55.765 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.890 10.640 80.490 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.615 10.640 105.215 98.160 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 93.785 104.610 96.615 ;
        RECT 5.330 88.345 104.610 91.175 ;
        RECT 5.330 82.905 104.610 85.735 ;
        RECT 5.330 77.465 104.610 80.295 ;
        RECT 5.330 72.025 104.610 74.855 ;
        RECT 5.330 66.585 104.610 69.415 ;
        RECT 5.330 61.145 104.610 63.975 ;
        RECT 5.330 55.705 104.610 58.535 ;
        RECT 5.330 50.265 104.610 53.095 ;
        RECT 5.330 44.825 104.610 47.655 ;
        RECT 5.330 39.385 104.610 42.215 ;
        RECT 5.330 33.945 104.610 36.775 ;
        RECT 5.330 28.505 104.610 31.335 ;
        RECT 5.330 23.065 104.610 25.895 ;
        RECT 5.330 17.625 104.610 20.455 ;
        RECT 5.330 12.185 104.610 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 104.420 98.005 ;
      LAYER met1 ;
        RECT 5.520 10.640 105.215 98.560 ;
      LAYER met2 ;
        RECT 7.920 105.720 18.210 106.490 ;
        RECT 19.050 105.720 54.550 106.490 ;
        RECT 55.390 105.720 90.890 106.490 ;
        RECT 91.730 105.720 105.185 106.490 ;
        RECT 7.920 4.280 105.185 105.720 ;
        RECT 8.470 4.000 20.970 4.280 ;
        RECT 21.810 4.000 34.310 4.280 ;
        RECT 35.150 4.000 47.650 4.280 ;
        RECT 48.490 4.000 60.990 4.280 ;
        RECT 61.830 4.000 74.330 4.280 ;
        RECT 75.170 4.000 87.670 4.280 ;
        RECT 88.510 4.000 101.010 4.280 ;
        RECT 101.850 4.000 105.185 4.280 ;
      LAYER met3 ;
        RECT 17.090 10.715 105.205 98.085 ;
  END
END tt2_tholin_diceroll
END LIBRARY

