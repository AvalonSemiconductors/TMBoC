magic
tech sky130B
magscale 1 2
timestamp 1675976271
<< viali >>
rect 2145 19465 2179 19499
rect 1961 19329 1995 19363
rect 4905 16065 4939 16099
rect 4997 16065 5031 16099
rect 5089 16065 5123 16099
rect 5733 16065 5767 16099
rect 5917 16065 5951 16099
rect 6837 16065 6871 16099
rect 7021 16065 7055 16099
rect 4721 15861 4755 15895
rect 5825 15861 5859 15895
rect 7021 15861 7055 15895
rect 8493 15657 8527 15691
rect 9873 15589 9907 15623
rect 5917 15521 5951 15555
rect 6745 15521 6779 15555
rect 8309 15521 8343 15555
rect 5089 15453 5123 15487
rect 5273 15453 5307 15487
rect 5457 15453 5491 15487
rect 6929 15453 6963 15487
rect 7021 15453 7055 15487
rect 7849 15453 7883 15487
rect 8585 15453 8619 15487
rect 5181 15385 5215 15419
rect 6101 15385 6135 15419
rect 6285 15385 6319 15419
rect 7573 15385 7607 15419
rect 7757 15385 7791 15419
rect 8309 15385 8343 15419
rect 9321 15385 9355 15419
rect 9873 15385 9907 15419
rect 4905 15317 4939 15351
rect 6745 15317 6779 15351
rect 7665 15317 7699 15351
rect 9137 15317 9171 15351
rect 9413 15317 9447 15351
rect 4721 15113 4755 15147
rect 7757 15113 7791 15147
rect 10609 15113 10643 15147
rect 4629 15045 4663 15079
rect 5825 15045 5859 15079
rect 9873 15045 9907 15079
rect 2237 14977 2271 15011
rect 3433 14977 3467 15011
rect 5641 14977 5675 15011
rect 7113 14977 7147 15011
rect 7205 14977 7239 15011
rect 7941 14977 7975 15011
rect 8769 14977 8803 15011
rect 9045 14977 9079 15011
rect 10057 14977 10091 15011
rect 10517 14977 10551 15011
rect 10701 14977 10735 15011
rect 2329 14909 2363 14943
rect 2421 14909 2455 14943
rect 3525 14909 3559 14943
rect 3709 14909 3743 14943
rect 4905 14909 4939 14943
rect 6929 14909 6963 14943
rect 7021 14909 7055 14943
rect 8125 14909 8159 14943
rect 9137 14909 9171 14943
rect 8953 14841 8987 14875
rect 1869 14773 1903 14807
rect 3065 14773 3099 14807
rect 4261 14773 4295 14807
rect 5457 14773 5491 14807
rect 6745 14773 6779 14807
rect 8861 14773 8895 14807
rect 9689 14773 9723 14807
rect 4721 14569 4755 14603
rect 8493 14569 8527 14603
rect 9229 14569 9263 14603
rect 9321 14569 9355 14603
rect 9965 14569 9999 14603
rect 2789 14433 2823 14467
rect 2973 14433 3007 14467
rect 9413 14433 9447 14467
rect 2053 14365 2087 14399
rect 3065 14365 3099 14399
rect 3985 14365 4019 14399
rect 4905 14365 4939 14399
rect 4997 14365 5031 14399
rect 5365 14365 5399 14399
rect 6837 14365 6871 14399
rect 6929 14365 6963 14399
rect 7113 14365 7147 14399
rect 7205 14365 7239 14399
rect 8401 14365 8435 14399
rect 8585 14365 8619 14399
rect 9137 14365 9171 14399
rect 9873 14365 9907 14399
rect 10057 14365 10091 14399
rect 5089 14297 5123 14331
rect 5207 14297 5241 14331
rect 2237 14229 2271 14263
rect 3433 14229 3467 14263
rect 4169 14229 4203 14263
rect 6653 14229 6687 14263
rect 2789 14025 2823 14059
rect 3249 14025 3283 14059
rect 8217 13957 8251 13991
rect 2145 13889 2179 13923
rect 3157 13889 3191 13923
rect 6837 13889 6871 13923
rect 8401 13889 8435 13923
rect 8953 13889 8987 13923
rect 10333 13889 10367 13923
rect 10517 13889 10551 13923
rect 3433 13821 3467 13855
rect 6561 13821 6595 13855
rect 9045 13821 9079 13855
rect 6653 13753 6687 13787
rect 1961 13685 1995 13719
rect 6745 13685 6779 13719
rect 10425 13685 10459 13719
rect 11069 13685 11103 13719
rect 10885 13481 10919 13515
rect 12541 13481 12575 13515
rect 4721 13413 4755 13447
rect 5273 13413 5307 13447
rect 10425 13413 10459 13447
rect 2697 13345 2731 13379
rect 8217 13345 8251 13379
rect 10701 13345 10735 13379
rect 11989 13345 12023 13379
rect 2513 13277 2547 13311
rect 3985 13277 4019 13311
rect 6193 13277 6227 13311
rect 6377 13277 6411 13311
rect 8125 13277 8159 13311
rect 10609 13277 10643 13311
rect 10885 13277 10919 13311
rect 11713 13277 11747 13311
rect 11805 13277 11839 13311
rect 11897 13277 11931 13311
rect 12547 13277 12581 13311
rect 12725 13277 12759 13311
rect 13461 13277 13495 13311
rect 2605 13209 2639 13243
rect 7941 13209 7975 13243
rect 9873 13209 9907 13243
rect 13369 13209 13403 13243
rect 2145 13141 2179 13175
rect 3341 13141 3375 13175
rect 4077 13141 4111 13175
rect 6285 13141 6319 13175
rect 8585 13141 8619 13175
rect 11529 13141 11563 13175
rect 1869 12937 1903 12971
rect 5181 12937 5215 12971
rect 6561 12937 6595 12971
rect 6929 12937 6963 12971
rect 7021 12937 7055 12971
rect 7941 12937 7975 12971
rect 12725 12937 12759 12971
rect 3157 12869 3191 12903
rect 3985 12869 4019 12903
rect 12449 12869 12483 12903
rect 2053 12801 2087 12835
rect 2881 12801 2915 12835
rect 2973 12801 3007 12835
rect 3617 12801 3651 12835
rect 3709 12801 3743 12835
rect 3893 12801 3927 12835
rect 4077 12801 4111 12835
rect 5089 12801 5123 12835
rect 7941 12801 7975 12835
rect 9229 12801 9263 12835
rect 9689 12801 9723 12835
rect 9873 12801 9907 12835
rect 10149 12801 10183 12835
rect 10333 12801 10367 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 12081 12801 12115 12835
rect 12173 12801 12207 12835
rect 12357 12801 12391 12835
rect 12541 12801 12575 12835
rect 13553 12801 13587 12835
rect 14197 12801 14231 12835
rect 14381 12801 14415 12835
rect 2237 12733 2271 12767
rect 5273 12733 5307 12767
rect 7205 12733 7239 12767
rect 8953 12733 8987 12767
rect 9137 12733 9171 12767
rect 13737 12733 13771 12767
rect 3157 12665 3191 12699
rect 11069 12665 11103 12699
rect 4261 12597 4295 12631
rect 4721 12597 4755 12631
rect 9229 12597 9263 12631
rect 13369 12597 13403 12631
rect 14289 12597 14323 12631
rect 3433 12393 3467 12427
rect 4077 12393 4111 12427
rect 5181 12393 5215 12427
rect 9597 12393 9631 12427
rect 10517 12393 10551 12427
rect 13093 12393 13127 12427
rect 12541 12325 12575 12359
rect 1961 12257 1995 12291
rect 2145 12257 2179 12291
rect 4353 12257 4387 12291
rect 11161 12257 11195 12291
rect 13001 12257 13035 12291
rect 14289 12257 14323 12291
rect 3249 12189 3283 12223
rect 4445 12189 4479 12223
rect 5365 12189 5399 12223
rect 5549 12189 5583 12223
rect 6009 12189 6043 12223
rect 6377 12189 6411 12223
rect 7297 12189 7331 12223
rect 7481 12189 7515 12223
rect 7665 12189 7699 12223
rect 8401 12189 8435 12223
rect 9321 12189 9355 12223
rect 9413 12189 9447 12223
rect 9689 12189 9723 12223
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 12725 12189 12759 12223
rect 13277 12189 13311 12223
rect 14565 12189 14599 12223
rect 14749 12189 14783 12223
rect 2237 12121 2271 12155
rect 3065 12121 3099 12155
rect 3985 12121 4019 12155
rect 7389 12121 7423 12155
rect 12817 12121 12851 12155
rect 14427 12121 14461 12155
rect 14657 12121 14691 12155
rect 2605 12053 2639 12087
rect 4629 12053 4663 12087
rect 7113 12053 7147 12087
rect 8217 12053 8251 12087
rect 9137 12053 9171 12087
rect 11253 12053 11287 12087
rect 11345 12053 11379 12087
rect 11713 12053 11747 12087
rect 14933 12053 14967 12087
rect 4261 11849 4295 11883
rect 5641 11849 5675 11883
rect 8953 11849 8987 11883
rect 11069 11849 11103 11883
rect 11713 11849 11747 11883
rect 14105 11849 14139 11883
rect 14565 11849 14599 11883
rect 8309 11781 8343 11815
rect 1961 11713 1995 11747
rect 2697 11713 2731 11747
rect 5457 11713 5491 11747
rect 7113 11713 7147 11747
rect 8769 11713 8803 11747
rect 9781 11713 9815 11747
rect 10977 11713 11011 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 12265 11713 12299 11747
rect 13553 11713 13587 11747
rect 13921 11713 13955 11747
rect 14749 11713 14783 11747
rect 14933 11713 14967 11747
rect 2237 11645 2271 11679
rect 3801 11645 3835 11679
rect 3893 11645 3927 11679
rect 5181 11645 5215 11679
rect 7205 11645 7239 11679
rect 7389 11645 7423 11679
rect 8677 11645 8711 11679
rect 9413 11645 9447 11679
rect 9689 11645 9723 11679
rect 2053 11577 2087 11611
rect 2881 11577 2915 11611
rect 2145 11509 2179 11543
rect 3617 11509 3651 11543
rect 5273 11509 5307 11543
rect 6745 11509 6779 11543
rect 8769 11509 8803 11543
rect 12173 11509 12207 11543
rect 13921 11509 13955 11543
rect 2973 11305 3007 11339
rect 6469 11305 6503 11339
rect 11345 11305 11379 11339
rect 14381 11305 14415 11339
rect 1777 11237 1811 11271
rect 8309 11237 8343 11271
rect 11805 11237 11839 11271
rect 7297 11169 7331 11203
rect 7757 11169 7791 11203
rect 1777 11101 1811 11135
rect 2053 11101 2087 11135
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 4537 11101 4571 11135
rect 5181 11101 5215 11135
rect 5825 11101 5859 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 7389 11101 7423 11135
rect 8401 11101 8435 11135
rect 9965 11101 9999 11135
rect 10232 11101 10266 11135
rect 11989 11101 12023 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 1961 11033 1995 11067
rect 7665 11033 7699 11067
rect 4353 10965 4387 10999
rect 4997 10965 5031 10999
rect 6009 10965 6043 10999
rect 7113 10965 7147 10999
rect 2973 10761 3007 10795
rect 4813 10761 4847 10795
rect 7941 10761 7975 10795
rect 11161 10761 11195 10795
rect 11897 10761 11931 10795
rect 13553 10761 13587 10795
rect 14749 10761 14783 10795
rect 3678 10693 3712 10727
rect 6828 10693 6862 10727
rect 10048 10693 10082 10727
rect 13645 10693 13679 10727
rect 1860 10625 1894 10659
rect 8585 10625 8619 10659
rect 8677 10625 8711 10659
rect 8953 10625 8987 10659
rect 12081 10625 12115 10659
rect 12725 10625 12759 10659
rect 14381 10625 14415 10659
rect 14565 10625 14599 10659
rect 15209 10625 15243 10659
rect 15393 10625 15427 10659
rect 1593 10557 1627 10591
rect 3433 10557 3467 10591
rect 6561 10557 6595 10591
rect 8861 10557 8895 10591
rect 9781 10557 9815 10591
rect 13737 10557 13771 10591
rect 13185 10489 13219 10523
rect 8401 10421 8435 10455
rect 12541 10421 12575 10455
rect 15301 10421 15335 10455
rect 1593 10217 1627 10251
rect 5733 10217 5767 10251
rect 7573 10217 7607 10251
rect 12817 10217 12851 10251
rect 11529 10149 11563 10183
rect 6193 10081 6227 10115
rect 13461 10081 13495 10115
rect 14381 10081 14415 10115
rect 2973 10013 3007 10047
rect 4353 10013 4387 10047
rect 4620 10013 4654 10047
rect 10149 10013 10183 10047
rect 10416 10013 10450 10047
rect 14657 10013 14691 10047
rect 14749 10013 14783 10047
rect 16221 10013 16255 10047
rect 16589 10013 16623 10047
rect 16957 10013 16991 10047
rect 2728 9945 2762 9979
rect 6438 9945 6472 9979
rect 13185 9945 13219 9979
rect 14289 9945 14323 9979
rect 13277 9877 13311 9911
rect 14933 9877 14967 9911
rect 15669 9877 15703 9911
rect 1860 9605 1894 9639
rect 4252 9605 4286 9639
rect 9422 9605 9456 9639
rect 13369 9605 13403 9639
rect 15577 9605 15611 9639
rect 3985 9537 4019 9571
rect 13461 9537 13495 9571
rect 14197 9537 14231 9571
rect 14381 9537 14415 9571
rect 16865 9537 16899 9571
rect 1593 9469 1627 9503
rect 9689 9469 9723 9503
rect 13553 9469 13587 9503
rect 14657 9469 14691 9503
rect 2973 9401 3007 9435
rect 5365 9401 5399 9435
rect 14565 9401 14599 9435
rect 17141 9401 17175 9435
rect 8309 9333 8343 9367
rect 13001 9333 13035 9367
rect 17325 9333 17359 9367
rect 5365 9129 5399 9163
rect 8585 9129 8619 9163
rect 13369 9129 13403 9163
rect 11529 9061 11563 9095
rect 16037 9061 16071 9095
rect 16681 9061 16715 9095
rect 18337 9061 18371 9095
rect 19625 9061 19659 9095
rect 7205 8993 7239 9027
rect 10149 8993 10183 9027
rect 15899 8993 15933 9027
rect 3985 8925 4019 8959
rect 4252 8925 4286 8959
rect 7472 8925 7506 8959
rect 12909 8925 12943 8959
rect 13645 8925 13679 8959
rect 15761 8925 15795 8959
rect 16221 8925 16255 8959
rect 16681 8925 16715 8959
rect 16865 8925 16899 8959
rect 17417 8925 17451 8959
rect 17601 8925 17635 8959
rect 18061 8925 18095 8959
rect 19809 8925 19843 8959
rect 10416 8857 10450 8891
rect 13369 8857 13403 8891
rect 13553 8857 13587 8891
rect 18153 8857 18187 8891
rect 18337 8857 18371 8891
rect 12725 8789 12759 8823
rect 16221 8789 16255 8823
rect 17417 8789 17451 8823
rect 3617 8585 3651 8619
rect 7481 8585 7515 8619
rect 11161 8585 11195 8619
rect 16865 8585 16899 8619
rect 18061 8585 18095 8619
rect 2482 8517 2516 8551
rect 10048 8517 10082 8551
rect 19993 8517 20027 8551
rect 20913 8517 20947 8551
rect 4077 8449 4111 8483
rect 8605 8449 8639 8483
rect 8861 8449 8895 8483
rect 9781 8449 9815 8483
rect 13829 8449 13863 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 14197 8449 14231 8483
rect 14841 8449 14875 8483
rect 15761 8449 15795 8483
rect 15945 8449 15979 8483
rect 17049 8449 17083 8483
rect 17233 8449 17267 8483
rect 17877 8449 17911 8483
rect 18061 8449 18095 8483
rect 18797 8449 18831 8483
rect 18981 8449 19015 8483
rect 19073 8449 19107 8483
rect 19257 8449 19291 8483
rect 19717 8449 19751 8483
rect 19810 8449 19844 8483
rect 20085 8449 20119 8483
rect 20223 8449 20257 8483
rect 20821 8449 20855 8483
rect 21005 8449 21039 8483
rect 2237 8381 2271 8415
rect 14657 8381 14691 8415
rect 15025 8381 15059 8415
rect 17141 8381 17175 8415
rect 17325 8381 17359 8415
rect 18613 8381 18647 8415
rect 4169 8313 4203 8347
rect 15853 8313 15887 8347
rect 18889 8313 18923 8347
rect 20361 8313 20395 8347
rect 5089 8245 5123 8279
rect 13645 8245 13679 8279
rect 6561 8041 6595 8075
rect 8585 8041 8619 8075
rect 11529 8041 11563 8075
rect 15209 8041 15243 8075
rect 17785 8041 17819 8075
rect 18613 8041 18647 8075
rect 18797 8041 18831 8075
rect 19625 8041 19659 8075
rect 14473 7973 14507 8007
rect 1593 7905 1627 7939
rect 7205 7905 7239 7939
rect 10149 7905 10183 7939
rect 14289 7905 14323 7939
rect 15669 7905 15703 7939
rect 15853 7905 15887 7939
rect 19717 7905 19751 7939
rect 4077 7837 4111 7871
rect 4261 7831 4295 7865
rect 4356 7837 4390 7871
rect 4445 7837 4479 7871
rect 5181 7837 5215 7871
rect 12357 7837 12391 7871
rect 13277 7837 13311 7871
rect 13369 7837 13403 7871
rect 13645 7837 13679 7871
rect 13737 7837 13771 7871
rect 14565 7837 14599 7871
rect 16405 7837 16439 7871
rect 16589 7837 16623 7871
rect 19441 7837 19475 7871
rect 19533 7837 19567 7871
rect 20361 7837 20395 7871
rect 1860 7769 1894 7803
rect 5448 7769 5482 7803
rect 7472 7769 7506 7803
rect 10416 7769 10450 7803
rect 13461 7769 13495 7803
rect 17601 7769 17635 7803
rect 17801 7769 17835 7803
rect 18429 7769 18463 7803
rect 2973 7701 3007 7735
rect 4721 7701 4755 7735
rect 12449 7701 12483 7735
rect 13001 7701 13035 7735
rect 14565 7701 14599 7735
rect 15577 7701 15611 7735
rect 16773 7701 16807 7735
rect 17969 7701 18003 7735
rect 18629 7701 18663 7735
rect 20269 7701 20303 7735
rect 1961 7497 1995 7531
rect 5273 7497 5307 7531
rect 14013 7497 14047 7531
rect 16313 7497 16347 7531
rect 17417 7497 17451 7531
rect 2605 7429 2639 7463
rect 4353 7429 4387 7463
rect 7849 7429 7883 7463
rect 9597 7429 9631 7463
rect 15301 7429 15335 7463
rect 19901 7429 19935 7463
rect 2145 7361 2179 7395
rect 5181 7361 5215 7395
rect 6561 7361 6595 7395
rect 13093 7361 13127 7395
rect 13277 7361 13311 7395
rect 13369 7361 13403 7395
rect 14105 7361 14139 7395
rect 15209 7361 15243 7395
rect 15485 7361 15519 7395
rect 15945 7361 15979 7395
rect 16129 7361 16163 7395
rect 17693 7361 17727 7395
rect 18429 7361 18463 7395
rect 18613 7361 18647 7395
rect 18705 7361 18739 7395
rect 18889 7361 18923 7395
rect 18981 7361 19015 7395
rect 5457 7293 5491 7327
rect 13185 7293 13219 7327
rect 17601 7293 17635 7327
rect 17785 7293 17819 7327
rect 17877 7293 17911 7327
rect 4813 7225 4847 7259
rect 15485 7225 15519 7259
rect 20177 7225 20211 7259
rect 6653 7157 6687 7191
rect 7205 7157 7239 7191
rect 12909 7157 12943 7191
rect 16037 7157 16071 7191
rect 20361 7157 20395 7191
rect 16405 6953 16439 6987
rect 15761 6885 15795 6919
rect 9781 6817 9815 6851
rect 15577 6817 15611 6851
rect 19625 6817 19659 6851
rect 19809 6817 19843 6851
rect 19901 6817 19935 6851
rect 3157 6749 3191 6783
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 4721 6749 4755 6783
rect 4813 6749 4847 6783
rect 10048 6749 10082 6783
rect 13277 6749 13311 6783
rect 14473 6749 14507 6783
rect 15853 6749 15887 6783
rect 16313 6749 16347 6783
rect 16497 6749 16531 6783
rect 19717 6749 19751 6783
rect 5089 6681 5123 6715
rect 5917 6681 5951 6715
rect 8125 6681 8159 6715
rect 13001 6681 13035 6715
rect 13185 6681 13219 6715
rect 15577 6681 15611 6715
rect 2973 6613 3007 6647
rect 7389 6613 7423 6647
rect 11161 6613 11195 6647
rect 13099 6613 13133 6647
rect 14381 6613 14415 6647
rect 19441 6613 19475 6647
rect 2973 6409 3007 6443
rect 6009 6409 6043 6443
rect 7849 6409 7883 6443
rect 11069 6409 11103 6443
rect 12725 6409 12759 6443
rect 17509 6409 17543 6443
rect 4874 6341 4908 6375
rect 7021 6341 7055 6375
rect 8984 6341 9018 6375
rect 13277 6341 13311 6375
rect 15393 6341 15427 6375
rect 17141 6341 17175 6375
rect 18889 6341 18923 6375
rect 20913 6341 20947 6375
rect 1860 6273 1894 6307
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 4629 6273 4663 6307
rect 6653 6273 6687 6307
rect 9956 6273 9990 6307
rect 13001 6273 13035 6307
rect 13829 6273 13863 6307
rect 14013 6273 14047 6307
rect 14105 6273 14139 6307
rect 14381 6273 14415 6307
rect 15577 6273 15611 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 15945 6273 15979 6307
rect 16865 6273 16899 6307
rect 16958 6273 16992 6307
rect 17233 6273 17267 6307
rect 17330 6273 17364 6307
rect 18797 6273 18831 6307
rect 18981 6273 19015 6307
rect 19165 6273 19199 6307
rect 20085 6273 20119 6307
rect 20821 6273 20855 6307
rect 21005 6273 21039 6307
rect 1593 6205 1627 6239
rect 4169 6205 4203 6239
rect 9229 6205 9263 6239
rect 9689 6205 9723 6239
rect 12909 6205 12943 6239
rect 13369 6205 13403 6239
rect 20361 6205 20395 6239
rect 20269 6137 20303 6171
rect 3617 6069 3651 6103
rect 14289 6069 14323 6103
rect 18613 6069 18647 6103
rect 20177 6069 20211 6103
rect 2697 5865 2731 5899
rect 4813 5865 4847 5899
rect 12725 5865 12759 5899
rect 14289 5865 14323 5899
rect 16865 5865 16899 5899
rect 19441 5865 19475 5899
rect 19809 5865 19843 5899
rect 11437 5797 11471 5831
rect 15853 5797 15887 5831
rect 19993 5797 20027 5831
rect 21005 5797 21039 5831
rect 4629 5729 4663 5763
rect 14657 5729 14691 5763
rect 14749 5729 14783 5763
rect 16313 5729 16347 5763
rect 20913 5729 20947 5763
rect 2881 5661 2915 5695
rect 3157 5661 3191 5695
rect 3341 5661 3375 5695
rect 4169 5661 4203 5695
rect 4537 5661 4571 5695
rect 6561 5661 6595 5695
rect 6828 5661 6862 5695
rect 10057 5661 10091 5695
rect 12081 5661 12115 5695
rect 12265 5661 12299 5695
rect 12906 5661 12940 5695
rect 13277 5661 13311 5695
rect 13369 5661 13403 5695
rect 14473 5661 14507 5695
rect 14841 5661 14875 5695
rect 15025 5661 15059 5695
rect 16037 5661 16071 5695
rect 16129 5661 16163 5695
rect 16405 5661 16439 5695
rect 16865 5661 16899 5695
rect 17049 5661 17083 5695
rect 17693 5661 17727 5695
rect 17877 5661 17911 5695
rect 17969 5661 18003 5695
rect 18061 5661 18095 5695
rect 19717 5661 19751 5695
rect 19901 5661 19935 5695
rect 20177 5661 20211 5695
rect 20821 5661 20855 5695
rect 21097 5661 21131 5695
rect 5733 5593 5767 5627
rect 10324 5593 10358 5627
rect 12173 5593 12207 5627
rect 4261 5525 4295 5559
rect 4353 5525 4387 5559
rect 6009 5525 6043 5559
rect 7941 5525 7975 5559
rect 12909 5525 12943 5559
rect 18337 5525 18371 5559
rect 20637 5525 20671 5559
rect 4537 5321 4571 5355
rect 4721 5321 4755 5355
rect 5181 5321 5215 5355
rect 7849 5321 7883 5355
rect 12909 5321 12943 5355
rect 14105 5321 14139 5355
rect 18797 5321 18831 5355
rect 19257 5321 19291 5355
rect 5333 5253 5367 5287
rect 5549 5253 5583 5287
rect 8984 5253 9018 5287
rect 13553 5253 13587 5287
rect 16313 5253 16347 5287
rect 17785 5253 17819 5287
rect 19809 5253 19843 5287
rect 19901 5253 19935 5287
rect 1860 5185 1894 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4353 5185 4387 5219
rect 4445 5185 4479 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 10048 5185 10082 5219
rect 13093 5185 13127 5219
rect 13185 5185 13219 5219
rect 14473 5185 14507 5219
rect 14565 5185 14599 5219
rect 16037 5185 16071 5219
rect 17601 5185 17635 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 19441 5185 19475 5219
rect 19533 5185 19567 5219
rect 1593 5117 1627 5151
rect 3893 5117 3927 5151
rect 4721 5117 4755 5151
rect 9229 5117 9263 5151
rect 9781 5117 9815 5151
rect 13461 5117 13495 5151
rect 14749 5117 14783 5151
rect 17417 5117 17451 5151
rect 2973 5049 3007 5083
rect 3801 4981 3835 5015
rect 5365 4981 5399 5015
rect 6561 4981 6595 5015
rect 7297 4981 7331 5015
rect 11161 4981 11195 5015
rect 16957 4981 16991 5015
rect 18521 4981 18555 5015
rect 7389 4777 7423 4811
rect 13553 4777 13587 4811
rect 14289 4777 14323 4811
rect 15853 4777 15887 4811
rect 16037 4777 16071 4811
rect 16773 4777 16807 4811
rect 17969 4777 18003 4811
rect 18705 4777 18739 4811
rect 19441 4777 19475 4811
rect 3985 4709 4019 4743
rect 6009 4641 6043 4675
rect 15485 4641 15519 4675
rect 4261 4573 4295 4607
rect 13737 4573 13771 4607
rect 14565 4573 14599 4607
rect 14657 4573 14691 4607
rect 14749 4573 14783 4607
rect 14933 4573 14967 4607
rect 16589 4573 16623 4607
rect 16773 4573 16807 4607
rect 17417 4573 17451 4607
rect 17877 4573 17911 4607
rect 18061 4573 18095 4607
rect 18705 4573 18739 4607
rect 18889 4573 18923 4607
rect 19441 4573 19475 4607
rect 19625 4573 19659 4607
rect 3985 4505 4019 4539
rect 6276 4505 6310 4539
rect 15853 4505 15887 4539
rect 17325 4505 17359 4539
rect 4169 4437 4203 4471
rect 5549 4437 5583 4471
rect 15393 4233 15427 4267
rect 17693 4233 17727 4267
rect 18981 4233 19015 4267
rect 14013 4165 14047 4199
rect 2688 4097 2722 4131
rect 4629 4097 4663 4131
rect 4896 4097 4930 4131
rect 7113 4097 7147 4131
rect 7389 4097 7423 4131
rect 8962 4097 8996 4131
rect 9229 4097 9263 4131
rect 9689 4097 9723 4131
rect 9956 4097 9990 4131
rect 12081 4097 12115 4131
rect 13001 4097 13035 4131
rect 14197 4097 14231 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 15853 4097 15887 4131
rect 17325 4097 17359 4131
rect 17509 4097 17543 4131
rect 18984 4097 19018 4131
rect 19625 4097 19659 4131
rect 19809 4097 19843 4131
rect 2421 4029 2455 4063
rect 13093 4029 13127 4063
rect 14933 4029 14967 4063
rect 18521 4029 18555 4063
rect 19717 4029 19751 4063
rect 7297 3961 7331 3995
rect 12265 3961 12299 3995
rect 13369 3961 13403 3995
rect 3801 3893 3835 3927
rect 6009 3893 6043 3927
rect 7205 3893 7239 3927
rect 7849 3893 7883 3927
rect 11069 3893 11103 3927
rect 14289 3893 14323 3927
rect 17325 3893 17359 3927
rect 18613 3893 18647 3927
rect 19165 3893 19199 3927
rect 3065 3689 3099 3723
rect 5549 3689 5583 3723
rect 6101 3689 6135 3723
rect 6469 3689 6503 3723
rect 12449 3689 12483 3723
rect 14381 3689 14415 3723
rect 14749 3689 14783 3723
rect 16589 3689 16623 3723
rect 19625 3689 19659 3723
rect 19809 3689 19843 3723
rect 11897 3621 11931 3655
rect 15853 3621 15887 3655
rect 18613 3621 18647 3655
rect 20269 3621 20303 3655
rect 4169 3553 4203 3587
rect 6561 3553 6595 3587
rect 7021 3553 7055 3587
rect 9965 3553 9999 3587
rect 13001 3553 13035 3587
rect 13093 3553 13127 3587
rect 13277 3553 13311 3587
rect 13461 3553 13495 3587
rect 16497 3553 16531 3587
rect 18521 3553 18555 3587
rect 21005 3553 21039 3587
rect 3249 3485 3283 3519
rect 3433 3485 3467 3519
rect 6285 3485 6319 3519
rect 7277 3485 7311 3519
rect 10232 3485 10266 3519
rect 13185 3485 13219 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 16589 3485 16623 3519
rect 17509 3485 17543 3519
rect 18153 3485 18187 3519
rect 18337 3485 18371 3519
rect 18429 3485 18463 3519
rect 19441 3485 19475 3519
rect 19625 3485 19659 3519
rect 20545 3485 20579 3519
rect 4436 3417 4470 3451
rect 12081 3417 12115 3451
rect 12173 3417 12207 3451
rect 12265 3417 12299 3451
rect 15669 3417 15703 3451
rect 16313 3417 16347 3451
rect 17325 3417 17359 3451
rect 17693 3417 17727 3451
rect 20269 3417 20303 3451
rect 20453 3417 20487 3451
rect 8401 3349 8435 3383
rect 11345 3349 11379 3383
rect 16773 3349 16807 3383
rect 18889 3349 18923 3383
rect 4813 3145 4847 3179
rect 7113 3145 7147 3179
rect 7205 3145 7239 3179
rect 10241 3145 10275 3179
rect 15777 3145 15811 3179
rect 18429 3145 18463 3179
rect 19625 3145 19659 3179
rect 2697 3077 2731 3111
rect 4353 3077 4387 3111
rect 7849 3077 7883 3111
rect 9505 3077 9539 3111
rect 11161 3077 11195 3111
rect 15577 3077 15611 3111
rect 4997 3009 5031 3043
rect 5181 3009 5215 3043
rect 5273 3009 5307 3043
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 7021 3009 7055 3043
rect 10057 3009 10091 3043
rect 10333 3009 10367 3043
rect 10885 3009 10919 3043
rect 10977 3009 11011 3043
rect 11989 3009 12023 3043
rect 12081 3009 12115 3043
rect 12173 3009 12207 3043
rect 13461 3009 13495 3043
rect 14933 3009 14967 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 18797 3009 18831 3043
rect 18889 3009 18923 3043
rect 19073 3009 19107 3043
rect 19717 3009 19751 3043
rect 5733 2941 5767 2975
rect 7389 2941 7423 2975
rect 11897 2941 11931 2975
rect 13185 2941 13219 2975
rect 15025 2941 15059 2975
rect 16957 2941 16991 2975
rect 17693 2941 17727 2975
rect 14565 2873 14599 2907
rect 10057 2805 10091 2839
rect 11161 2805 11195 2839
rect 11713 2805 11747 2839
rect 12909 2805 12943 2839
rect 13093 2805 13127 2839
rect 15761 2805 15795 2839
rect 15945 2805 15979 2839
rect 16865 2805 16899 2839
rect 17233 2805 17267 2839
rect 3065 2601 3099 2635
rect 3985 2601 4019 2635
rect 5089 2601 5123 2635
rect 5733 2601 5767 2635
rect 7205 2601 7239 2635
rect 7389 2601 7423 2635
rect 8033 2601 8067 2635
rect 9137 2601 9171 2635
rect 9505 2601 9539 2635
rect 11069 2601 11103 2635
rect 12081 2601 12115 2635
rect 12725 2601 12759 2635
rect 15209 2601 15243 2635
rect 15945 2601 15979 2635
rect 16957 2601 16991 2635
rect 18613 2601 18647 2635
rect 3157 2533 3191 2567
rect 4353 2465 4387 2499
rect 3249 2397 3283 2431
rect 4169 2397 4203 2431
rect 4813 2397 4847 2431
rect 4905 2397 4939 2431
rect 5733 2397 5767 2431
rect 5917 2397 5951 2431
rect 8033 2397 8067 2431
rect 8293 2375 8327 2409
rect 9321 2397 9355 2431
rect 9597 2397 9631 2431
rect 11713 2397 11747 2431
rect 13369 2397 13403 2431
rect 15669 2397 15703 2431
rect 17049 2397 17083 2431
rect 18337 2397 18371 2431
rect 2973 2329 3007 2363
rect 5089 2329 5123 2363
rect 7573 2329 7607 2363
rect 11897 2329 11931 2363
rect 15761 2329 15795 2363
rect 15945 2329 15979 2363
rect 17601 2329 17635 2363
rect 18613 2329 18647 2363
rect 7373 2261 7407 2295
rect 8217 2261 8251 2295
rect 13553 2261 13587 2295
rect 18429 2261 18463 2295
<< metal1 >>
rect 1104 21786 22976 21808
rect 1104 21734 6378 21786
rect 6430 21734 6442 21786
rect 6494 21734 6506 21786
rect 6558 21734 6570 21786
rect 6622 21734 6634 21786
rect 6686 21734 11806 21786
rect 11858 21734 11870 21786
rect 11922 21734 11934 21786
rect 11986 21734 11998 21786
rect 12050 21734 12062 21786
rect 12114 21734 17234 21786
rect 17286 21734 17298 21786
rect 17350 21734 17362 21786
rect 17414 21734 17426 21786
rect 17478 21734 17490 21786
rect 17542 21734 22662 21786
rect 22714 21734 22726 21786
rect 22778 21734 22790 21786
rect 22842 21734 22854 21786
rect 22906 21734 22918 21786
rect 22970 21734 22976 21786
rect 1104 21712 22976 21734
rect 1104 21242 22816 21264
rect 1104 21190 3664 21242
rect 3716 21190 3728 21242
rect 3780 21190 3792 21242
rect 3844 21190 3856 21242
rect 3908 21190 3920 21242
rect 3972 21190 9092 21242
rect 9144 21190 9156 21242
rect 9208 21190 9220 21242
rect 9272 21190 9284 21242
rect 9336 21190 9348 21242
rect 9400 21190 14520 21242
rect 14572 21190 14584 21242
rect 14636 21190 14648 21242
rect 14700 21190 14712 21242
rect 14764 21190 14776 21242
rect 14828 21190 19948 21242
rect 20000 21190 20012 21242
rect 20064 21190 20076 21242
rect 20128 21190 20140 21242
rect 20192 21190 20204 21242
rect 20256 21190 22816 21242
rect 1104 21168 22816 21190
rect 1104 20698 22976 20720
rect 1104 20646 6378 20698
rect 6430 20646 6442 20698
rect 6494 20646 6506 20698
rect 6558 20646 6570 20698
rect 6622 20646 6634 20698
rect 6686 20646 11806 20698
rect 11858 20646 11870 20698
rect 11922 20646 11934 20698
rect 11986 20646 11998 20698
rect 12050 20646 12062 20698
rect 12114 20646 17234 20698
rect 17286 20646 17298 20698
rect 17350 20646 17362 20698
rect 17414 20646 17426 20698
rect 17478 20646 17490 20698
rect 17542 20646 22662 20698
rect 22714 20646 22726 20698
rect 22778 20646 22790 20698
rect 22842 20646 22854 20698
rect 22906 20646 22918 20698
rect 22970 20646 22976 20698
rect 1104 20624 22976 20646
rect 1104 20154 22816 20176
rect 1104 20102 3664 20154
rect 3716 20102 3728 20154
rect 3780 20102 3792 20154
rect 3844 20102 3856 20154
rect 3908 20102 3920 20154
rect 3972 20102 9092 20154
rect 9144 20102 9156 20154
rect 9208 20102 9220 20154
rect 9272 20102 9284 20154
rect 9336 20102 9348 20154
rect 9400 20102 14520 20154
rect 14572 20102 14584 20154
rect 14636 20102 14648 20154
rect 14700 20102 14712 20154
rect 14764 20102 14776 20154
rect 14828 20102 19948 20154
rect 20000 20102 20012 20154
rect 20064 20102 20076 20154
rect 20128 20102 20140 20154
rect 20192 20102 20204 20154
rect 20256 20102 22816 20154
rect 1104 20080 22816 20102
rect 1104 19610 22976 19632
rect 1104 19558 6378 19610
rect 6430 19558 6442 19610
rect 6494 19558 6506 19610
rect 6558 19558 6570 19610
rect 6622 19558 6634 19610
rect 6686 19558 11806 19610
rect 11858 19558 11870 19610
rect 11922 19558 11934 19610
rect 11986 19558 11998 19610
rect 12050 19558 12062 19610
rect 12114 19558 17234 19610
rect 17286 19558 17298 19610
rect 17350 19558 17362 19610
rect 17414 19558 17426 19610
rect 17478 19558 17490 19610
rect 17542 19558 22662 19610
rect 22714 19558 22726 19610
rect 22778 19558 22790 19610
rect 22842 19558 22854 19610
rect 22906 19558 22918 19610
rect 22970 19558 22976 19610
rect 1104 19536 22976 19558
rect 2130 19496 2136 19508
rect 2091 19468 2136 19496
rect 2130 19456 2136 19468
rect 2188 19456 2194 19508
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 1949 19363 2007 19369
rect 1949 19360 1961 19363
rect 1912 19332 1961 19360
rect 1912 19320 1918 19332
rect 1949 19329 1961 19332
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 1104 19066 22816 19088
rect 1104 19014 3664 19066
rect 3716 19014 3728 19066
rect 3780 19014 3792 19066
rect 3844 19014 3856 19066
rect 3908 19014 3920 19066
rect 3972 19014 9092 19066
rect 9144 19014 9156 19066
rect 9208 19014 9220 19066
rect 9272 19014 9284 19066
rect 9336 19014 9348 19066
rect 9400 19014 14520 19066
rect 14572 19014 14584 19066
rect 14636 19014 14648 19066
rect 14700 19014 14712 19066
rect 14764 19014 14776 19066
rect 14828 19014 19948 19066
rect 20000 19014 20012 19066
rect 20064 19014 20076 19066
rect 20128 19014 20140 19066
rect 20192 19014 20204 19066
rect 20256 19014 22816 19066
rect 1104 18992 22816 19014
rect 1104 18522 22976 18544
rect 1104 18470 6378 18522
rect 6430 18470 6442 18522
rect 6494 18470 6506 18522
rect 6558 18470 6570 18522
rect 6622 18470 6634 18522
rect 6686 18470 11806 18522
rect 11858 18470 11870 18522
rect 11922 18470 11934 18522
rect 11986 18470 11998 18522
rect 12050 18470 12062 18522
rect 12114 18470 17234 18522
rect 17286 18470 17298 18522
rect 17350 18470 17362 18522
rect 17414 18470 17426 18522
rect 17478 18470 17490 18522
rect 17542 18470 22662 18522
rect 22714 18470 22726 18522
rect 22778 18470 22790 18522
rect 22842 18470 22854 18522
rect 22906 18470 22918 18522
rect 22970 18470 22976 18522
rect 1104 18448 22976 18470
rect 1104 17978 22816 18000
rect 1104 17926 3664 17978
rect 3716 17926 3728 17978
rect 3780 17926 3792 17978
rect 3844 17926 3856 17978
rect 3908 17926 3920 17978
rect 3972 17926 9092 17978
rect 9144 17926 9156 17978
rect 9208 17926 9220 17978
rect 9272 17926 9284 17978
rect 9336 17926 9348 17978
rect 9400 17926 14520 17978
rect 14572 17926 14584 17978
rect 14636 17926 14648 17978
rect 14700 17926 14712 17978
rect 14764 17926 14776 17978
rect 14828 17926 19948 17978
rect 20000 17926 20012 17978
rect 20064 17926 20076 17978
rect 20128 17926 20140 17978
rect 20192 17926 20204 17978
rect 20256 17926 22816 17978
rect 1104 17904 22816 17926
rect 1104 17434 22976 17456
rect 1104 17382 6378 17434
rect 6430 17382 6442 17434
rect 6494 17382 6506 17434
rect 6558 17382 6570 17434
rect 6622 17382 6634 17434
rect 6686 17382 11806 17434
rect 11858 17382 11870 17434
rect 11922 17382 11934 17434
rect 11986 17382 11998 17434
rect 12050 17382 12062 17434
rect 12114 17382 17234 17434
rect 17286 17382 17298 17434
rect 17350 17382 17362 17434
rect 17414 17382 17426 17434
rect 17478 17382 17490 17434
rect 17542 17382 22662 17434
rect 22714 17382 22726 17434
rect 22778 17382 22790 17434
rect 22842 17382 22854 17434
rect 22906 17382 22918 17434
rect 22970 17382 22976 17434
rect 1104 17360 22976 17382
rect 1104 16890 22816 16912
rect 1104 16838 3664 16890
rect 3716 16838 3728 16890
rect 3780 16838 3792 16890
rect 3844 16838 3856 16890
rect 3908 16838 3920 16890
rect 3972 16838 9092 16890
rect 9144 16838 9156 16890
rect 9208 16838 9220 16890
rect 9272 16838 9284 16890
rect 9336 16838 9348 16890
rect 9400 16838 14520 16890
rect 14572 16838 14584 16890
rect 14636 16838 14648 16890
rect 14700 16838 14712 16890
rect 14764 16838 14776 16890
rect 14828 16838 19948 16890
rect 20000 16838 20012 16890
rect 20064 16838 20076 16890
rect 20128 16838 20140 16890
rect 20192 16838 20204 16890
rect 20256 16838 22816 16890
rect 1104 16816 22816 16838
rect 1104 16346 22976 16368
rect 1104 16294 6378 16346
rect 6430 16294 6442 16346
rect 6494 16294 6506 16346
rect 6558 16294 6570 16346
rect 6622 16294 6634 16346
rect 6686 16294 11806 16346
rect 11858 16294 11870 16346
rect 11922 16294 11934 16346
rect 11986 16294 11998 16346
rect 12050 16294 12062 16346
rect 12114 16294 17234 16346
rect 17286 16294 17298 16346
rect 17350 16294 17362 16346
rect 17414 16294 17426 16346
rect 17478 16294 17490 16346
rect 17542 16294 22662 16346
rect 22714 16294 22726 16346
rect 22778 16294 22790 16346
rect 22842 16294 22854 16346
rect 22906 16294 22918 16346
rect 22970 16294 22976 16346
rect 1104 16272 22976 16294
rect 5534 16164 5540 16176
rect 5000 16136 5540 16164
rect 5000 16105 5028 16136
rect 5534 16124 5540 16136
rect 5592 16124 5598 16176
rect 4893 16099 4951 16105
rect 4893 16065 4905 16099
rect 4939 16065 4951 16099
rect 4893 16059 4951 16065
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16065 5043 16099
rect 4985 16059 5043 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5166 16096 5172 16108
rect 5123 16068 5172 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 4908 16028 4936 16059
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 6086 16096 6092 16108
rect 5951 16068 6092 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 5258 16028 5264 16040
rect 4908 16000 5264 16028
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 5736 16028 5764 16059
rect 6086 16056 6092 16068
rect 6144 16096 6150 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6144 16068 6837 16096
rect 6144 16056 6150 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16096 7067 16099
rect 8202 16096 8208 16108
rect 7055 16068 8208 16096
rect 7055 16065 7067 16068
rect 7009 16059 7067 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 6270 16028 6276 16040
rect 5736 16000 6276 16028
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 4709 15895 4767 15901
rect 4709 15892 4721 15895
rect 4120 15864 4721 15892
rect 4120 15852 4126 15864
rect 4709 15861 4721 15864
rect 4755 15861 4767 15895
rect 4709 15855 4767 15861
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 5813 15895 5871 15901
rect 5813 15892 5825 15895
rect 5592 15864 5825 15892
rect 5592 15852 5598 15864
rect 5813 15861 5825 15864
rect 5859 15861 5871 15895
rect 7006 15892 7012 15904
rect 6967 15864 7012 15892
rect 5813 15855 5871 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 1104 15802 22816 15824
rect 1104 15750 3664 15802
rect 3716 15750 3728 15802
rect 3780 15750 3792 15802
rect 3844 15750 3856 15802
rect 3908 15750 3920 15802
rect 3972 15750 9092 15802
rect 9144 15750 9156 15802
rect 9208 15750 9220 15802
rect 9272 15750 9284 15802
rect 9336 15750 9348 15802
rect 9400 15750 14520 15802
rect 14572 15750 14584 15802
rect 14636 15750 14648 15802
rect 14700 15750 14712 15802
rect 14764 15750 14776 15802
rect 14828 15750 19948 15802
rect 20000 15750 20012 15802
rect 20064 15750 20076 15802
rect 20128 15750 20140 15802
rect 20192 15750 20204 15802
rect 20256 15750 22816 15802
rect 1104 15728 22816 15750
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 8260 15660 8493 15688
rect 8260 15648 8266 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 8481 15651 8539 15657
rect 6086 15580 6092 15632
rect 6144 15620 6150 15632
rect 8110 15620 8116 15632
rect 6144 15592 8116 15620
rect 6144 15580 6150 15592
rect 8110 15580 8116 15592
rect 8168 15620 8174 15632
rect 8168 15592 8340 15620
rect 8168 15580 8174 15592
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5276 15524 5917 15552
rect 5276 15496 5304 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15552 6791 15555
rect 6822 15552 6828 15564
rect 6779 15524 6828 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15453 5135 15487
rect 5258 15484 5264 15496
rect 5219 15456 5264 15484
rect 5077 15447 5135 15453
rect 4890 15348 4896 15360
rect 4851 15320 4896 15348
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5092 15348 5120 15447
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 5445 15487 5503 15493
rect 5445 15453 5457 15487
rect 5491 15484 5503 15487
rect 5534 15484 5540 15496
rect 5491 15456 5540 15484
rect 5491 15453 5503 15456
rect 5445 15447 5503 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 6748 15484 6776 15515
rect 6822 15512 6828 15524
rect 6880 15552 6886 15564
rect 8312 15561 8340 15592
rect 8297 15555 8355 15561
rect 6880 15524 7972 15552
rect 6880 15512 6886 15524
rect 6914 15484 6920 15496
rect 5920 15456 6776 15484
rect 6875 15456 6920 15484
rect 5166 15376 5172 15428
rect 5224 15416 5230 15428
rect 5920 15416 5948 15456
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7837 15487 7895 15493
rect 7064 15456 7109 15484
rect 7208 15456 7788 15484
rect 7064 15444 7070 15456
rect 6086 15416 6092 15428
rect 5224 15388 5948 15416
rect 6047 15388 6092 15416
rect 5224 15376 5230 15388
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 6270 15376 6276 15428
rect 6328 15416 6334 15428
rect 7208 15416 7236 15456
rect 7760 15428 7788 15456
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7944 15484 7972 15524
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8496 15552 8524 15651
rect 8754 15580 8760 15632
rect 8812 15620 8818 15632
rect 9861 15623 9919 15629
rect 9861 15620 9873 15623
rect 8812 15592 9873 15620
rect 8812 15580 8818 15592
rect 9861 15589 9873 15592
rect 9907 15589 9919 15623
rect 9861 15583 9919 15589
rect 8496 15524 9904 15552
rect 8297 15515 8355 15521
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 7944 15456 8585 15484
rect 7837 15447 7895 15453
rect 8573 15453 8585 15456
rect 8619 15484 8631 15487
rect 8754 15484 8760 15496
rect 8619 15456 8760 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 7558 15416 7564 15428
rect 6328 15388 7236 15416
rect 7519 15388 7564 15416
rect 6328 15376 6334 15388
rect 7558 15376 7564 15388
rect 7616 15376 7622 15428
rect 7742 15416 7748 15428
rect 7703 15388 7748 15416
rect 7742 15376 7748 15388
rect 7800 15376 7806 15428
rect 7852 15416 7880 15447
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 7852 15388 8309 15416
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 9309 15419 9367 15425
rect 9309 15385 9321 15419
rect 9355 15416 9367 15419
rect 9582 15416 9588 15428
rect 9355 15388 9588 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 9876 15425 9904 15524
rect 9861 15419 9919 15425
rect 9861 15385 9873 15419
rect 9907 15416 9919 15419
rect 10594 15416 10600 15428
rect 9907 15388 10600 15416
rect 9907 15385 9919 15388
rect 9861 15379 9919 15385
rect 10594 15376 10600 15388
rect 10652 15376 10658 15428
rect 6288 15348 6316 15376
rect 6730 15348 6736 15360
rect 5092 15320 6316 15348
rect 6691 15320 6736 15348
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 9122 15348 9128 15360
rect 9083 15320 9128 15348
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 9398 15348 9404 15360
rect 9359 15320 9404 15348
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 1104 15258 22976 15280
rect 1104 15206 6378 15258
rect 6430 15206 6442 15258
rect 6494 15206 6506 15258
rect 6558 15206 6570 15258
rect 6622 15206 6634 15258
rect 6686 15206 11806 15258
rect 11858 15206 11870 15258
rect 11922 15206 11934 15258
rect 11986 15206 11998 15258
rect 12050 15206 12062 15258
rect 12114 15206 17234 15258
rect 17286 15206 17298 15258
rect 17350 15206 17362 15258
rect 17414 15206 17426 15258
rect 17478 15206 17490 15258
rect 17542 15206 22662 15258
rect 22714 15206 22726 15258
rect 22778 15206 22790 15258
rect 22842 15206 22854 15258
rect 22906 15206 22918 15258
rect 22970 15206 22976 15258
rect 1104 15184 22976 15206
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4890 15144 4896 15156
rect 4755 15116 4896 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7098 15144 7104 15156
rect 6972 15116 7104 15144
rect 6972 15104 6978 15116
rect 7098 15104 7104 15116
rect 7156 15144 7162 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7156 15116 7757 15144
rect 7156 15104 7162 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 7745 15107 7803 15113
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 10594 15144 10600 15156
rect 8168 15116 9904 15144
rect 10555 15116 10600 15144
rect 8168 15104 8174 15116
rect 9876 15088 9904 15116
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 4617 15079 4675 15085
rect 4617 15045 4629 15079
rect 4663 15076 4675 15079
rect 5718 15076 5724 15088
rect 4663 15048 5724 15076
rect 4663 15045 4675 15048
rect 4617 15039 4675 15045
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6270 15076 6276 15088
rect 5859 15048 6276 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 9122 15076 9128 15088
rect 7208 15048 9128 15076
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 15008 2283 15011
rect 2498 15008 2504 15020
rect 2271 14980 2504 15008
rect 2271 14977 2283 14980
rect 2225 14971 2283 14977
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 4246 15008 4252 15020
rect 3467 14980 4252 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 5166 14968 5172 15020
rect 5224 15008 5230 15020
rect 5629 15011 5687 15017
rect 5629 15008 5641 15011
rect 5224 14980 5641 15008
rect 5224 14968 5230 14980
rect 5629 14977 5641 14980
rect 5675 14977 5687 15011
rect 5629 14971 5687 14977
rect 6822 14968 6828 15020
rect 6880 15008 6886 15020
rect 7208 15017 7236 15048
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 9858 15076 9864 15088
rect 9771 15048 9864 15076
rect 9858 15036 9864 15048
rect 9916 15036 9922 15088
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 6880 14980 7113 15008
rect 6880 14968 6886 14980
rect 7101 14977 7113 14980
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 15008 7987 15011
rect 8202 15008 8208 15020
rect 7975 14980 8208 15008
rect 7975 14977 7987 14980
rect 7929 14971 7987 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8754 15008 8760 15020
rect 8715 14980 8760 15008
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9582 15008 9588 15020
rect 9079 14980 9588 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 10042 15008 10048 15020
rect 10003 14980 10048 15008
rect 10042 14968 10048 14980
rect 10100 15008 10106 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10100 14980 10517 15008
rect 10100 14968 10106 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10686 15008 10692 15020
rect 10647 14980 10692 15008
rect 10505 14971 10563 14977
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 2314 14940 2320 14952
rect 2275 14912 2320 14940
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2409 14943 2467 14949
rect 2409 14909 2421 14943
rect 2455 14940 2467 14943
rect 2774 14940 2780 14952
rect 2455 14912 2780 14940
rect 2455 14909 2467 14912
rect 2409 14903 2467 14909
rect 2774 14900 2780 14912
rect 2832 14940 2838 14952
rect 2832 14912 3464 14940
rect 2832 14900 2838 14912
rect 3436 14884 3464 14912
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 3697 14943 3755 14949
rect 3568 14912 3613 14940
rect 3568 14900 3574 14912
rect 3697 14909 3709 14943
rect 3743 14940 3755 14943
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 3743 14912 4905 14940
rect 3743 14909 3755 14912
rect 3697 14903 3755 14909
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5074 14940 5080 14952
rect 4939 14912 5080 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7742 14940 7748 14952
rect 7055 14912 7748 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 3418 14832 3424 14884
rect 3476 14832 3482 14884
rect 1857 14807 1915 14813
rect 1857 14773 1869 14807
rect 1903 14804 1915 14807
rect 2130 14804 2136 14816
rect 1903 14776 2136 14804
rect 1903 14773 1915 14776
rect 1857 14767 1915 14773
rect 2130 14764 2136 14776
rect 2188 14764 2194 14816
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3053 14807 3111 14813
rect 3053 14804 3065 14807
rect 3016 14776 3065 14804
rect 3016 14764 3022 14776
rect 3053 14773 3065 14776
rect 3099 14773 3111 14807
rect 3053 14767 3111 14773
rect 3234 14764 3240 14816
rect 3292 14804 3298 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3292 14776 4261 14804
rect 3292 14764 3298 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 4249 14767 4307 14773
rect 4890 14764 4896 14816
rect 4948 14804 4954 14816
rect 5445 14807 5503 14813
rect 5445 14804 5457 14807
rect 4948 14776 5457 14804
rect 4948 14764 4954 14776
rect 5445 14773 5457 14776
rect 5491 14773 5503 14807
rect 5445 14767 5503 14773
rect 6733 14807 6791 14813
rect 6733 14773 6745 14807
rect 6779 14804 6791 14807
rect 6822 14804 6828 14816
rect 6779 14776 6828 14804
rect 6779 14773 6791 14776
rect 6733 14767 6791 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 6932 14804 6960 14903
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 8110 14940 8116 14952
rect 8071 14912 8116 14940
rect 8110 14900 8116 14912
rect 8168 14900 8174 14952
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 9490 14940 9496 14952
rect 9171 14912 9496 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 8938 14872 8944 14884
rect 8899 14844 8944 14872
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 7006 14804 7012 14816
rect 6932 14776 7012 14804
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7558 14764 7564 14816
rect 7616 14804 7622 14816
rect 8849 14807 8907 14813
rect 8849 14804 8861 14807
rect 7616 14776 8861 14804
rect 7616 14764 7622 14776
rect 8849 14773 8861 14776
rect 8895 14804 8907 14807
rect 9398 14804 9404 14816
rect 8895 14776 9404 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 9398 14764 9404 14776
rect 9456 14804 9462 14816
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 9456 14776 9689 14804
rect 9456 14764 9462 14776
rect 9677 14773 9689 14776
rect 9723 14773 9735 14807
rect 9677 14767 9735 14773
rect 1104 14714 22816 14736
rect 1104 14662 3664 14714
rect 3716 14662 3728 14714
rect 3780 14662 3792 14714
rect 3844 14662 3856 14714
rect 3908 14662 3920 14714
rect 3972 14662 9092 14714
rect 9144 14662 9156 14714
rect 9208 14662 9220 14714
rect 9272 14662 9284 14714
rect 9336 14662 9348 14714
rect 9400 14662 14520 14714
rect 14572 14662 14584 14714
rect 14636 14662 14648 14714
rect 14700 14662 14712 14714
rect 14764 14662 14776 14714
rect 14828 14662 19948 14714
rect 20000 14662 20012 14714
rect 20064 14662 20076 14714
rect 20128 14662 20140 14714
rect 20192 14662 20204 14714
rect 20256 14662 22816 14714
rect 1104 14640 22816 14662
rect 2314 14560 2320 14612
rect 2372 14600 2378 14612
rect 4709 14603 4767 14609
rect 4709 14600 4721 14603
rect 2372 14572 4721 14600
rect 2372 14560 2378 14572
rect 4709 14569 4721 14572
rect 4755 14569 4767 14603
rect 4709 14563 4767 14569
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 7800 14572 8493 14600
rect 7800 14560 7806 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 8481 14563 8539 14569
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 8812 14572 9229 14600
rect 8812 14560 8818 14572
rect 9217 14569 9229 14572
rect 9263 14569 9275 14603
rect 9217 14563 9275 14569
rect 9309 14603 9367 14609
rect 9309 14569 9321 14603
rect 9355 14600 9367 14603
rect 9490 14600 9496 14612
rect 9355 14572 9496 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9640 14572 9965 14600
rect 9640 14560 9646 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 2958 14464 2964 14476
rect 2832 14436 2877 14464
rect 2919 14436 2964 14464
rect 2832 14424 2838 14436
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 6730 14464 6736 14476
rect 3068 14436 4476 14464
rect 2038 14396 2044 14408
rect 1999 14368 2044 14396
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 3068 14405 3096 14436
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14365 3111 14399
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3053 14359 3111 14365
rect 3436 14368 3985 14396
rect 2222 14260 2228 14272
rect 2183 14232 2228 14260
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 3436 14269 3464 14368
rect 3973 14365 3985 14368
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 3421 14263 3479 14269
rect 3421 14229 3433 14263
rect 3467 14229 3479 14263
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 3421 14223 3479 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4448 14260 4476 14436
rect 5000 14436 6736 14464
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5000 14405 5028 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7558 14464 7564 14476
rect 6932 14436 7564 14464
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 5350 14396 5356 14408
rect 5311 14368 5356 14396
rect 4985 14359 5043 14365
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 6932 14405 6960 14436
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 8404 14436 9413 14464
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 5592 14368 6837 14396
rect 5592 14356 5598 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 7098 14396 7104 14408
rect 7059 14368 7104 14396
rect 6917 14359 6975 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 5074 14328 5080 14340
rect 5035 14300 5080 14328
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 5195 14331 5253 14337
rect 5195 14328 5207 14331
rect 5184 14297 5207 14328
rect 5241 14297 5253 14331
rect 5184 14291 5253 14297
rect 4890 14260 4896 14272
rect 4448 14232 4896 14260
rect 4890 14220 4896 14232
rect 4948 14260 4954 14272
rect 5184 14260 5212 14291
rect 7006 14288 7012 14340
rect 7064 14328 7070 14340
rect 7208 14328 7236 14359
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8404 14405 8432 14436
rect 9401 14433 9413 14436
rect 9447 14464 9459 14467
rect 10686 14464 10692 14476
rect 9447 14436 10692 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8352 14368 8401 14396
rect 8352 14356 8358 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8662 14396 8668 14408
rect 8619 14368 8668 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8904 14368 9137 14396
rect 8904 14356 8910 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9125 14359 9183 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10042 14356 10048 14408
rect 10100 14396 10106 14408
rect 10100 14368 10193 14396
rect 10100 14356 10106 14368
rect 7064 14300 7236 14328
rect 8680 14328 8708 14356
rect 10060 14328 10088 14356
rect 8680 14300 10088 14328
rect 7064 14288 7070 14300
rect 4948 14232 5212 14260
rect 6641 14263 6699 14269
rect 4948 14220 4954 14232
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 6730 14260 6736 14272
rect 6687 14232 6736 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 1104 14170 22976 14192
rect 1104 14118 6378 14170
rect 6430 14118 6442 14170
rect 6494 14118 6506 14170
rect 6558 14118 6570 14170
rect 6622 14118 6634 14170
rect 6686 14118 11806 14170
rect 11858 14118 11870 14170
rect 11922 14118 11934 14170
rect 11986 14118 11998 14170
rect 12050 14118 12062 14170
rect 12114 14118 17234 14170
rect 17286 14118 17298 14170
rect 17350 14118 17362 14170
rect 17414 14118 17426 14170
rect 17478 14118 17490 14170
rect 17542 14118 22662 14170
rect 22714 14118 22726 14170
rect 22778 14118 22790 14170
rect 22842 14118 22854 14170
rect 22906 14118 22918 14170
rect 22970 14118 22976 14170
rect 1104 14096 22976 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2096 14028 2789 14056
rect 2096 14016 2102 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 3234 14056 3240 14068
rect 3195 14028 3240 14056
rect 2777 14019 2835 14025
rect 3234 14016 3240 14028
rect 3292 14016 3298 14068
rect 7006 13948 7012 14000
rect 7064 13988 7070 14000
rect 8205 13991 8263 13997
rect 8205 13988 8217 13991
rect 7064 13960 8217 13988
rect 7064 13948 7070 13960
rect 8205 13957 8217 13960
rect 8251 13957 8263 13991
rect 8205 13951 8263 13957
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 4246 13920 4252 13932
rect 3191 13892 4252 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 4246 13880 4252 13892
rect 4304 13920 4310 13932
rect 4614 13920 4620 13932
rect 4304 13892 4620 13920
rect 4304 13880 4310 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7098 13920 7104 13932
rect 6871 13892 7104 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8386 13920 8392 13932
rect 8347 13892 8392 13920
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9858 13920 9864 13932
rect 8987 13892 9864 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 10318 13920 10324 13932
rect 10279 13892 10324 13920
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 14274 13920 14280 13932
rect 10551 13892 14280 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 3418 13852 3424 13864
rect 3379 13824 3424 13852
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13852 6607 13855
rect 6730 13852 6736 13864
rect 6595 13824 6736 13852
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8904 13824 9045 13852
rect 8904 13812 8910 13824
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9674 13812 9680 13864
rect 9732 13852 9738 13864
rect 10520 13852 10548 13883
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 9732 13824 10548 13852
rect 9732 13812 9738 13824
rect 6641 13787 6699 13793
rect 6641 13753 6653 13787
rect 6687 13784 6699 13787
rect 7098 13784 7104 13796
rect 6687 13756 7104 13784
rect 6687 13753 6699 13756
rect 6641 13747 6699 13753
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 6730 13716 6736 13728
rect 6691 13688 6736 13716
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 10413 13719 10471 13725
rect 10413 13685 10425 13719
rect 10459 13716 10471 13719
rect 10778 13716 10784 13728
rect 10459 13688 10784 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 11057 13719 11115 13725
rect 11057 13685 11069 13719
rect 11103 13716 11115 13719
rect 11146 13716 11152 13728
rect 11103 13688 11152 13716
rect 11103 13685 11115 13688
rect 11057 13679 11115 13685
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 1104 13626 22816 13648
rect 1104 13574 3664 13626
rect 3716 13574 3728 13626
rect 3780 13574 3792 13626
rect 3844 13574 3856 13626
rect 3908 13574 3920 13626
rect 3972 13574 9092 13626
rect 9144 13574 9156 13626
rect 9208 13574 9220 13626
rect 9272 13574 9284 13626
rect 9336 13574 9348 13626
rect 9400 13574 14520 13626
rect 14572 13574 14584 13626
rect 14636 13574 14648 13626
rect 14700 13574 14712 13626
rect 14764 13574 14776 13626
rect 14828 13574 19948 13626
rect 20000 13574 20012 13626
rect 20064 13574 20076 13626
rect 20128 13574 20140 13626
rect 20192 13574 20204 13626
rect 20256 13574 22816 13626
rect 1104 13552 22816 13574
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 12308 13484 12541 13512
rect 12308 13472 12314 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 4709 13447 4767 13453
rect 4709 13413 4721 13447
rect 4755 13444 4767 13447
rect 5261 13447 5319 13453
rect 5261 13444 5273 13447
rect 4755 13416 5273 13444
rect 4755 13413 4767 13416
rect 4709 13407 4767 13413
rect 5261 13413 5273 13416
rect 5307 13444 5319 13447
rect 5442 13444 5448 13456
rect 5307 13416 5448 13444
rect 5307 13413 5319 13416
rect 5261 13407 5319 13413
rect 2682 13376 2688 13388
rect 2643 13348 2688 13376
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13308 2562 13320
rect 3234 13308 3240 13320
rect 2556 13280 3240 13308
rect 2556 13268 2562 13280
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3602 13268 3608 13320
rect 3660 13308 3666 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3660 13280 3985 13308
rect 3660 13268 3666 13280
rect 3973 13277 3985 13280
rect 4019 13308 4031 13311
rect 4724 13308 4752 13407
rect 5442 13404 5448 13416
rect 5500 13444 5506 13456
rect 5500 13416 8064 13444
rect 5500 13404 5506 13416
rect 7650 13376 7656 13388
rect 4019 13280 4752 13308
rect 5184 13348 7656 13376
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 2593 13243 2651 13249
rect 2593 13209 2605 13243
rect 2639 13240 2651 13243
rect 5184 13240 5212 13348
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 6178 13308 6184 13320
rect 6139 13280 6184 13308
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13308 6423 13311
rect 6822 13308 6828 13320
rect 6411 13280 6828 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 2639 13212 5212 13240
rect 2639 13209 2651 13212
rect 2593 13203 2651 13209
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 7929 13243 7987 13249
rect 7929 13240 7941 13243
rect 6788 13212 7941 13240
rect 6788 13200 6794 13212
rect 7929 13209 7941 13212
rect 7975 13209 7987 13243
rect 8036 13240 8064 13416
rect 8938 13404 8944 13456
rect 8996 13444 9002 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 8996 13416 10425 13444
rect 8996 13404 9002 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 11054 13444 11060 13456
rect 10413 13407 10471 13413
rect 10704 13416 11060 13444
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13376 8263 13379
rect 8846 13376 8852 13388
rect 8251 13348 8852 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 10704 13385 10732 13416
rect 11054 13404 11060 13416
rect 11112 13444 11118 13456
rect 12268 13444 12296 13472
rect 11112 13416 12296 13444
rect 11112 13404 11118 13416
rect 10689 13379 10747 13385
rect 10689 13345 10701 13379
rect 10735 13345 10747 13379
rect 10689 13339 10747 13345
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 12158 13376 12164 13388
rect 12023 13348 12164 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12158 13336 12164 13348
rect 12216 13376 12222 13388
rect 12216 13348 12756 13376
rect 12216 13336 12222 13348
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8294 13308 8300 13320
rect 8159 13280 8300 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 8294 13268 8300 13280
rect 8352 13308 8358 13320
rect 8478 13308 8484 13320
rect 8352 13280 8484 13308
rect 8352 13268 8358 13280
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 9861 13243 9919 13249
rect 9861 13240 9873 13243
rect 8036 13212 9873 13240
rect 7929 13203 7987 13209
rect 9861 13209 9873 13212
rect 9907 13240 9919 13243
rect 10612 13240 10640 13271
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10836 13280 10885 13308
rect 10836 13268 10842 13280
rect 10873 13277 10885 13280
rect 10919 13308 10931 13311
rect 10962 13308 10968 13320
rect 10919 13280 10968 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 12342 13308 12348 13320
rect 11931 13280 12348 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 11146 13240 11152 13252
rect 9907 13212 11152 13240
rect 9907 13209 9919 13212
rect 9861 13203 9919 13209
rect 10796 13184 10824 13212
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 11808 13240 11836 13271
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12728 13317 12756 13348
rect 12535 13311 12593 13317
rect 12535 13277 12547 13311
rect 12581 13277 12593 13311
rect 12535 13271 12593 13277
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 13262 13308 13268 13320
rect 12759 13280 13268 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 12434 13240 12440 13252
rect 11808 13212 12440 13240
rect 12434 13200 12440 13212
rect 12492 13240 12498 13252
rect 12544 13240 12572 13271
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 14182 13308 14188 13320
rect 13495 13280 14188 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 13357 13243 13415 13249
rect 13357 13240 13369 13243
rect 12492 13212 13369 13240
rect 12492 13200 12498 13212
rect 13357 13209 13369 13212
rect 13403 13209 13415 13243
rect 13357 13203 13415 13209
rect 2130 13172 2136 13184
rect 2091 13144 2136 13172
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 2832 13144 3341 13172
rect 2832 13132 2838 13144
rect 3329 13141 3341 13144
rect 3375 13141 3387 13175
rect 3329 13135 3387 13141
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 3970 13172 3976 13184
rect 3476 13144 3976 13172
rect 3476 13132 3482 13144
rect 3970 13132 3976 13144
rect 4028 13172 4034 13184
rect 4065 13175 4123 13181
rect 4065 13172 4077 13175
rect 4028 13144 4077 13172
rect 4028 13132 4034 13144
rect 4065 13141 4077 13144
rect 4111 13141 4123 13175
rect 4065 13135 4123 13141
rect 6273 13175 6331 13181
rect 6273 13141 6285 13175
rect 6319 13172 6331 13175
rect 7466 13172 7472 13184
rect 6319 13144 7472 13172
rect 6319 13141 6331 13144
rect 6273 13135 6331 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 8573 13175 8631 13181
rect 8573 13172 8585 13175
rect 8444 13144 8585 13172
rect 8444 13132 8450 13144
rect 8573 13141 8585 13144
rect 8619 13172 8631 13175
rect 9582 13172 9588 13184
rect 8619 13144 9588 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10778 13132 10784 13184
rect 10836 13132 10842 13184
rect 11514 13172 11520 13184
rect 11475 13144 11520 13172
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 1104 13082 22976 13104
rect 1104 13030 6378 13082
rect 6430 13030 6442 13082
rect 6494 13030 6506 13082
rect 6558 13030 6570 13082
rect 6622 13030 6634 13082
rect 6686 13030 11806 13082
rect 11858 13030 11870 13082
rect 11922 13030 11934 13082
rect 11986 13030 11998 13082
rect 12050 13030 12062 13082
rect 12114 13030 17234 13082
rect 17286 13030 17298 13082
rect 17350 13030 17362 13082
rect 17414 13030 17426 13082
rect 17478 13030 17490 13082
rect 17542 13030 22662 13082
rect 22714 13030 22726 13082
rect 22778 13030 22790 13082
rect 22842 13030 22854 13082
rect 22906 13030 22918 13082
rect 22970 13030 22976 13082
rect 1104 13008 22976 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 5074 12968 5080 12980
rect 2746 12940 5080 12968
rect 2746 12900 2774 12940
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 5215 12940 6561 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 6917 12971 6975 12977
rect 6917 12968 6929 12971
rect 6880 12940 6929 12968
rect 6880 12928 6886 12940
rect 6917 12937 6929 12940
rect 6963 12937 6975 12971
rect 6917 12931 6975 12937
rect 7009 12971 7067 12977
rect 7009 12937 7021 12971
rect 7055 12968 7067 12971
rect 7098 12968 7104 12980
rect 7055 12940 7104 12968
rect 7055 12937 7067 12940
rect 7009 12931 7067 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7929 12971 7987 12977
rect 7929 12968 7941 12971
rect 7800 12940 7941 12968
rect 7800 12928 7806 12940
rect 7929 12937 7941 12940
rect 7975 12968 7987 12971
rect 9674 12968 9680 12980
rect 7975 12940 9680 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 11054 12968 11060 12980
rect 10244 12940 11060 12968
rect 2056 12872 2774 12900
rect 3145 12903 3203 12909
rect 2056 12841 2084 12872
rect 3145 12869 3157 12903
rect 3191 12900 3203 12903
rect 3973 12903 4031 12909
rect 3191 12872 3924 12900
rect 3191 12869 3203 12872
rect 3145 12863 3203 12869
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 2866 12832 2872 12844
rect 2827 12804 2872 12832
rect 2041 12795 2099 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3016 12804 3061 12832
rect 3016 12792 3022 12804
rect 2225 12767 2283 12773
rect 2225 12764 2237 12767
rect 2056 12736 2237 12764
rect 2056 12708 2084 12736
rect 2225 12733 2237 12736
rect 2271 12733 2283 12767
rect 2225 12727 2283 12733
rect 2314 12724 2320 12776
rect 2372 12764 2378 12776
rect 2682 12764 2688 12776
rect 2372 12736 2688 12764
rect 2372 12724 2378 12736
rect 2682 12724 2688 12736
rect 2740 12764 2746 12776
rect 3252 12764 3280 12872
rect 3602 12832 3608 12844
rect 3563 12804 3608 12832
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 3896 12841 3924 12872
rect 3973 12869 3985 12903
rect 4019 12900 4031 12903
rect 6730 12900 6736 12912
rect 4019 12872 6736 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 9766 12900 9772 12912
rect 6932 12872 9772 12900
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 2740 12736 3280 12764
rect 2740 12724 2746 12736
rect 2038 12656 2044 12708
rect 2096 12656 2102 12708
rect 3145 12699 3203 12705
rect 3145 12665 3157 12699
rect 3191 12696 3203 12699
rect 3712 12696 3740 12795
rect 3896 12764 3924 12795
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 5077 12835 5135 12841
rect 4120 12804 4165 12832
rect 4120 12792 4126 12804
rect 5077 12801 5089 12835
rect 5123 12832 5135 12835
rect 5534 12832 5540 12844
rect 5123 12804 5540 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 5718 12832 5724 12844
rect 5592 12804 5724 12832
rect 5592 12792 5598 12804
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 4430 12764 4436 12776
rect 3896 12736 4436 12764
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 4540 12736 5273 12764
rect 3191 12668 3740 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 4540 12696 4568 12736
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 6932 12764 6960 12872
rect 9766 12860 9772 12872
rect 9824 12900 9830 12912
rect 9824 12872 9904 12900
rect 9824 12860 9830 12872
rect 9876 12841 9904 12872
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 5261 12727 5319 12733
rect 6656 12736 6960 12764
rect 7024 12804 7941 12832
rect 4028 12668 4568 12696
rect 4028 12656 4034 12668
rect 5074 12656 5080 12708
rect 5132 12696 5138 12708
rect 6656 12696 6684 12736
rect 5132 12668 6684 12696
rect 5132 12656 5138 12668
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7024 12696 7052 12804
rect 7929 12801 7941 12804
rect 7975 12832 7987 12835
rect 9217 12835 9275 12841
rect 7975 12804 8156 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 6788 12668 7052 12696
rect 6788 12656 6794 12668
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4580 12600 4721 12628
rect 4580 12588 4586 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 4709 12591 4767 12597
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 6178 12628 6184 12640
rect 5224 12600 6184 12628
rect 5224 12588 5230 12600
rect 6178 12588 6184 12600
rect 6236 12628 6242 12640
rect 7208 12628 7236 12727
rect 8128 12696 8156 12804
rect 9217 12801 9229 12835
rect 9263 12832 9275 12835
rect 9677 12835 9735 12841
rect 9677 12832 9689 12835
rect 9263 12804 9689 12832
rect 9263 12801 9275 12804
rect 9217 12795 9275 12801
rect 9677 12801 9689 12804
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10244 12832 10272 12940
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 12618 12968 12624 12980
rect 12084 12940 12624 12968
rect 10502 12900 10508 12912
rect 10336 12872 10508 12900
rect 10336 12841 10364 12872
rect 10502 12860 10508 12872
rect 10560 12900 10566 12912
rect 10560 12872 10916 12900
rect 10560 12860 10566 12872
rect 10888 12844 10916 12872
rect 10183 12804 10272 12832
rect 10321 12835 10379 12841
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10321 12795 10379 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10928 12804 10977 12832
rect 10928 12792 10934 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11698 12832 11704 12844
rect 11112 12804 11704 12832
rect 11112 12792 11118 12804
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12084 12841 12112 12940
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12968 12771 12971
rect 12759 12940 16574 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 12434 12900 12440 12912
rect 12395 12872 12440 12900
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 16546 12900 16574 12940
rect 16942 12900 16948 12912
rect 16546 12872 16948 12900
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12158 12792 12164 12844
rect 12216 12832 12222 12844
rect 12342 12832 12348 12844
rect 12216 12804 12261 12832
rect 12303 12804 12348 12832
rect 12216 12792 12222 12804
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12801 13599 12835
rect 14182 12832 14188 12844
rect 14143 12804 14188 12832
rect 13541 12795 13599 12801
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8352 12736 8953 12764
rect 8352 12724 8358 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9125 12767 9183 12773
rect 9125 12733 9137 12767
rect 9171 12764 9183 12767
rect 11514 12764 11520 12776
rect 9171 12736 11520 12764
rect 9171 12733 9183 12736
rect 9125 12727 9183 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11716 12764 11744 12792
rect 12544 12764 12572 12795
rect 11716 12736 12572 12764
rect 9858 12696 9864 12708
rect 8128 12668 9864 12696
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 11057 12699 11115 12705
rect 11057 12665 11069 12699
rect 11103 12696 11115 12699
rect 11146 12696 11152 12708
rect 11103 12668 11152 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 11146 12656 11152 12668
rect 11204 12696 11210 12708
rect 13446 12696 13452 12708
rect 11204 12668 13452 12696
rect 11204 12656 11210 12668
rect 13446 12656 13452 12668
rect 13504 12696 13510 12708
rect 13556 12696 13584 12795
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 14332 12804 14381 12832
rect 14332 12792 14338 12804
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 13725 12767 13783 12773
rect 13725 12733 13737 12767
rect 13771 12764 13783 12767
rect 13771 12736 14320 12764
rect 13771 12733 13783 12736
rect 13725 12727 13783 12733
rect 13504 12668 13584 12696
rect 13504 12656 13510 12668
rect 6236 12600 7236 12628
rect 9217 12631 9275 12637
rect 6236 12588 6242 12600
rect 9217 12597 9229 12631
rect 9263 12628 9275 12631
rect 9490 12628 9496 12640
rect 9263 12600 9496 12628
rect 9263 12597 9275 12600
rect 9217 12591 9275 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 14292 12637 14320 12736
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 9732 12600 13369 12628
rect 9732 12588 9738 12600
rect 13357 12597 13369 12600
rect 13403 12597 13415 12631
rect 13357 12591 13415 12597
rect 14277 12631 14335 12637
rect 14277 12597 14289 12631
rect 14323 12628 14335 12631
rect 14366 12628 14372 12640
rect 14323 12600 14372 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 1104 12538 22816 12560
rect 1104 12486 3664 12538
rect 3716 12486 3728 12538
rect 3780 12486 3792 12538
rect 3844 12486 3856 12538
rect 3908 12486 3920 12538
rect 3972 12486 9092 12538
rect 9144 12486 9156 12538
rect 9208 12486 9220 12538
rect 9272 12486 9284 12538
rect 9336 12486 9348 12538
rect 9400 12486 14520 12538
rect 14572 12486 14584 12538
rect 14636 12486 14648 12538
rect 14700 12486 14712 12538
rect 14764 12486 14776 12538
rect 14828 12486 19948 12538
rect 20000 12486 20012 12538
rect 20064 12486 20076 12538
rect 20128 12486 20140 12538
rect 20192 12486 20204 12538
rect 20256 12486 22816 12538
rect 1104 12464 22816 12486
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 3016 12396 3433 12424
rect 3016 12384 3022 12396
rect 3421 12393 3433 12396
rect 3467 12424 3479 12427
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3467 12396 4077 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 4065 12387 4123 12393
rect 4430 12384 4436 12436
rect 4488 12424 4494 12436
rect 5166 12424 5172 12436
rect 4488 12396 5172 12424
rect 4488 12384 4494 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5350 12384 5356 12436
rect 5408 12424 5414 12436
rect 7742 12424 7748 12436
rect 5408 12396 7748 12424
rect 5408 12384 5414 12396
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 8904 12396 9597 12424
rect 8904 12384 8910 12396
rect 9585 12393 9597 12396
rect 9631 12424 9643 12427
rect 9674 12424 9680 12436
rect 9631 12396 9680 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10502 12424 10508 12436
rect 10463 12396 10508 12424
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12400 12396 13093 12424
rect 12400 12384 12406 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 12529 12359 12587 12365
rect 11020 12328 12434 12356
rect 11020 12316 11026 12328
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12257 2007 12291
rect 2130 12288 2136 12300
rect 2091 12260 2136 12288
rect 1949 12251 2007 12257
rect 1964 12220 1992 12251
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12288 4399 12291
rect 4614 12288 4620 12300
rect 4387 12260 4620 12288
rect 4387 12257 4399 12260
rect 4341 12251 4399 12257
rect 4614 12248 4620 12260
rect 4672 12288 4678 12300
rect 4890 12288 4896 12300
rect 4672 12260 4896 12288
rect 4672 12248 4678 12260
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 11146 12288 11152 12300
rect 11107 12260 11152 12288
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 12406 12288 12434 12328
rect 12529 12325 12541 12359
rect 12575 12356 12587 12359
rect 16206 12356 16212 12368
rect 12575 12328 16212 12356
rect 12575 12325 12587 12328
rect 12529 12319 12587 12325
rect 16206 12316 16212 12328
rect 16264 12316 16270 12368
rect 12989 12291 13047 12297
rect 12406 12260 12848 12288
rect 1964 12192 2176 12220
rect 2148 12164 2176 12192
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3234 12220 3240 12232
rect 3016 12192 3240 12220
rect 3016 12180 3022 12192
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4706 12220 4712 12232
rect 4479 12192 4712 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5350 12220 5356 12232
rect 5311 12192 5356 12220
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 2130 12112 2136 12164
rect 2188 12112 2194 12164
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 2682 12152 2688 12164
rect 2271 12124 2688 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 2682 12112 2688 12124
rect 2740 12152 2746 12164
rect 3053 12155 3111 12161
rect 3053 12152 3065 12155
rect 2740 12124 3065 12152
rect 2740 12112 2746 12124
rect 3053 12121 3065 12124
rect 3099 12121 3111 12155
rect 3053 12115 3111 12121
rect 3973 12155 4031 12161
rect 3973 12121 3985 12155
rect 4019 12152 4031 12155
rect 4338 12152 4344 12164
rect 4019 12124 4344 12152
rect 4019 12121 4031 12124
rect 3973 12115 4031 12121
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 2590 12084 2596 12096
rect 2551 12056 2596 12084
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 4617 12087 4675 12093
rect 4617 12053 4629 12087
rect 4663 12084 4675 12087
rect 5552 12084 5580 12183
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5902 12220 5908 12232
rect 5684 12192 5908 12220
rect 5684 12180 5690 12192
rect 5902 12180 5908 12192
rect 5960 12220 5966 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5960 12192 6009 12220
rect 5960 12180 5966 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 6144 12192 6377 12220
rect 6144 12180 6150 12192
rect 6365 12189 6377 12192
rect 6411 12220 6423 12223
rect 6914 12220 6920 12232
rect 6411 12192 6920 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6914 12180 6920 12192
rect 6972 12220 6978 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6972 12192 7297 12220
rect 6972 12180 6978 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 7285 12183 7343 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7650 12220 7656 12232
rect 7611 12192 7656 12220
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 8294 12220 8300 12232
rect 7944 12192 8300 12220
rect 7006 12112 7012 12164
rect 7064 12152 7070 12164
rect 7377 12155 7435 12161
rect 7377 12152 7389 12155
rect 7064 12124 7389 12152
rect 7064 12112 7070 12124
rect 7377 12121 7389 12124
rect 7423 12152 7435 12155
rect 7944 12152 7972 12192
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8570 12220 8576 12232
rect 8435 12192 8576 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8570 12180 8576 12192
rect 8628 12220 8634 12232
rect 8938 12220 8944 12232
rect 8628 12192 8944 12220
rect 8628 12180 8634 12192
rect 8938 12180 8944 12192
rect 8996 12220 9002 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8996 12192 9321 12220
rect 8996 12180 9002 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9677 12223 9735 12229
rect 9456 12192 9501 12220
rect 9456 12180 9462 12192
rect 9677 12189 9689 12223
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 7423 12124 7972 12152
rect 7423 12121 7435 12124
rect 7377 12115 7435 12121
rect 8018 12112 8024 12164
rect 8076 12152 8082 12164
rect 9692 12152 9720 12183
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 9916 12192 10333 12220
rect 9916 12180 9922 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10321 12183 10379 12189
rect 8076 12124 9720 12152
rect 10336 12152 10364 12183
rect 10502 12180 10508 12192
rect 10560 12220 10566 12232
rect 12342 12220 12348 12232
rect 10560 12192 12348 12220
rect 10560 12180 10566 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12710 12220 12716 12232
rect 12671 12192 12716 12220
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 12434 12152 12440 12164
rect 10336 12124 12440 12152
rect 8076 12112 8082 12124
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 12820 12161 12848 12260
rect 12989 12257 13001 12291
rect 13035 12288 13047 12291
rect 14274 12288 14280 12300
rect 13035 12260 14136 12288
rect 14235 12260 14280 12288
rect 13035 12257 13047 12260
rect 12989 12251 13047 12257
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 14108 12220 14136 12260
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 14366 12248 14372 12300
rect 14424 12288 14430 12300
rect 15010 12288 15016 12300
rect 14424 12260 15016 12288
rect 14424 12248 14430 12260
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 14384 12220 14412 12248
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14108 12192 14565 12220
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14734 12220 14740 12232
rect 14695 12192 14740 12220
rect 14553 12183 14611 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 12805 12155 12863 12161
rect 12805 12121 12817 12155
rect 12851 12121 12863 12155
rect 12805 12115 12863 12121
rect 13906 12112 13912 12164
rect 13964 12152 13970 12164
rect 14415 12155 14473 12161
rect 14415 12152 14427 12155
rect 13964 12124 14427 12152
rect 13964 12112 13970 12124
rect 14415 12121 14427 12124
rect 14461 12121 14473 12155
rect 14415 12115 14473 12121
rect 14645 12155 14703 12161
rect 14645 12121 14657 12155
rect 14691 12121 14703 12155
rect 14645 12115 14703 12121
rect 4663 12056 5580 12084
rect 4663 12053 4675 12056
rect 4617 12047 4675 12053
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 5776 12056 7113 12084
rect 5776 12044 5782 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7800 12056 8217 12084
rect 7800 12044 7806 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8205 12047 8263 12053
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8812 12056 9137 12084
rect 8812 12044 8818 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 11238 12084 11244 12096
rect 11199 12056 11244 12084
rect 9125 12047 9183 12053
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11698 12084 11704 12096
rect 11388 12056 11433 12084
rect 11659 12056 11704 12084
rect 11388 12044 11394 12056
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 14660 12084 14688 12115
rect 14918 12084 14924 12096
rect 14332 12056 14688 12084
rect 14879 12056 14924 12084
rect 14332 12044 14338 12056
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 1104 11994 22976 12016
rect 1104 11942 6378 11994
rect 6430 11942 6442 11994
rect 6494 11942 6506 11994
rect 6558 11942 6570 11994
rect 6622 11942 6634 11994
rect 6686 11942 11806 11994
rect 11858 11942 11870 11994
rect 11922 11942 11934 11994
rect 11986 11942 11998 11994
rect 12050 11942 12062 11994
rect 12114 11942 17234 11994
rect 17286 11942 17298 11994
rect 17350 11942 17362 11994
rect 17414 11942 17426 11994
rect 17478 11942 17490 11994
rect 17542 11942 22662 11994
rect 22714 11942 22726 11994
rect 22778 11942 22790 11994
rect 22842 11942 22854 11994
rect 22906 11942 22918 11994
rect 22970 11942 22976 11994
rect 1104 11920 22976 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 4246 11880 4252 11892
rect 2188 11852 3372 11880
rect 4207 11852 4252 11880
rect 2188 11840 2194 11852
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2038 11744 2044 11756
rect 1995 11716 2044 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2240 11685 2268 11852
rect 3344 11756 3372 11852
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 7650 11880 7656 11892
rect 5675 11852 7656 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8941 11883 8999 11889
rect 8941 11849 8953 11883
rect 8987 11849 8999 11883
rect 11054 11880 11060 11892
rect 11015 11852 11060 11880
rect 8941 11843 8999 11849
rect 7466 11772 7472 11824
rect 7524 11812 7530 11824
rect 8018 11812 8024 11824
rect 7524 11784 8024 11812
rect 7524 11772 7530 11784
rect 8018 11772 8024 11784
rect 8076 11812 8082 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 8076 11784 8309 11812
rect 8076 11772 8082 11784
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 8956 11812 8984 11843
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 11296 11852 11713 11880
rect 11296 11840 11302 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 11701 11843 11759 11849
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14182 11880 14188 11892
rect 14139 11852 14188 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 14553 11883 14611 11889
rect 14553 11849 14565 11883
rect 14599 11880 14611 11883
rect 14734 11880 14740 11892
rect 14599 11852 14740 11880
rect 14599 11849 14611 11852
rect 14553 11843 14611 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 10318 11812 10324 11824
rect 8956 11784 10324 11812
rect 8297 11775 8355 11781
rect 10318 11772 10324 11784
rect 10376 11812 10382 11824
rect 10376 11784 11008 11812
rect 10376 11772 10382 11784
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11744 2743 11747
rect 2774 11744 2780 11756
rect 2731 11716 2780 11744
rect 2731 11713 2743 11716
rect 2685 11707 2743 11713
rect 2774 11704 2780 11716
rect 2832 11704 2838 11756
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 4062 11744 4068 11756
rect 3384 11716 4068 11744
rect 3384 11704 3390 11716
rect 4062 11704 4068 11716
rect 4120 11744 4126 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 4120 11716 5457 11744
rect 4120 11704 4126 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 8202 11744 8208 11756
rect 7147 11716 8208 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 10980 11753 11008 11784
rect 8757 11747 8815 11753
rect 8757 11744 8769 11747
rect 8444 11716 8769 11744
rect 8444 11704 8450 11716
rect 8757 11713 8769 11716
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11645 2283 11679
rect 2225 11639 2283 11645
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 5169 11679 5227 11685
rect 3927 11648 5120 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2314 11608 2320 11620
rect 2087 11580 2320 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 3804 11608 3832 11639
rect 4338 11608 4344 11620
rect 2915 11580 3740 11608
rect 3804 11580 4344 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2188 11512 2233 11540
rect 2188 11500 2194 11512
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 3605 11543 3663 11549
rect 3605 11540 3617 11543
rect 3568 11512 3617 11540
rect 3568 11500 3574 11512
rect 3605 11509 3617 11512
rect 3651 11509 3663 11543
rect 3712 11540 3740 11580
rect 4338 11568 4344 11580
rect 4396 11608 4402 11620
rect 5092 11608 5120 11648
rect 5169 11645 5181 11679
rect 5215 11676 5227 11679
rect 6270 11676 6276 11688
rect 5215 11648 6276 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 6512 11648 7205 11676
rect 6512 11636 6518 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 8938 11676 8944 11688
rect 8711 11648 8944 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 7006 11608 7012 11620
rect 4396 11580 4844 11608
rect 5092 11580 7012 11608
rect 4396 11568 4402 11580
rect 4816 11552 4844 11580
rect 7006 11568 7012 11580
rect 7064 11568 7070 11620
rect 7392 11608 7420 11639
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9398 11676 9404 11688
rect 9359 11648 9404 11676
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 8846 11608 8852 11620
rect 7392 11580 8852 11608
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 8956 11608 8984 11636
rect 9692 11608 9720 11639
rect 8956 11580 9720 11608
rect 4246 11540 4252 11552
rect 3712 11512 4252 11540
rect 3605 11503 3663 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 4856 11512 5273 11540
rect 4856 11500 4862 11512
rect 5261 11509 5273 11512
rect 5307 11509 5319 11543
rect 5261 11503 5319 11509
rect 5810 11500 5816 11552
rect 5868 11540 5874 11552
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 5868 11512 6745 11540
rect 5868 11500 5874 11512
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 6733 11503 6791 11509
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8260 11512 8769 11540
rect 8260 11500 8266 11512
rect 8757 11509 8769 11512
rect 8803 11540 8815 11543
rect 9784 11540 9812 11707
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11664 11716 11897 11744
rect 11664 11704 11670 11716
rect 11885 11713 11897 11716
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12158 11744 12164 11756
rect 12023 11716 12164 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12434 11744 12440 11756
rect 12299 11716 12440 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12434 11704 12440 11716
rect 12492 11744 12498 11756
rect 13262 11744 13268 11756
rect 12492 11716 13268 11744
rect 12492 11704 12498 11716
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 14366 11744 14372 11756
rect 13955 11716 14372 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 13556 11676 13584 11707
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15194 11744 15200 11756
rect 14967 11716 15200 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 12124 11648 13584 11676
rect 12124 11636 12130 11648
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14752 11676 14780 11707
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 14240 11648 14780 11676
rect 14240 11636 14246 11648
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 11388 11580 12434 11608
rect 11388 11568 11394 11580
rect 8803 11512 9812 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 12066 11540 12072 11552
rect 11204 11512 12072 11540
rect 11204 11500 11210 11512
rect 12066 11500 12072 11512
rect 12124 11540 12130 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 12124 11512 12173 11540
rect 12124 11500 12130 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12406 11540 12434 11580
rect 13906 11540 13912 11552
rect 12406 11512 13912 11540
rect 12161 11503 12219 11509
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 1104 11450 22816 11472
rect 1104 11398 3664 11450
rect 3716 11398 3728 11450
rect 3780 11398 3792 11450
rect 3844 11398 3856 11450
rect 3908 11398 3920 11450
rect 3972 11398 9092 11450
rect 9144 11398 9156 11450
rect 9208 11398 9220 11450
rect 9272 11398 9284 11450
rect 9336 11398 9348 11450
rect 9400 11398 14520 11450
rect 14572 11398 14584 11450
rect 14636 11398 14648 11450
rect 14700 11398 14712 11450
rect 14764 11398 14776 11450
rect 14828 11398 19948 11450
rect 20000 11398 20012 11450
rect 20064 11398 20076 11450
rect 20128 11398 20140 11450
rect 20192 11398 20204 11450
rect 20256 11398 22816 11450
rect 1104 11376 22816 11398
rect 2866 11296 2872 11348
rect 2924 11336 2930 11348
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2924 11308 2973 11336
rect 2924 11296 2930 11308
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 2961 11299 3019 11305
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 5442 11336 5448 11348
rect 4304 11308 5448 11336
rect 4304 11296 4310 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11756 11308 12020 11336
rect 11756 11296 11762 11308
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 1854 11268 1860 11280
rect 1811 11240 1860 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 1854 11228 1860 11240
rect 1912 11228 1918 11280
rect 8297 11271 8355 11277
rect 8297 11268 8309 11271
rect 7300 11240 8309 11268
rect 2130 11200 2136 11212
rect 1780 11172 2136 11200
rect 1780 11141 1808 11172
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 7300 11209 7328 11240
rect 8297 11237 8309 11240
rect 8343 11237 8355 11271
rect 8297 11231 8355 11237
rect 11793 11271 11851 11277
rect 11793 11237 11805 11271
rect 11839 11237 11851 11271
rect 11793 11231 11851 11237
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 2648 11172 5212 11200
rect 2648 11160 2654 11172
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11101 1823 11135
rect 1765 11095 1823 11101
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2314 11132 2320 11144
rect 2087 11104 2320 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 4522 11132 4528 11144
rect 4483 11104 4528 11132
rect 3053 11095 3111 11101
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 2130 11064 2136 11076
rect 1995 11036 2136 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 2130 11024 2136 11036
rect 2188 11024 2194 11076
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 3068 11064 3096 11095
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 5184 11141 5212 11172
rect 6656 11172 7297 11200
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5810 11132 5816 11144
rect 5771 11104 5816 11132
rect 5169 11095 5227 11101
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 6656 11141 6684 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7742 11200 7748 11212
rect 7703 11172 7748 11200
rect 7285 11163 7343 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 6328 11104 6469 11132
rect 6328 11092 6334 11104
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 8386 11132 8392 11144
rect 7423 11104 8248 11132
rect 8347 11104 8392 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 2740 11036 3096 11064
rect 6472 11064 6500 11095
rect 6730 11064 6736 11076
rect 6472 11036 6736 11064
rect 2740 11024 2746 11036
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 7653 11067 7711 11073
rect 7653 11064 7665 11067
rect 7524 11036 7665 11064
rect 7524 11024 7530 11036
rect 7653 11033 7665 11036
rect 7699 11033 7711 11067
rect 8220 11064 8248 11104
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9732 11104 9965 11132
rect 9732 11092 9738 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10220 11135 10278 11141
rect 10220 11101 10232 11135
rect 10266 11132 10278 11135
rect 11808 11132 11836 11231
rect 11992 11141 12020 11308
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 14332 11308 14381 11336
rect 14332 11296 14338 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 15194 11200 15200 11212
rect 14292 11172 15200 11200
rect 14292 11141 14320 11172
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 10266 11104 11836 11132
rect 11977 11135 12035 11141
rect 10266 11101 10278 11104
rect 10220 11095 10278 11101
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 8846 11064 8852 11076
rect 8220 11036 8852 11064
rect 7653 11027 7711 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 11606 11024 11612 11076
rect 11664 11064 11670 11076
rect 14182 11064 14188 11076
rect 11664 11036 14188 11064
rect 11664 11024 11670 11036
rect 14182 11024 14188 11036
rect 14240 11064 14246 11076
rect 14476 11064 14504 11095
rect 14240 11036 14504 11064
rect 14240 11024 14246 11036
rect 4338 10996 4344 11008
rect 4299 10968 4344 10996
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 4985 10999 5043 11005
rect 4985 10996 4997 10999
rect 4488 10968 4997 10996
rect 4488 10956 4494 10968
rect 4985 10965 4997 10968
rect 5031 10965 5043 10999
rect 5994 10996 6000 11008
rect 5955 10968 6000 10996
rect 4985 10959 5043 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 7098 10996 7104 11008
rect 7059 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 1104 10906 22976 10928
rect 1104 10854 6378 10906
rect 6430 10854 6442 10906
rect 6494 10854 6506 10906
rect 6558 10854 6570 10906
rect 6622 10854 6634 10906
rect 6686 10854 11806 10906
rect 11858 10854 11870 10906
rect 11922 10854 11934 10906
rect 11986 10854 11998 10906
rect 12050 10854 12062 10906
rect 12114 10854 17234 10906
rect 17286 10854 17298 10906
rect 17350 10854 17362 10906
rect 17414 10854 17426 10906
rect 17478 10854 17490 10906
rect 17542 10854 22662 10906
rect 22714 10854 22726 10906
rect 22778 10854 22790 10906
rect 22842 10854 22854 10906
rect 22906 10854 22918 10906
rect 22970 10854 22976 10906
rect 1104 10832 22976 10854
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 2188 10764 2973 10792
rect 2188 10752 2194 10764
rect 2961 10761 2973 10764
rect 3007 10761 3019 10795
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 2961 10755 3019 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8386 10792 8392 10804
rect 7975 10764 8392 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 11146 10792 11152 10804
rect 11107 10764 11152 10792
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10761 11943 10795
rect 11885 10755 11943 10761
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13814 10792 13820 10804
rect 13587 10764 13820 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 3510 10684 3516 10736
rect 3568 10724 3574 10736
rect 3666 10727 3724 10733
rect 3666 10724 3678 10727
rect 3568 10696 3678 10724
rect 3568 10684 3574 10696
rect 3666 10693 3678 10696
rect 3712 10693 3724 10727
rect 3666 10687 3724 10693
rect 6816 10727 6874 10733
rect 6816 10693 6828 10727
rect 6862 10724 6874 10727
rect 7098 10724 7104 10736
rect 6862 10696 7104 10724
rect 6862 10693 6874 10696
rect 6816 10687 6874 10693
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 10036 10727 10094 10733
rect 8260 10696 8708 10724
rect 8260 10684 8266 10696
rect 1854 10665 1860 10668
rect 1848 10656 1860 10665
rect 1815 10628 1860 10656
rect 1848 10619 1860 10628
rect 1854 10616 1860 10619
rect 1912 10616 1918 10668
rect 8570 10656 8576 10668
rect 8531 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8680 10665 8708 10696
rect 10036 10693 10048 10727
rect 10082 10724 10094 10727
rect 11900 10724 11928 10755
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 14366 10752 14372 10804
rect 14424 10792 14430 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 14424 10764 14749 10792
rect 14424 10752 14430 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 14737 10755 14795 10761
rect 10082 10696 11928 10724
rect 13633 10727 13691 10733
rect 10082 10693 10094 10696
rect 10036 10687 10094 10693
rect 13633 10693 13645 10727
rect 13679 10724 13691 10727
rect 14918 10724 14924 10736
rect 13679 10696 14924 10724
rect 13679 10693 13691 10696
rect 13633 10687 13691 10693
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 15010 10684 15016 10736
rect 15068 10724 15074 10736
rect 15068 10696 15424 10724
rect 15068 10684 15074 10696
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8938 10656 8944 10668
rect 8899 10628 8944 10656
rect 8665 10619 8723 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 12066 10656 12072 10668
rect 12027 10628 12072 10656
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 12713 10659 12771 10665
rect 12713 10625 12725 10659
rect 12759 10656 12771 10659
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 12759 10628 13216 10656
rect 12759 10625 12771 10628
rect 12713 10619 12771 10625
rect 1578 10588 1584 10600
rect 1539 10560 1584 10588
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 3418 10588 3424 10600
rect 3379 10560 3424 10588
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6236 10560 6561 10588
rect 6236 10548 6242 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 8846 10588 8852 10600
rect 8807 10560 8852 10588
rect 6549 10551 6607 10557
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9732 10560 9781 10588
rect 9732 10548 9738 10560
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 13188 10529 13216 10628
rect 13648 10628 14381 10656
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13648 10588 13676 10628
rect 14369 10625 14381 10628
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10625 14611 10659
rect 15194 10656 15200 10668
rect 15155 10628 15200 10656
rect 14553 10619 14611 10625
rect 13412 10560 13676 10588
rect 13725 10591 13783 10597
rect 13412 10548 13418 10560
rect 13725 10557 13737 10591
rect 13771 10557 13783 10591
rect 13725 10551 13783 10557
rect 13173 10523 13231 10529
rect 13173 10489 13185 10523
rect 13219 10489 13231 10523
rect 13173 10483 13231 10489
rect 13446 10480 13452 10532
rect 13504 10520 13510 10532
rect 13740 10520 13768 10551
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14568 10588 14596 10619
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15396 10665 15424 10696
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 13872 10560 14596 10588
rect 13872 10548 13878 10560
rect 13504 10492 13768 10520
rect 13504 10480 13510 10492
rect 8386 10452 8392 10464
rect 8347 10424 8392 10452
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 14918 10412 14924 10464
rect 14976 10452 14982 10464
rect 15289 10455 15347 10461
rect 15289 10452 15301 10455
rect 14976 10424 15301 10452
rect 14976 10412 14982 10424
rect 15289 10421 15301 10424
rect 15335 10421 15347 10455
rect 15289 10415 15347 10421
rect 1104 10362 22816 10384
rect 1104 10310 3664 10362
rect 3716 10310 3728 10362
rect 3780 10310 3792 10362
rect 3844 10310 3856 10362
rect 3908 10310 3920 10362
rect 3972 10310 9092 10362
rect 9144 10310 9156 10362
rect 9208 10310 9220 10362
rect 9272 10310 9284 10362
rect 9336 10310 9348 10362
rect 9400 10310 14520 10362
rect 14572 10310 14584 10362
rect 14636 10310 14648 10362
rect 14700 10310 14712 10362
rect 14764 10310 14776 10362
rect 14828 10310 19948 10362
rect 20000 10310 20012 10362
rect 20064 10310 20076 10362
rect 20128 10310 20140 10362
rect 20192 10310 20204 10362
rect 20256 10310 22816 10362
rect 1104 10288 22816 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2682 10248 2688 10260
rect 1627 10220 2688 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 6086 10248 6092 10260
rect 5767 10220 6092 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 8202 10248 8208 10260
rect 7607 10220 8208 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12124 10220 12817 10248
rect 12124 10208 12130 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 11517 10183 11575 10189
rect 11517 10149 11529 10183
rect 11563 10180 11575 10183
rect 13814 10180 13820 10192
rect 11563 10152 13820 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 6178 10112 6184 10124
rect 6139 10084 6184 10112
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 13446 10112 13452 10124
rect 13407 10084 13452 10112
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 14366 10112 14372 10124
rect 14327 10084 14372 10112
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 14918 10112 14924 10124
rect 14660 10084 14924 10112
rect 1578 10004 1584 10056
rect 1636 10044 1642 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 1636 10016 2973 10044
rect 1636 10004 1642 10016
rect 2961 10013 2973 10016
rect 3007 10044 3019 10047
rect 3418 10044 3424 10056
rect 3007 10016 3424 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3418 10004 3424 10016
rect 3476 10044 3482 10056
rect 4062 10044 4068 10056
rect 3476 10016 4068 10044
rect 3476 10004 3482 10016
rect 4062 10004 4068 10016
rect 4120 10044 4126 10056
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 4120 10016 4353 10044
rect 4120 10004 4126 10016
rect 4341 10013 4353 10016
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 4608 10047 4666 10053
rect 4608 10013 4620 10047
rect 4654 10044 4666 10047
rect 5718 10044 5724 10056
rect 4654 10016 5724 10044
rect 4654 10013 4666 10016
rect 4608 10007 4666 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 6196 10044 6224 10072
rect 7190 10044 7196 10056
rect 6196 10016 7196 10044
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9732 10016 10149 10044
rect 9732 10004 9738 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10404 10047 10462 10053
rect 10404 10013 10416 10047
rect 10450 10044 10462 10047
rect 12526 10044 12532 10056
rect 10450 10016 12532 10044
rect 10450 10013 10462 10016
rect 10404 10007 10462 10013
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14660 10053 14688 10084
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 14645 10047 14703 10053
rect 14240 10016 14596 10044
rect 14240 10004 14246 10016
rect 2716 9979 2774 9985
rect 2716 9945 2728 9979
rect 2762 9976 2774 9979
rect 4430 9976 4436 9988
rect 2762 9948 4436 9976
rect 2762 9945 2774 9948
rect 2716 9939 2774 9945
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 5994 9936 6000 9988
rect 6052 9976 6058 9988
rect 6426 9979 6484 9985
rect 6426 9976 6438 9979
rect 6052 9948 6438 9976
rect 6052 9936 6058 9948
rect 6426 9945 6438 9948
rect 6472 9945 6484 9979
rect 6426 9939 6484 9945
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 13173 9979 13231 9985
rect 13173 9976 13185 9979
rect 11204 9948 13185 9976
rect 11204 9936 11210 9948
rect 13173 9945 13185 9948
rect 13219 9945 13231 9979
rect 14274 9976 14280 9988
rect 14235 9948 14280 9976
rect 13173 9939 13231 9945
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14568 9976 14596 10016
rect 14645 10013 14657 10047
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 16206 10044 16212 10056
rect 16167 10016 16212 10044
rect 14737 10007 14795 10013
rect 14752 9976 14780 10007
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 16574 10044 16580 10056
rect 16535 10016 16580 10044
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 14568 9948 14780 9976
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 13311 9880 14933 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 15654 9908 15660 9920
rect 15615 9880 15660 9908
rect 14921 9871 14979 9877
rect 15654 9868 15660 9880
rect 15712 9868 15718 9920
rect 1104 9818 22976 9840
rect 1104 9766 6378 9818
rect 6430 9766 6442 9818
rect 6494 9766 6506 9818
rect 6558 9766 6570 9818
rect 6622 9766 6634 9818
rect 6686 9766 11806 9818
rect 11858 9766 11870 9818
rect 11922 9766 11934 9818
rect 11986 9766 11998 9818
rect 12050 9766 12062 9818
rect 12114 9766 17234 9818
rect 17286 9766 17298 9818
rect 17350 9766 17362 9818
rect 17414 9766 17426 9818
rect 17478 9766 17490 9818
rect 17542 9766 22662 9818
rect 22714 9766 22726 9818
rect 22778 9766 22790 9818
rect 22842 9766 22854 9818
rect 22906 9766 22918 9818
rect 22970 9766 22976 9818
rect 1104 9744 22976 9766
rect 1848 9639 1906 9645
rect 1848 9605 1860 9639
rect 1894 9636 1906 9639
rect 1946 9636 1952 9648
rect 1894 9608 1952 9636
rect 1894 9605 1906 9608
rect 1848 9599 1906 9605
rect 1946 9596 1952 9608
rect 2004 9596 2010 9648
rect 4240 9639 4298 9645
rect 4240 9605 4252 9639
rect 4286 9636 4298 9639
rect 4338 9636 4344 9648
rect 4286 9608 4344 9636
rect 4286 9605 4298 9608
rect 4240 9599 4298 9605
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 9398 9636 9404 9648
rect 9456 9645 9462 9648
rect 9368 9608 9404 9636
rect 9398 9596 9404 9608
rect 9456 9599 9468 9645
rect 13354 9636 13360 9648
rect 13315 9608 13360 9636
rect 9456 9596 9462 9599
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 15565 9639 15623 9645
rect 15565 9605 15577 9639
rect 15611 9636 15623 9639
rect 16574 9636 16580 9648
rect 15611 9608 16580 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9568 4031 9571
rect 4062 9568 4068 9580
rect 4019 9540 4068 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13495 9540 14197 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14918 9568 14924 9580
rect 14415 9540 14924 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 16206 9568 16212 9580
rect 15344 9540 16212 9568
rect 15344 9528 15350 9540
rect 16206 9528 16212 9540
rect 16264 9568 16270 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16264 9540 16865 9568
rect 16264 9528 16270 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 9674 9500 9680 9512
rect 9635 9472 9680 9500
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 13538 9500 13544 9512
rect 13499 9472 13544 9500
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 13872 9472 14657 9500
rect 13872 9460 13878 9472
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 14645 9463 14703 9469
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 2961 9435 3019 9441
rect 2961 9432 2973 9435
rect 2924 9404 2973 9432
rect 2924 9392 2930 9404
rect 2961 9401 2973 9404
rect 3007 9401 3019 9435
rect 2961 9395 3019 9401
rect 5353 9435 5411 9441
rect 5353 9401 5365 9435
rect 5399 9432 5411 9435
rect 5902 9432 5908 9444
rect 5399 9404 5908 9432
rect 5399 9401 5411 9404
rect 5353 9395 5411 9401
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 14553 9435 14611 9441
rect 14553 9401 14565 9435
rect 14599 9432 14611 9435
rect 15010 9432 15016 9444
rect 14599 9404 15016 9432
rect 14599 9401 14611 9404
rect 14553 9395 14611 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 16942 9392 16948 9444
rect 17000 9432 17006 9444
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 17000 9404 17141 9432
rect 17000 9392 17006 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 17129 9395 17187 9401
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 9766 9364 9772 9376
rect 8343 9336 9772 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12952 9336 13001 9364
rect 12952 9324 12958 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17313 9367 17371 9373
rect 17313 9364 17325 9367
rect 17092 9336 17325 9364
rect 17092 9324 17098 9336
rect 17313 9333 17325 9336
rect 17359 9333 17371 9367
rect 17313 9327 17371 9333
rect 1104 9274 22816 9296
rect 1104 9222 3664 9274
rect 3716 9222 3728 9274
rect 3780 9222 3792 9274
rect 3844 9222 3856 9274
rect 3908 9222 3920 9274
rect 3972 9222 9092 9274
rect 9144 9222 9156 9274
rect 9208 9222 9220 9274
rect 9272 9222 9284 9274
rect 9336 9222 9348 9274
rect 9400 9222 14520 9274
rect 14572 9222 14584 9274
rect 14636 9222 14648 9274
rect 14700 9222 14712 9274
rect 14764 9222 14776 9274
rect 14828 9222 19948 9274
rect 20000 9222 20012 9274
rect 20064 9222 20076 9274
rect 20128 9222 20140 9274
rect 20192 9222 20204 9274
rect 20256 9222 22816 9274
rect 1104 9200 22816 9222
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 4672 9132 5365 9160
rect 4672 9120 4678 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5353 9123 5411 9129
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 8938 9160 8944 9172
rect 8619 9132 8944 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 14274 9160 14280 9172
rect 13403 9132 14280 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14366 9120 14372 9172
rect 14424 9160 14430 9172
rect 17678 9160 17684 9172
rect 14424 9132 17684 9160
rect 14424 9120 14430 9132
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 11517 9095 11575 9101
rect 11517 9061 11529 9095
rect 11563 9092 11575 9095
rect 16025 9095 16083 9101
rect 11563 9064 12434 9092
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 9732 8996 10149 9024
rect 9732 8984 9738 8996
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 12406 9024 12434 9064
rect 16025 9061 16037 9095
rect 16071 9092 16083 9095
rect 16669 9095 16727 9101
rect 16669 9092 16681 9095
rect 16071 9064 16681 9092
rect 16071 9061 16083 9064
rect 16025 9055 16083 9061
rect 16669 9061 16681 9064
rect 16715 9061 16727 9095
rect 16669 9055 16727 9061
rect 18325 9095 18383 9101
rect 18325 9061 18337 9095
rect 18371 9092 18383 9095
rect 18598 9092 18604 9104
rect 18371 9064 18604 9092
rect 18371 9061 18383 9064
rect 18325 9055 18383 9061
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 19610 9092 19616 9104
rect 19306 9064 19616 9092
rect 13354 9024 13360 9036
rect 12406 8996 13360 9024
rect 10137 8987 10195 8993
rect 13354 8984 13360 8996
rect 13412 9024 13418 9036
rect 13412 8996 13676 9024
rect 13412 8984 13418 8996
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 4062 8956 4068 8968
rect 4019 8928 4068 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4246 8965 4252 8968
rect 4240 8919 4252 8965
rect 4304 8956 4310 8968
rect 7460 8959 7518 8965
rect 4304 8928 4340 8956
rect 4246 8916 4252 8919
rect 4304 8916 4310 8928
rect 7460 8925 7472 8959
rect 7506 8956 7518 8959
rect 8386 8956 8392 8968
rect 7506 8928 8392 8956
rect 7506 8925 7518 8928
rect 7460 8919 7518 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 12894 8956 12900 8968
rect 12855 8928 12900 8956
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 13648 8965 13676 8996
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 15887 9027 15945 9033
rect 15887 9024 15899 9027
rect 15712 8996 15899 9024
rect 15712 8984 15718 8996
rect 15887 8993 15899 8996
rect 15933 8993 15945 9027
rect 19306 9024 19334 9064
rect 19610 9052 19616 9064
rect 19668 9052 19674 9104
rect 15887 8987 15945 8993
rect 16776 8996 19334 9024
rect 16776 8968 16804 8996
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 10404 8891 10462 8897
rect 10404 8857 10416 8891
rect 10450 8888 10462 8891
rect 10450 8860 12434 8888
rect 10450 8857 10462 8860
rect 10404 8851 10462 8857
rect 12406 8820 12434 8860
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 13320 8860 13369 8888
rect 13320 8848 13326 8860
rect 13357 8857 13369 8860
rect 13403 8857 13415 8891
rect 13357 8851 13415 8857
rect 13541 8891 13599 8897
rect 13541 8857 13553 8891
rect 13587 8888 13599 8891
rect 13814 8888 13820 8900
rect 13587 8860 13820 8888
rect 13587 8857 13599 8860
rect 13541 8851 13599 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 15764 8888 15792 8919
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 16209 8959 16267 8965
rect 16209 8956 16221 8959
rect 16172 8928 16221 8956
rect 16172 8916 16178 8928
rect 16209 8925 16221 8928
rect 16255 8925 16267 8959
rect 16209 8919 16267 8925
rect 16669 8959 16727 8965
rect 16669 8925 16681 8959
rect 16715 8956 16727 8959
rect 16758 8956 16764 8968
rect 16715 8928 16764 8956
rect 16715 8925 16727 8928
rect 16669 8919 16727 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 16899 8928 17417 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17770 8956 17776 8968
rect 17635 8928 17776 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 16390 8888 16396 8900
rect 15764 8860 16396 8888
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 16868 8888 16896 8919
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 18046 8956 18052 8968
rect 18007 8928 18052 8956
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 19702 8916 19708 8968
rect 19760 8956 19766 8968
rect 19797 8959 19855 8965
rect 19797 8956 19809 8959
rect 19760 8928 19809 8956
rect 19760 8916 19766 8928
rect 19797 8925 19809 8928
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 16540 8860 16896 8888
rect 16540 8848 16546 8860
rect 16942 8848 16948 8900
rect 17000 8888 17006 8900
rect 18141 8891 18199 8897
rect 18141 8888 18153 8891
rect 17000 8860 18153 8888
rect 17000 8848 17006 8860
rect 18141 8857 18153 8860
rect 18187 8857 18199 8891
rect 18141 8851 18199 8857
rect 18325 8891 18383 8897
rect 18325 8857 18337 8891
rect 18371 8888 18383 8891
rect 18966 8888 18972 8900
rect 18371 8860 18972 8888
rect 18371 8857 18383 8860
rect 18325 8851 18383 8857
rect 18966 8848 18972 8860
rect 19024 8848 19030 8900
rect 12713 8823 12771 8829
rect 12713 8820 12725 8823
rect 12406 8792 12725 8820
rect 12713 8789 12725 8792
rect 12759 8789 12771 8823
rect 16206 8820 16212 8832
rect 16167 8792 16212 8820
rect 12713 8783 12771 8789
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 16356 8792 17417 8820
rect 16356 8780 16362 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 17405 8783 17463 8789
rect 1104 8730 22976 8752
rect 1104 8678 6378 8730
rect 6430 8678 6442 8730
rect 6494 8678 6506 8730
rect 6558 8678 6570 8730
rect 6622 8678 6634 8730
rect 6686 8678 11806 8730
rect 11858 8678 11870 8730
rect 11922 8678 11934 8730
rect 11986 8678 11998 8730
rect 12050 8678 12062 8730
rect 12114 8678 17234 8730
rect 17286 8678 17298 8730
rect 17350 8678 17362 8730
rect 17414 8678 17426 8730
rect 17478 8678 17490 8730
rect 17542 8678 22662 8730
rect 22714 8678 22726 8730
rect 22778 8678 22790 8730
rect 22842 8678 22854 8730
rect 22906 8678 22918 8730
rect 22970 8678 22976 8730
rect 1104 8656 22976 8678
rect 3605 8619 3663 8625
rect 3605 8585 3617 8619
rect 3651 8616 3663 8619
rect 4706 8616 4712 8628
rect 3651 8588 4712 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 7466 8616 7472 8628
rect 7427 8588 7472 8616
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11606 8616 11612 8628
rect 11195 8588 11612 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11606 8576 11612 8588
rect 11664 8576 11670 8628
rect 16853 8619 16911 8625
rect 16853 8616 16865 8619
rect 12406 8588 16865 8616
rect 2222 8508 2228 8560
rect 2280 8548 2286 8560
rect 2470 8551 2528 8557
rect 2470 8548 2482 8551
rect 2280 8520 2482 8548
rect 2280 8508 2286 8520
rect 2470 8517 2482 8520
rect 2516 8517 2528 8551
rect 2470 8511 2528 8517
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 10036 8551 10094 8557
rect 7248 8520 8892 8548
rect 7248 8508 7254 8520
rect 4062 8480 4068 8492
rect 4023 8452 4068 8480
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 8593 8483 8651 8489
rect 8593 8449 8605 8483
rect 8639 8480 8651 8483
rect 8754 8480 8760 8492
rect 8639 8452 8760 8480
rect 8639 8449 8651 8452
rect 8593 8443 8651 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 8864 8489 8892 8520
rect 10036 8517 10048 8551
rect 10082 8548 10094 8551
rect 12406 8548 12434 8588
rect 16853 8585 16865 8588
rect 16899 8585 16911 8619
rect 18046 8616 18052 8628
rect 18007 8588 18052 8616
rect 16853 8579 16911 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 19610 8576 19616 8628
rect 19668 8616 19674 8628
rect 19668 8588 20024 8616
rect 19668 8576 19674 8588
rect 10082 8520 12434 8548
rect 10082 8517 10094 8520
rect 10036 8511 10094 8517
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 15654 8548 15660 8560
rect 13320 8520 15660 8548
rect 13320 8508 13326 8520
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9674 8480 9680 8492
rect 8895 8452 9680 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9674 8440 9680 8452
rect 9732 8480 9738 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9732 8452 9781 8480
rect 9732 8440 9738 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 13817 8443 13875 8449
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 1636 8384 2237 8412
rect 1636 8372 1642 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4430 8344 4436 8356
rect 4203 8316 4436 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4430 8304 4436 8316
rect 4488 8304 4494 8356
rect 13832 8344 13860 8443
rect 13906 8440 13912 8492
rect 13964 8480 13970 8492
rect 14090 8480 14096 8492
rect 13964 8452 14009 8480
rect 14051 8452 14096 8480
rect 13964 8440 13970 8452
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 14366 8480 14372 8492
rect 14240 8452 14372 8480
rect 14240 8440 14246 8452
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 14844 8489 14872 8520
rect 15654 8508 15660 8520
rect 15712 8548 15718 8560
rect 15712 8520 15976 8548
rect 15712 8508 15718 8520
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15948 8489 15976 8520
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 19886 8548 19892 8560
rect 16448 8520 17908 8548
rect 16448 8508 16454 8520
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15528 8452 15761 8480
rect 15528 8440 15534 8452
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 13998 8372 14004 8424
rect 14056 8412 14062 8424
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14056 8384 14657 8412
rect 14056 8372 14062 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8412 15071 8415
rect 15654 8412 15660 8424
rect 15059 8384 15660 8412
rect 15059 8381 15071 8384
rect 15013 8375 15071 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15948 8412 15976 8443
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 16264 8452 17049 8480
rect 16264 8440 16270 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17678 8480 17684 8492
rect 17267 8452 17684 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 17880 8489 17908 8520
rect 18800 8520 19892 8548
rect 18800 8489 18828 8520
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 19996 8557 20024 8588
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20128 8588 20944 8616
rect 20128 8576 20134 8588
rect 20916 8557 20944 8588
rect 19981 8551 20039 8557
rect 19981 8517 19993 8551
rect 20027 8517 20039 8551
rect 19981 8511 20039 8517
rect 20901 8551 20959 8557
rect 20901 8517 20913 8551
rect 20947 8517 20959 8551
rect 20901 8511 20959 8517
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18785 8483 18843 8489
rect 18095 8452 18736 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 16666 8412 16672 8424
rect 15948 8384 16672 8412
rect 16666 8372 16672 8384
rect 16724 8412 16730 8424
rect 16942 8412 16948 8424
rect 16724 8384 16948 8412
rect 16724 8372 16730 8384
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 17359 8384 18613 8412
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18708 8412 18736 8452
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18966 8480 18972 8492
rect 18927 8452 18972 8480
rect 18785 8443 18843 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19150 8480 19156 8492
rect 19107 8452 19156 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19260 8412 19288 8443
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19576 8452 19717 8480
rect 19576 8440 19582 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 19852 8452 19897 8480
rect 19852 8440 19858 8452
rect 20070 8440 20076 8492
rect 20128 8480 20134 8492
rect 20211 8483 20269 8489
rect 20128 8452 20173 8480
rect 20128 8440 20134 8452
rect 20211 8449 20223 8483
rect 20257 8480 20269 8483
rect 20346 8480 20352 8492
rect 20257 8452 20352 8480
rect 20257 8449 20269 8452
rect 20211 8443 20269 8449
rect 20346 8440 20352 8452
rect 20404 8480 20410 8492
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20404 8452 20821 8480
rect 20404 8440 20410 8452
rect 20809 8449 20821 8452
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 20993 8483 21051 8489
rect 20993 8449 21005 8483
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 18708 8384 19012 8412
rect 19260 8384 20392 8412
rect 18601 8375 18659 8381
rect 15194 8344 15200 8356
rect 13832 8316 15200 8344
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 15841 8347 15899 8353
rect 15841 8313 15853 8347
rect 15887 8344 15899 8347
rect 18414 8344 18420 8356
rect 15887 8316 18420 8344
rect 15887 8313 15899 8316
rect 15841 8307 15899 8313
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 18874 8344 18880 8356
rect 18835 8316 18880 8344
rect 18874 8304 18880 8316
rect 18932 8304 18938 8356
rect 18984 8344 19012 8384
rect 19610 8344 19616 8356
rect 18984 8316 19616 8344
rect 19610 8304 19616 8316
rect 19668 8344 19674 8356
rect 20070 8344 20076 8356
rect 19668 8316 20076 8344
rect 19668 8304 19674 8316
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 20364 8353 20392 8384
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 21008 8412 21036 8443
rect 20496 8384 21036 8412
rect 20496 8372 20502 8384
rect 20349 8347 20407 8353
rect 20349 8313 20361 8347
rect 20395 8313 20407 8347
rect 20349 8307 20407 8313
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5442 8276 5448 8288
rect 5123 8248 5448 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 13412 8248 13645 8276
rect 13412 8236 13418 8248
rect 13633 8245 13645 8248
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 19058 8276 19064 8288
rect 17736 8248 19064 8276
rect 17736 8236 17742 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 1104 8186 22816 8208
rect 1104 8134 3664 8186
rect 3716 8134 3728 8186
rect 3780 8134 3792 8186
rect 3844 8134 3856 8186
rect 3908 8134 3920 8186
rect 3972 8134 9092 8186
rect 9144 8134 9156 8186
rect 9208 8134 9220 8186
rect 9272 8134 9284 8186
rect 9336 8134 9348 8186
rect 9400 8134 14520 8186
rect 14572 8134 14584 8186
rect 14636 8134 14648 8186
rect 14700 8134 14712 8186
rect 14764 8134 14776 8186
rect 14828 8134 19948 8186
rect 20000 8134 20012 8186
rect 20064 8134 20076 8186
rect 20128 8134 20140 8186
rect 20192 8134 20204 8186
rect 20256 8134 22816 8186
rect 1104 8112 22816 8134
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 6328 8044 6561 8072
rect 6328 8032 6334 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8536 8044 8585 8072
rect 8536 8032 8542 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 12710 8072 12716 8084
rect 11563 8044 12716 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 15194 8072 15200 8084
rect 15155 8044 15200 8072
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 16540 8044 17785 8072
rect 16540 8032 16546 8044
rect 17773 8041 17785 8044
rect 17819 8072 17831 8075
rect 18601 8075 18659 8081
rect 18601 8072 18613 8075
rect 17819 8044 18613 8072
rect 17819 8041 17831 8044
rect 17773 8035 17831 8041
rect 18601 8041 18613 8044
rect 18647 8041 18659 8075
rect 18601 8035 18659 8041
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 18966 8072 18972 8084
rect 18831 8044 18972 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19794 8072 19800 8084
rect 19659 8044 19800 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 19794 8032 19800 8044
rect 19852 8032 19858 8084
rect 14461 8007 14519 8013
rect 14461 7973 14473 8007
rect 14507 8004 14519 8007
rect 14507 7976 17448 8004
rect 14507 7973 14519 7976
rect 14461 7967 14519 7973
rect 1578 7936 1584 7948
rect 1539 7908 1584 7936
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 4798 7936 4804 7948
rect 4359 7908 4804 7936
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4359 7877 4387 7908
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 7190 7936 7196 7948
rect 7151 7908 7196 7936
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10137 7939 10195 7945
rect 10137 7936 10149 7939
rect 9732 7908 10149 7936
rect 9732 7896 9738 7908
rect 10137 7905 10149 7908
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13044 7908 14289 7936
rect 13044 7896 13050 7908
rect 4065 7871 4123 7877
rect 4344 7871 4402 7877
rect 4065 7868 4077 7871
rect 3384 7840 4077 7868
rect 3384 7828 3390 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4249 7865 4307 7871
rect 4249 7831 4261 7865
rect 4295 7831 4307 7865
rect 4344 7837 4356 7871
rect 4390 7837 4402 7871
rect 4344 7831 4402 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4249 7825 4307 7831
rect 1848 7803 1906 7809
rect 1848 7769 1860 7803
rect 1894 7800 1906 7803
rect 1946 7800 1952 7812
rect 1894 7772 1952 7800
rect 1894 7769 1906 7772
rect 1848 7763 1906 7769
rect 1946 7760 1952 7772
rect 2004 7760 2010 7812
rect 2961 7735 3019 7741
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 4062 7732 4068 7744
rect 3007 7704 4068 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4264 7732 4292 7825
rect 4448 7800 4476 7831
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4672 7840 5181 7868
rect 4672 7828 4678 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 12894 7868 12900 7880
rect 12391 7840 12900 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13262 7868 13268 7880
rect 13223 7840 13268 7868
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13372 7877 13400 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 15654 7936 15660 7948
rect 15615 7908 15660 7936
rect 14277 7899 14335 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15804 7908 15853 7936
rect 15804 7896 15810 7908
rect 15841 7905 15853 7908
rect 15887 7936 15899 7939
rect 16298 7936 16304 7948
rect 15887 7908 16304 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 17420 7936 17448 7976
rect 17494 7964 17500 8016
rect 17552 8004 17558 8016
rect 17552 7976 19472 8004
rect 17552 7964 17558 7976
rect 17678 7936 17684 7948
rect 17420 7908 17684 7936
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7837 13415 7871
rect 13630 7868 13636 7880
rect 13591 7840 13636 7868
rect 13357 7831 13415 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14553 7871 14611 7877
rect 13780 7840 13825 7868
rect 13780 7828 13786 7840
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15194 7868 15200 7880
rect 14599 7840 15200 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 15528 7840 16405 7868
rect 15528 7828 15534 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16666 7868 16672 7880
rect 16623 7840 16672 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 19334 7868 19340 7880
rect 17604 7840 19340 7868
rect 4890 7800 4896 7812
rect 4448 7772 4896 7800
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 5442 7809 5448 7812
rect 5436 7800 5448 7809
rect 5403 7772 5448 7800
rect 5436 7763 5448 7772
rect 5442 7760 5448 7763
rect 5500 7760 5506 7812
rect 7460 7803 7518 7809
rect 7460 7769 7472 7803
rect 7506 7800 7518 7803
rect 10226 7800 10232 7812
rect 7506 7772 10232 7800
rect 7506 7769 7518 7772
rect 7460 7763 7518 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 10404 7803 10462 7809
rect 10404 7769 10416 7803
rect 10450 7800 10462 7803
rect 13280 7800 13308 7828
rect 10450 7772 13308 7800
rect 13449 7803 13507 7809
rect 10450 7769 10462 7772
rect 10404 7763 10462 7769
rect 13449 7769 13461 7803
rect 13495 7800 13507 7803
rect 13998 7800 14004 7812
rect 13495 7772 14004 7800
rect 13495 7769 13507 7772
rect 13449 7763 13507 7769
rect 13998 7760 14004 7772
rect 14056 7760 14062 7812
rect 15654 7760 15660 7812
rect 15712 7800 15718 7812
rect 17604 7809 17632 7840
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 19444 7877 19472 7976
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7936 19763 7939
rect 19794 7936 19800 7948
rect 19751 7908 19800 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 19794 7896 19800 7908
rect 19852 7896 19858 7948
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7868 19579 7871
rect 20162 7868 20168 7880
rect 19567 7840 20168 7868
rect 19567 7837 19579 7840
rect 19521 7831 19579 7837
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20530 7868 20536 7880
rect 20395 7840 20536 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 15712 7772 17601 7800
rect 15712 7760 15718 7772
rect 17589 7769 17601 7772
rect 17635 7769 17647 7803
rect 17589 7763 17647 7769
rect 17770 7760 17776 7812
rect 17828 7809 17834 7812
rect 17828 7803 17847 7809
rect 17835 7800 17847 7803
rect 17835 7772 18368 7800
rect 17835 7769 17847 7772
rect 17828 7763 17847 7769
rect 17828 7760 17834 7763
rect 4522 7732 4528 7744
rect 4264 7704 4528 7732
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7732 12495 7735
rect 12618 7732 12624 7744
rect 12483 7704 12624 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12989 7735 13047 7741
rect 12989 7701 13001 7735
rect 13035 7732 13047 7735
rect 13262 7732 13268 7744
rect 13035 7704 13268 7732
rect 13035 7701 13047 7704
rect 12989 7695 13047 7701
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 13596 7704 14565 7732
rect 13596 7692 13602 7704
rect 14553 7701 14565 7704
rect 14599 7701 14611 7735
rect 14553 7695 14611 7701
rect 15010 7692 15016 7744
rect 15068 7732 15074 7744
rect 15470 7732 15476 7744
rect 15068 7704 15476 7732
rect 15068 7692 15074 7704
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 15930 7732 15936 7744
rect 15611 7704 15936 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 15930 7692 15936 7704
rect 15988 7732 15994 7744
rect 16761 7735 16819 7741
rect 16761 7732 16773 7735
rect 15988 7704 16773 7732
rect 15988 7692 15994 7704
rect 16761 7701 16773 7704
rect 16807 7732 16819 7735
rect 17494 7732 17500 7744
rect 16807 7704 17500 7732
rect 16807 7701 16819 7704
rect 16761 7695 16819 7701
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18340 7732 18368 7772
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 18472 7772 18517 7800
rect 18472 7760 18478 7772
rect 18617 7735 18675 7741
rect 18617 7732 18629 7735
rect 18340 7704 18629 7732
rect 18617 7701 18629 7704
rect 18663 7732 18675 7735
rect 19702 7732 19708 7744
rect 18663 7704 19708 7732
rect 18663 7701 18675 7704
rect 18617 7695 18675 7701
rect 19702 7692 19708 7704
rect 19760 7732 19766 7744
rect 20257 7735 20315 7741
rect 20257 7732 20269 7735
rect 19760 7704 20269 7732
rect 19760 7692 19766 7704
rect 20257 7701 20269 7704
rect 20303 7701 20315 7735
rect 20257 7695 20315 7701
rect 1104 7642 22976 7664
rect 1104 7590 6378 7642
rect 6430 7590 6442 7642
rect 6494 7590 6506 7642
rect 6558 7590 6570 7642
rect 6622 7590 6634 7642
rect 6686 7590 11806 7642
rect 11858 7590 11870 7642
rect 11922 7590 11934 7642
rect 11986 7590 11998 7642
rect 12050 7590 12062 7642
rect 12114 7590 17234 7642
rect 17286 7590 17298 7642
rect 17350 7590 17362 7642
rect 17414 7590 17426 7642
rect 17478 7590 17490 7642
rect 17542 7590 22662 7642
rect 22714 7590 22726 7642
rect 22778 7590 22790 7642
rect 22842 7590 22854 7642
rect 22906 7590 22918 7642
rect 22970 7590 22976 7642
rect 1104 7568 22976 7590
rect 1946 7528 1952 7540
rect 1907 7500 1952 7528
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5261 7531 5319 7537
rect 5261 7528 5273 7531
rect 4120 7500 5273 7528
rect 4120 7488 4126 7500
rect 5261 7497 5273 7500
rect 5307 7497 5319 7531
rect 13998 7528 14004 7540
rect 13959 7500 14004 7528
rect 5261 7491 5319 7497
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 17126 7528 17132 7540
rect 16347 7500 17132 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 17126 7488 17132 7500
rect 17184 7488 17190 7540
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 1636 7432 2605 7460
rect 1636 7420 1642 7432
rect 2593 7429 2605 7432
rect 2639 7429 2651 7463
rect 2593 7423 2651 7429
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 7374 7460 7380 7472
rect 4387 7432 7380 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 7374 7420 7380 7432
rect 7432 7460 7438 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7432 7432 7849 7460
rect 7432 7420 7438 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 9674 7460 9680 7472
rect 9631 7432 9680 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 15289 7463 15347 7469
rect 15289 7429 15301 7463
rect 15335 7460 15347 7463
rect 16022 7460 16028 7472
rect 15335 7432 16028 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 16022 7420 16028 7432
rect 16080 7420 16086 7472
rect 17954 7420 17960 7472
rect 18012 7460 18018 7472
rect 18506 7460 18512 7472
rect 18012 7432 18512 7460
rect 18012 7420 18018 7432
rect 18506 7420 18512 7432
rect 18564 7460 18570 7472
rect 18564 7432 18920 7460
rect 18564 7420 18570 7432
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 5166 7392 5172 7404
rect 2179 7364 2774 7392
rect 5127 7364 5172 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2746 7256 2774 7364
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5316 7364 6561 7392
rect 5316 7352 5322 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12676 7364 13093 7392
rect 12676 7352 12682 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13262 7392 13268 7404
rect 13223 7364 13268 7392
rect 13081 7355 13139 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13354 7352 13360 7404
rect 13412 7392 13418 7404
rect 14093 7395 14151 7401
rect 13412 7364 13457 7392
rect 13412 7352 13418 7364
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 15010 7392 15016 7404
rect 14139 7364 15016 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 5445 7327 5503 7333
rect 5445 7324 5457 7327
rect 5408 7296 5457 7324
rect 5408 7284 5414 7296
rect 5445 7293 5457 7296
rect 5491 7324 5503 7327
rect 13173 7327 13231 7333
rect 5491 7296 6960 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 2746 7228 4813 7256
rect 4801 7225 4813 7228
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 6932 7200 6960 7296
rect 13173 7293 13185 7327
rect 13219 7324 13231 7327
rect 13538 7324 13544 7336
rect 13219 7296 13544 7324
rect 13219 7293 13231 7296
rect 13173 7287 13231 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 14108 7256 14136 7355
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 15194 7392 15200 7404
rect 15155 7364 15200 7392
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15304 7364 15485 7392
rect 12400 7228 14136 7256
rect 12400 7216 12406 7228
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 4948 7160 6653 7188
rect 4948 7148 4954 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 6972 7160 7205 7188
rect 6972 7148 6978 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 11296 7160 12909 7188
rect 11296 7148 11302 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 13630 7148 13636 7200
rect 13688 7188 13694 7200
rect 15304 7188 15332 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7361 15991 7395
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 15933 7355 15991 7361
rect 15948 7324 15976 7355
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 18417 7395 18475 7401
rect 18417 7392 18429 7395
rect 17727 7364 18429 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 18417 7361 18429 7364
rect 18463 7361 18475 7395
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18417 7355 18475 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 18690 7352 18696 7404
rect 18748 7392 18754 7404
rect 18892 7401 18920 7432
rect 19334 7420 19340 7472
rect 19392 7460 19398 7472
rect 19889 7463 19947 7469
rect 19889 7460 19901 7463
rect 19392 7432 19901 7460
rect 19392 7420 19398 7432
rect 19889 7429 19901 7432
rect 19935 7460 19947 7463
rect 20346 7460 20352 7472
rect 19935 7432 20352 7460
rect 19935 7429 19947 7432
rect 19889 7423 19947 7429
rect 20346 7420 20352 7432
rect 20404 7420 20410 7472
rect 18877 7395 18935 7401
rect 18748 7364 18793 7392
rect 18748 7352 18754 7364
rect 18877 7361 18889 7395
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7392 19027 7395
rect 19058 7392 19064 7404
rect 19015 7364 19064 7392
rect 19015 7361 19027 7364
rect 18969 7355 19027 7361
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 15488 7296 15976 7324
rect 15488 7265 15516 7296
rect 16022 7284 16028 7336
rect 16080 7324 16086 7336
rect 17586 7324 17592 7336
rect 16080 7296 16896 7324
rect 17547 7296 17592 7324
rect 16080 7284 16086 7296
rect 15473 7259 15531 7265
rect 15473 7225 15485 7259
rect 15519 7225 15531 7259
rect 16758 7256 16764 7268
rect 15473 7219 15531 7225
rect 15856 7228 16764 7256
rect 15856 7188 15884 7228
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 16868 7256 16896 7296
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 17770 7324 17776 7336
rect 17731 7296 17776 7324
rect 17770 7284 17776 7296
rect 17828 7284 17834 7336
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7324 17923 7327
rect 18230 7324 18236 7336
rect 17911 7296 18236 7324
rect 17911 7293 17923 7296
rect 17865 7287 17923 7293
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 18690 7256 18696 7268
rect 16868 7228 18696 7256
rect 18690 7216 18696 7228
rect 18748 7216 18754 7268
rect 20162 7256 20168 7268
rect 20123 7228 20168 7256
rect 20162 7216 20168 7228
rect 20220 7216 20226 7268
rect 16022 7188 16028 7200
rect 13688 7160 15884 7188
rect 15983 7160 16028 7188
rect 13688 7148 13694 7160
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 16776 7188 16804 7216
rect 16942 7188 16948 7200
rect 16776 7160 16948 7188
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 20180 7188 20208 7216
rect 20346 7188 20352 7200
rect 17920 7160 20208 7188
rect 20307 7160 20352 7188
rect 17920 7148 17926 7160
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 1104 7098 22816 7120
rect 1104 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 9092 7098
rect 9144 7046 9156 7098
rect 9208 7046 9220 7098
rect 9272 7046 9284 7098
rect 9336 7046 9348 7098
rect 9400 7046 14520 7098
rect 14572 7046 14584 7098
rect 14636 7046 14648 7098
rect 14700 7046 14712 7098
rect 14764 7046 14776 7098
rect 14828 7046 19948 7098
rect 20000 7046 20012 7098
rect 20064 7046 20076 7098
rect 20128 7046 20140 7098
rect 20192 7046 20204 7098
rect 20256 7046 22816 7098
rect 1104 7024 22816 7046
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 15252 6956 16405 6984
rect 15252 6944 15258 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 15746 6916 15752 6928
rect 15707 6888 15752 6916
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 17770 6916 17776 6928
rect 16172 6888 17776 6916
rect 16172 6876 16178 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 19150 6876 19156 6928
rect 19208 6916 19214 6928
rect 19208 6888 19932 6916
rect 19208 6876 19214 6888
rect 5258 6848 5264 6860
rect 3344 6820 5264 6848
rect 3344 6792 3372 6820
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9732 6820 9781 6848
rect 9732 6808 9738 6820
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 9769 6811 9827 6817
rect 13832 6820 15577 6848
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6749 3203 6783
rect 3326 6780 3332 6792
rect 3239 6752 3332 6780
rect 3145 6743 3203 6749
rect 3160 6712 3188 6743
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 4246 6780 4252 6792
rect 3467 6752 4252 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4430 6780 4436 6792
rect 4391 6752 4436 6780
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4580 6752 4629 6780
rect 4580 6740 4586 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 4890 6780 4896 6792
rect 4847 6752 4896 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 4154 6712 4160 6724
rect 3160 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 4724 6712 4752 6743
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 10036 6783 10094 6789
rect 5092 6752 9996 6780
rect 5092 6721 5120 6752
rect 5077 6715 5135 6721
rect 4724 6684 4844 6712
rect 4816 6656 4844 6684
rect 5077 6681 5089 6715
rect 5123 6681 5135 6715
rect 5902 6712 5908 6724
rect 5863 6684 5908 6712
rect 5077 6675 5135 6681
rect 5902 6672 5908 6684
rect 5960 6712 5966 6724
rect 8113 6715 8171 6721
rect 8113 6712 8125 6715
rect 5960 6684 8125 6712
rect 5960 6672 5966 6684
rect 8113 6681 8125 6684
rect 8159 6681 8171 6715
rect 9968 6712 9996 6752
rect 10036 6749 10048 6783
rect 10082 6780 10094 6783
rect 11238 6780 11244 6792
rect 10082 6752 11244 6780
rect 10082 6749 10094 6752
rect 10036 6743 10094 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 13262 6780 13268 6792
rect 13223 6752 13268 6780
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 10502 6712 10508 6724
rect 9968 6684 10508 6712
rect 8113 6675 8171 6681
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 12989 6715 13047 6721
rect 12989 6712 13001 6715
rect 12676 6684 13001 6712
rect 12676 6672 12682 6684
rect 12989 6681 13001 6684
rect 13035 6681 13047 6715
rect 12989 6675 13047 6681
rect 13173 6715 13231 6721
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 13538 6712 13544 6724
rect 13219 6684 13544 6712
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 13538 6672 13544 6684
rect 13596 6712 13602 6724
rect 13832 6712 13860 6820
rect 15565 6817 15577 6820
rect 15611 6848 15623 6851
rect 18414 6848 18420 6860
rect 15611 6820 15700 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 13964 6752 14473 6780
rect 13964 6740 13970 6752
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 15672 6724 15700 6820
rect 15856 6820 18420 6848
rect 15856 6789 15884 6820
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 19613 6851 19671 6857
rect 19613 6848 19625 6851
rect 18748 6820 19625 6848
rect 18748 6808 18754 6820
rect 19613 6817 19625 6820
rect 19659 6817 19671 6851
rect 19794 6848 19800 6860
rect 19755 6820 19800 6848
rect 19613 6811 19671 6817
rect 19794 6808 19800 6820
rect 19852 6808 19858 6860
rect 19904 6857 19932 6888
rect 19889 6851 19947 6857
rect 19889 6817 19901 6851
rect 19935 6817 19947 6851
rect 19889 6811 19947 6817
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16301 6783 16359 6789
rect 16301 6780 16313 6783
rect 15988 6752 16313 6780
rect 15988 6740 15994 6752
rect 16301 6749 16313 6752
rect 16347 6749 16359 6783
rect 16482 6780 16488 6792
rect 16443 6752 16488 6780
rect 16301 6743 16359 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 17770 6740 17776 6792
rect 17828 6780 17834 6792
rect 18874 6780 18880 6792
rect 17828 6752 18880 6780
rect 17828 6740 17834 6752
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19702 6740 19708 6792
rect 19760 6780 19766 6792
rect 19760 6752 19805 6780
rect 19760 6740 19766 6752
rect 13596 6684 13860 6712
rect 13596 6672 13602 6684
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 15565 6715 15623 6721
rect 15565 6712 15577 6715
rect 14056 6684 15577 6712
rect 14056 6672 14062 6684
rect 15565 6681 15577 6684
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 15654 6672 15660 6724
rect 15712 6712 15718 6724
rect 16114 6712 16120 6724
rect 15712 6684 16120 6712
rect 15712 6672 15718 6684
rect 16114 6672 16120 6684
rect 16172 6672 16178 6724
rect 16942 6672 16948 6724
rect 17000 6712 17006 6724
rect 20806 6712 20812 6724
rect 17000 6684 20812 6712
rect 17000 6672 17006 6684
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 2924 6616 2973 6644
rect 2924 6604 2930 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 4798 6604 4804 6656
rect 4856 6604 4862 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 11146 6644 11152 6656
rect 11107 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 13078 6644 13084 6656
rect 13136 6653 13142 6656
rect 13045 6616 13084 6644
rect 13078 6604 13084 6616
rect 13136 6607 13145 6653
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 15010 6644 15016 6656
rect 14415 6616 15016 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 13136 6604 13142 6607
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 19392 6616 19441 6644
rect 19392 6604 19398 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 1104 6554 22976 6576
rect 1104 6502 6378 6554
rect 6430 6502 6442 6554
rect 6494 6502 6506 6554
rect 6558 6502 6570 6554
rect 6622 6502 6634 6554
rect 6686 6502 11806 6554
rect 11858 6502 11870 6554
rect 11922 6502 11934 6554
rect 11986 6502 11998 6554
rect 12050 6502 12062 6554
rect 12114 6502 17234 6554
rect 17286 6502 17298 6554
rect 17350 6502 17362 6554
rect 17414 6502 17426 6554
rect 17478 6502 17490 6554
rect 17542 6502 22662 6554
rect 22714 6502 22726 6554
rect 22778 6502 22790 6554
rect 22842 6502 22854 6554
rect 22906 6502 22918 6554
rect 22970 6502 22976 6554
rect 1104 6480 22976 6502
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3326 6440 3332 6452
rect 3007 6412 3332 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 3436 6412 5028 6440
rect 1848 6307 1906 6313
rect 1848 6273 1860 6307
rect 1894 6304 1906 6307
rect 2682 6304 2688 6316
rect 1894 6276 2688 6304
rect 1894 6273 1906 6276
rect 1848 6267 1906 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3436 6313 3464 6412
rect 4706 6332 4712 6384
rect 4764 6372 4770 6384
rect 4862 6375 4920 6381
rect 4862 6372 4874 6375
rect 4764 6344 4874 6372
rect 4764 6332 4770 6344
rect 4862 6341 4874 6344
rect 4908 6341 4920 6375
rect 5000 6372 5028 6412
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5224 6412 6009 6440
rect 5224 6400 5230 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 7837 6443 7895 6449
rect 7837 6409 7849 6443
rect 7883 6440 7895 6443
rect 8110 6440 8116 6452
rect 7883 6412 8116 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6440 11115 6443
rect 12342 6440 12348 6452
rect 11103 6412 12348 6440
rect 11103 6409 11115 6412
rect 11057 6403 11115 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6409 12771 6443
rect 16390 6440 16396 6452
rect 12713 6403 12771 6409
rect 12912 6412 16396 6440
rect 7006 6372 7012 6384
rect 5000 6344 7012 6372
rect 4862 6335 4920 6341
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 8972 6375 9030 6381
rect 8972 6341 8984 6375
rect 9018 6372 9030 6375
rect 12728 6372 12756 6403
rect 9018 6344 12756 6372
rect 9018 6341 9030 6344
rect 8972 6335 9030 6341
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6304 3663 6307
rect 4246 6304 4252 6316
rect 3651 6276 4252 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 4724 6276 6653 6304
rect 1578 6236 1584 6248
rect 1539 6208 1584 6236
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 4154 6236 4160 6248
rect 4067 6208 4160 6236
rect 4154 6196 4160 6208
rect 4212 6236 4218 6248
rect 4724 6236 4752 6276
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 6822 6304 6828 6316
rect 6687 6276 6828 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 9944 6307 10002 6313
rect 9944 6273 9956 6307
rect 9990 6304 10002 6307
rect 12912 6304 12940 6412
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17586 6440 17592 6452
rect 17543 6412 17592 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 20070 6440 20076 6452
rect 17736 6412 20076 6440
rect 17736 6400 17742 6412
rect 20070 6400 20076 6412
rect 20128 6440 20134 6452
rect 20530 6440 20536 6452
rect 20128 6412 20536 6440
rect 20128 6400 20134 6412
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 15381 6375 15439 6381
rect 15381 6372 15393 6375
rect 13311 6344 15393 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 15381 6341 15393 6344
rect 15427 6341 15439 6375
rect 15746 6372 15752 6384
rect 15381 6335 15439 6341
rect 15580 6344 15752 6372
rect 9990 6276 12940 6304
rect 12989 6307 13047 6313
rect 9990 6273 10002 6276
rect 9944 6267 10002 6273
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13817 6307 13875 6313
rect 13817 6304 13829 6307
rect 13035 6276 13829 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13817 6273 13829 6276
rect 13863 6273 13875 6307
rect 13998 6304 14004 6316
rect 13959 6276 14004 6304
rect 13817 6267 13875 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 15580 6313 15608 6344
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 17129 6375 17187 6381
rect 17129 6341 17141 6375
rect 17175 6372 17187 6375
rect 17954 6372 17960 6384
rect 17175 6344 17960 6372
rect 17175 6341 17187 6344
rect 17129 6335 17187 6341
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 18874 6372 18880 6384
rect 18835 6344 18880 6372
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 20901 6375 20959 6381
rect 20901 6372 20913 6375
rect 19628 6344 20913 6372
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 14369 6307 14427 6313
rect 14139 6276 14320 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 4212 6208 4752 6236
rect 9217 6239 9275 6245
rect 4212 6196 4218 6208
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 9490 6236 9496 6248
rect 9263 6208 9496 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 9490 6196 9496 6208
rect 9548 6236 9554 6248
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 9548 6208 9689 6236
rect 9548 6196 9554 6208
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 12894 6236 12900 6248
rect 12807 6208 12900 6236
rect 9677 6199 9735 6205
rect 12894 6196 12900 6208
rect 12952 6236 12958 6248
rect 13078 6236 13084 6248
rect 12952 6208 13084 6236
rect 12952 6196 12958 6208
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13170 6196 13176 6248
rect 13228 6236 13234 6248
rect 13357 6239 13415 6245
rect 13357 6236 13369 6239
rect 13228 6208 13369 6236
rect 13228 6196 13234 6208
rect 13357 6205 13369 6208
rect 13403 6205 13415 6239
rect 13357 6199 13415 6205
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14292 6168 14320 6276
rect 14369 6273 14381 6307
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 14384 6236 14412 6267
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15841 6307 15899 6313
rect 15712 6276 15757 6304
rect 15712 6264 15718 6276
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 15672 6236 15700 6264
rect 14384 6208 15700 6236
rect 15856 6236 15884 6267
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 16850 6304 16856 6316
rect 15988 6276 16033 6304
rect 16811 6276 16856 6304
rect 15988 6264 15994 6276
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 17221 6307 17279 6313
rect 17000 6276 17045 6304
rect 17000 6264 17006 6276
rect 17221 6273 17233 6307
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17236 6236 17264 6267
rect 17310 6264 17316 6316
rect 17368 6313 17374 6316
rect 17368 6304 17376 6313
rect 18785 6307 18843 6313
rect 17368 6276 17413 6304
rect 17368 6267 17376 6276
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 17368 6264 17374 6267
rect 18414 6236 18420 6248
rect 15856 6208 17172 6236
rect 17236 6208 18420 6236
rect 14366 6168 14372 6180
rect 14056 6140 14228 6168
rect 14292 6140 14372 6168
rect 14056 6128 14062 6140
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3568 6072 3617 6100
rect 3568 6060 3574 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 3605 6063 3663 6069
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 13446 6100 13452 6112
rect 12676 6072 13452 6100
rect 12676 6060 12682 6072
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 14200 6100 14228 6140
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 17144 6168 17172 6208
rect 18414 6196 18420 6208
rect 18472 6236 18478 6248
rect 18690 6236 18696 6248
rect 18472 6208 18696 6236
rect 18472 6196 18478 6208
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 18800 6236 18828 6267
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19153 6307 19211 6313
rect 19024 6276 19069 6304
rect 19024 6264 19030 6276
rect 19153 6273 19165 6307
rect 19199 6304 19211 6307
rect 19426 6304 19432 6316
rect 19199 6276 19432 6304
rect 19199 6273 19211 6276
rect 19153 6267 19211 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19242 6236 19248 6248
rect 18800 6208 19248 6236
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 19628 6180 19656 6344
rect 20901 6341 20913 6344
rect 20947 6341 20959 6375
rect 20901 6335 20959 6341
rect 20070 6304 20076 6316
rect 20031 6276 20076 6304
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 20806 6304 20812 6316
rect 20767 6276 20812 6304
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 20993 6307 21051 6313
rect 20993 6273 21005 6307
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 20346 6236 20352 6248
rect 20307 6208 20352 6236
rect 20346 6196 20352 6208
rect 20404 6236 20410 6248
rect 21008 6236 21036 6267
rect 20404 6208 21036 6236
rect 20404 6196 20410 6208
rect 19610 6168 19616 6180
rect 17144 6140 19616 6168
rect 19610 6128 19616 6140
rect 19668 6128 19674 6180
rect 19794 6128 19800 6180
rect 19852 6168 19858 6180
rect 20257 6171 20315 6177
rect 20257 6168 20269 6171
rect 19852 6140 20269 6168
rect 19852 6128 19858 6140
rect 20257 6137 20269 6140
rect 20303 6137 20315 6171
rect 20257 6131 20315 6137
rect 14277 6103 14335 6109
rect 14277 6100 14289 6103
rect 14200 6072 14289 6100
rect 14277 6069 14289 6072
rect 14323 6069 14335 6103
rect 14277 6063 14335 6069
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 18046 6100 18052 6112
rect 16448 6072 18052 6100
rect 16448 6060 16454 6072
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 20165 6103 20223 6109
rect 20165 6069 20177 6103
rect 20211 6100 20223 6103
rect 20530 6100 20536 6112
rect 20211 6072 20536 6100
rect 20211 6069 20223 6072
rect 20165 6063 20223 6069
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 1104 6010 22816 6032
rect 1104 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 9092 6010
rect 9144 5958 9156 6010
rect 9208 5958 9220 6010
rect 9272 5958 9284 6010
rect 9336 5958 9348 6010
rect 9400 5958 14520 6010
rect 14572 5958 14584 6010
rect 14636 5958 14648 6010
rect 14700 5958 14712 6010
rect 14764 5958 14776 6010
rect 14828 5958 19948 6010
rect 20000 5958 20012 6010
rect 20064 5958 20076 6010
rect 20128 5958 20140 6010
rect 20192 5958 20204 6010
rect 20256 5958 22816 6010
rect 1104 5936 22816 5958
rect 2682 5896 2688 5908
rect 2643 5868 2688 5896
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 4522 5856 4528 5908
rect 4580 5896 4586 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4580 5868 4813 5896
rect 4580 5856 4586 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 12713 5899 12771 5905
rect 12713 5896 12725 5899
rect 4801 5859 4859 5865
rect 9416 5868 12725 5896
rect 4338 5760 4344 5772
rect 3344 5732 4344 5760
rect 3344 5704 3372 5732
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4488 5732 4629 5760
rect 4488 5720 4494 5732
rect 4617 5729 4629 5732
rect 4663 5760 4675 5763
rect 5166 5760 5172 5772
rect 4663 5732 5172 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 3145 5655 3203 5661
rect 3160 5624 3188 5655
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 4120 5664 4169 5692
rect 4120 5652 4126 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4246 5652 4252 5704
rect 4304 5652 4310 5704
rect 4522 5692 4528 5704
rect 4483 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6052 5664 6561 5692
rect 6052 5652 6058 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6816 5695 6874 5701
rect 6816 5661 6828 5695
rect 6862 5692 6874 5695
rect 9416 5692 9444 5868
rect 12713 5865 12725 5868
rect 12759 5865 12771 5899
rect 12713 5859 12771 5865
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 13538 5896 13544 5908
rect 12860 5868 13544 5896
rect 12860 5856 12866 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14090 5856 14096 5908
rect 14148 5896 14154 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14148 5868 14289 5896
rect 14148 5856 14154 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 16758 5896 16764 5908
rect 14424 5868 16764 5896
rect 14424 5856 14430 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 16853 5899 16911 5905
rect 16853 5865 16865 5899
rect 16899 5896 16911 5899
rect 17310 5896 17316 5908
rect 16899 5868 17316 5896
rect 16899 5865 16911 5868
rect 16853 5859 16911 5865
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 19426 5896 19432 5908
rect 19387 5868 19432 5896
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 19668 5868 19809 5896
rect 19668 5856 19674 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 19797 5859 19855 5865
rect 19996 5868 21128 5896
rect 11425 5831 11483 5837
rect 11425 5797 11437 5831
rect 11471 5828 11483 5831
rect 12986 5828 12992 5840
rect 11471 5800 12992 5828
rect 11471 5797 11483 5800
rect 11425 5791 11483 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13262 5788 13268 5840
rect 13320 5828 13326 5840
rect 15841 5831 15899 5837
rect 15841 5828 15853 5831
rect 13320 5800 15853 5828
rect 13320 5788 13326 5800
rect 15841 5797 15853 5800
rect 15887 5828 15899 5831
rect 15930 5828 15936 5840
rect 15887 5800 15936 5828
rect 15887 5797 15899 5800
rect 15841 5791 15899 5797
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 17862 5828 17868 5840
rect 16132 5800 17868 5828
rect 13630 5760 13636 5772
rect 12084 5732 13636 5760
rect 6862 5664 9444 5692
rect 6862 5661 6874 5664
rect 6816 5655 6874 5661
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9548 5664 10057 5692
rect 9548 5652 9554 5664
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 12084 5701 12112 5732
rect 13630 5720 13636 5732
rect 13688 5760 13694 5772
rect 13688 5732 14320 5760
rect 13688 5720 13694 5732
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11756 5664 12081 5692
rect 11756 5652 11762 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12710 5692 12716 5704
rect 12299 5664 12716 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 12894 5695 12952 5701
rect 12894 5661 12906 5695
rect 12940 5692 12952 5695
rect 13170 5692 13176 5704
rect 12940 5664 13176 5692
rect 12940 5661 12952 5664
rect 12894 5655 12952 5661
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5692 13415 5695
rect 14182 5692 14188 5704
rect 13403 5664 14188 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 4264 5624 4292 5652
rect 5166 5624 5172 5636
rect 3160 5596 5172 5624
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 5721 5627 5779 5633
rect 5721 5624 5733 5627
rect 5592 5596 5733 5624
rect 5592 5584 5598 5596
rect 5721 5593 5733 5596
rect 5767 5593 5779 5627
rect 5721 5587 5779 5593
rect 10312 5627 10370 5633
rect 10312 5593 10324 5627
rect 10358 5624 10370 5627
rect 12161 5627 12219 5633
rect 10358 5596 11560 5624
rect 10358 5593 10370 5596
rect 10312 5587 10370 5593
rect 4246 5556 4252 5568
rect 4207 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4338 5516 4344 5568
rect 4396 5556 4402 5568
rect 5997 5559 6055 5565
rect 4396 5528 4441 5556
rect 4396 5516 4402 5528
rect 5997 5525 6009 5559
rect 6043 5556 6055 5559
rect 6822 5556 6828 5568
rect 6043 5528 6828 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7929 5559 7987 5565
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 9582 5556 9588 5568
rect 7975 5528 9588 5556
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 11532 5556 11560 5596
rect 12161 5593 12173 5627
rect 12207 5624 12219 5627
rect 12207 5596 12940 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 12802 5556 12808 5568
rect 11532 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 12912 5565 12940 5596
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13280 5624 13308 5655
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14292 5692 14320 5732
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14424 5732 14657 5760
rect 14424 5720 14430 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5760 14795 5763
rect 14918 5760 14924 5772
rect 14783 5732 14924 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 14292 5664 14473 5692
rect 14461 5661 14473 5664
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 15010 5692 15016 5704
rect 14971 5664 15016 5692
rect 14829 5655 14887 5661
rect 14090 5624 14096 5636
rect 13136 5596 14096 5624
rect 13136 5584 13142 5596
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 14844 5624 14872 5655
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 16132 5701 16160 5800
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 19996 5837 20024 5868
rect 19981 5831 20039 5837
rect 19981 5797 19993 5831
rect 20027 5797 20039 5831
rect 19981 5791 20039 5797
rect 16301 5763 16359 5769
rect 16301 5729 16313 5763
rect 16347 5760 16359 5763
rect 16666 5760 16672 5772
rect 16347 5732 16672 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 16666 5720 16672 5732
rect 16724 5760 16730 5772
rect 16724 5732 18000 5760
rect 16724 5720 16730 5732
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 15804 5664 16037 5692
rect 15804 5652 15810 5664
rect 16025 5661 16037 5664
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16390 5692 16396 5704
rect 16351 5664 16396 5692
rect 16117 5655 16175 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 16853 5695 16911 5701
rect 16853 5692 16865 5695
rect 16816 5664 16865 5692
rect 16816 5652 16822 5664
rect 16853 5661 16865 5664
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 16942 5652 16948 5704
rect 17000 5692 17006 5704
rect 17037 5695 17095 5701
rect 17037 5692 17049 5695
rect 17000 5664 17049 5692
rect 17000 5652 17006 5664
rect 17037 5661 17049 5664
rect 17083 5661 17095 5695
rect 17678 5692 17684 5704
rect 17639 5664 17684 5692
rect 17037 5655 17095 5661
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 17972 5701 18000 5732
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 18874 5760 18880 5772
rect 18196 5732 18880 5760
rect 18196 5720 18202 5732
rect 18874 5720 18880 5732
rect 18932 5760 18938 5772
rect 19150 5760 19156 5772
rect 18932 5732 19156 5760
rect 18932 5720 18938 5732
rect 19150 5720 19156 5732
rect 19208 5760 19214 5772
rect 19996 5760 20024 5791
rect 20346 5788 20352 5840
rect 20404 5828 20410 5840
rect 20993 5831 21051 5837
rect 20993 5828 21005 5831
rect 20404 5800 21005 5828
rect 20404 5788 20410 5800
rect 20993 5797 21005 5800
rect 21039 5797 21051 5831
rect 20993 5791 21051 5797
rect 19208 5732 20024 5760
rect 19208 5720 19214 5732
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20588 5732 20913 5760
rect 20588 5720 20594 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17828 5664 17877 5692
rect 17828 5652 17834 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 17957 5695 18015 5701
rect 17957 5661 17969 5695
rect 18003 5661 18015 5695
rect 17957 5655 18015 5661
rect 18046 5652 18052 5704
rect 18104 5692 18110 5704
rect 18104 5664 18149 5692
rect 18104 5652 18110 5664
rect 19610 5652 19616 5704
rect 19668 5692 19674 5704
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19668 5664 19717 5692
rect 19668 5652 19674 5664
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5661 19947 5695
rect 19889 5655 19947 5661
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20438 5692 20444 5704
rect 20211 5664 20444 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 18414 5624 18420 5636
rect 14844 5596 18420 5624
rect 18414 5584 18420 5596
rect 18472 5624 18478 5636
rect 19904 5624 19932 5655
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 21100 5701 21128 5868
rect 20809 5695 20867 5701
rect 20809 5692 20821 5695
rect 20680 5664 20821 5692
rect 20680 5652 20686 5664
rect 20809 5661 20821 5664
rect 20855 5661 20867 5695
rect 20809 5655 20867 5661
rect 21085 5695 21143 5701
rect 21085 5661 21097 5695
rect 21131 5661 21143 5695
rect 21085 5655 21143 5661
rect 18472 5596 19932 5624
rect 18472 5584 18478 5596
rect 20346 5584 20352 5636
rect 20404 5624 20410 5636
rect 20640 5624 20668 5652
rect 20404 5596 20668 5624
rect 20404 5584 20410 5596
rect 12897 5559 12955 5565
rect 12897 5525 12909 5559
rect 12943 5525 12955 5559
rect 12897 5519 12955 5525
rect 13446 5516 13452 5568
rect 13504 5556 13510 5568
rect 16850 5556 16856 5568
rect 13504 5528 16856 5556
rect 13504 5516 13510 5528
rect 16850 5516 16856 5528
rect 16908 5556 16914 5568
rect 18138 5556 18144 5568
rect 16908 5528 18144 5556
rect 16908 5516 16914 5528
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18325 5559 18383 5565
rect 18325 5525 18337 5559
rect 18371 5556 18383 5559
rect 19518 5556 19524 5568
rect 18371 5528 19524 5556
rect 18371 5525 18383 5528
rect 18325 5519 18383 5525
rect 19518 5516 19524 5528
rect 19576 5516 19582 5568
rect 20622 5556 20628 5568
rect 20583 5528 20628 5556
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 1104 5466 22976 5488
rect 1104 5414 6378 5466
rect 6430 5414 6442 5466
rect 6494 5414 6506 5466
rect 6558 5414 6570 5466
rect 6622 5414 6634 5466
rect 6686 5414 11806 5466
rect 11858 5414 11870 5466
rect 11922 5414 11934 5466
rect 11986 5414 11998 5466
rect 12050 5414 12062 5466
rect 12114 5414 17234 5466
rect 17286 5414 17298 5466
rect 17350 5414 17362 5466
rect 17414 5414 17426 5466
rect 17478 5414 17490 5466
rect 17542 5414 22662 5466
rect 22714 5414 22726 5466
rect 22778 5414 22790 5466
rect 22842 5414 22854 5466
rect 22906 5414 22918 5466
rect 22970 5414 22976 5466
rect 1104 5392 22976 5414
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 4488 5324 4537 5352
rect 4488 5312 4494 5324
rect 4525 5321 4537 5324
rect 4571 5321 4583 5355
rect 4525 5315 4583 5321
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4798 5352 4804 5364
rect 4755 5324 4804 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5166 5352 5172 5364
rect 5127 5324 5172 5352
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8662 5352 8668 5364
rect 7883 5324 8668 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12768 5324 12909 5352
rect 12768 5312 12774 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 13998 5312 14004 5364
rect 14056 5352 14062 5364
rect 14093 5355 14151 5361
rect 14093 5352 14105 5355
rect 14056 5324 14105 5352
rect 14056 5312 14062 5324
rect 14093 5321 14105 5324
rect 14139 5321 14151 5355
rect 14093 5315 14151 5321
rect 18785 5355 18843 5361
rect 18785 5321 18797 5355
rect 18831 5352 18843 5355
rect 18966 5352 18972 5364
rect 18831 5324 18972 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 19242 5352 19248 5364
rect 19203 5324 19248 5352
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 5321 5287 5379 5293
rect 5321 5284 5333 5287
rect 4356 5256 5333 5284
rect 1848 5219 1906 5225
rect 1848 5185 1860 5219
rect 1894 5216 1906 5219
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 1894 5188 3433 5216
rect 1894 5185 1906 5188
rect 1848 5179 1906 5185
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3568 5188 3617 5216
rect 3568 5176 3574 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 4062 5216 4068 5228
rect 3605 5179 3663 5185
rect 3804 5188 4068 5216
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 3326 5108 3332 5160
rect 3384 5148 3390 5160
rect 3804 5148 3832 5188
rect 4062 5176 4068 5188
rect 4120 5216 4126 5228
rect 4356 5225 4384 5256
rect 5321 5253 5333 5256
rect 5367 5253 5379 5287
rect 5321 5247 5379 5253
rect 5537 5287 5595 5293
rect 5537 5253 5549 5287
rect 5583 5253 5595 5287
rect 7006 5284 7012 5296
rect 5537 5247 5595 5253
rect 6564 5256 7012 5284
rect 4341 5219 4399 5225
rect 4341 5216 4353 5219
rect 4120 5188 4353 5216
rect 4120 5176 4126 5188
rect 4341 5185 4353 5188
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4488 5188 4533 5216
rect 4488 5176 4494 5188
rect 3384 5120 3832 5148
rect 3881 5151 3939 5157
rect 3384 5108 3390 5120
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4522 5148 4528 5160
rect 3927 5120 4528 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 2961 5083 3019 5089
rect 2961 5049 2973 5083
rect 3007 5080 3019 5083
rect 3896 5080 3924 5111
rect 4522 5108 4528 5120
rect 4580 5148 4586 5160
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 4580 5120 4721 5148
rect 4580 5108 4586 5120
rect 4709 5117 4721 5120
rect 4755 5148 4767 5151
rect 5552 5148 5580 5247
rect 6564 5225 6592 5256
rect 7006 5244 7012 5256
rect 7064 5244 7070 5296
rect 8972 5287 9030 5293
rect 8972 5253 8984 5287
rect 9018 5284 9030 5287
rect 13541 5287 13599 5293
rect 9018 5256 12434 5284
rect 9018 5253 9030 5256
rect 8972 5247 9030 5253
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7282 5216 7288 5228
rect 6779 5188 7288 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 10036 5219 10094 5225
rect 10036 5185 10048 5219
rect 10082 5216 10094 5219
rect 11698 5216 11704 5228
rect 10082 5188 11704 5216
rect 10082 5185 10094 5188
rect 10036 5179 10094 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 4755 5120 5580 5148
rect 9217 5151 9275 5157
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 9217 5117 9229 5151
rect 9263 5148 9275 5151
rect 9490 5148 9496 5160
rect 9263 5120 9496 5148
rect 9263 5117 9275 5120
rect 9217 5111 9275 5117
rect 9490 5108 9496 5120
rect 9548 5148 9554 5160
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9548 5120 9781 5148
rect 9548 5108 9554 5120
rect 9769 5117 9781 5120
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 3007 5052 3924 5080
rect 12406 5080 12434 5256
rect 13541 5253 13553 5287
rect 13587 5284 13599 5287
rect 13814 5284 13820 5296
rect 13587 5256 13820 5284
rect 13587 5253 13599 5256
rect 13541 5247 13599 5253
rect 13814 5244 13820 5256
rect 13872 5284 13878 5296
rect 15010 5284 15016 5296
rect 13872 5256 15016 5284
rect 13872 5244 13878 5256
rect 15010 5244 15016 5256
rect 15068 5244 15074 5296
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 16390 5284 16396 5296
rect 16347 5256 16396 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 16758 5244 16764 5296
rect 16816 5284 16822 5296
rect 17678 5284 17684 5296
rect 16816 5256 17684 5284
rect 16816 5244 16822 5256
rect 17678 5244 17684 5256
rect 17736 5284 17742 5296
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 17736 5256 17785 5284
rect 17736 5244 17742 5256
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 19794 5284 19800 5296
rect 19755 5256 19800 5284
rect 17773 5247 17831 5253
rect 19794 5244 19800 5256
rect 19852 5244 19858 5296
rect 19889 5287 19947 5293
rect 19889 5253 19901 5287
rect 19935 5284 19947 5287
rect 20622 5284 20628 5296
rect 19935 5256 20628 5284
rect 19935 5253 19947 5256
rect 19889 5247 19947 5253
rect 20622 5244 20628 5256
rect 20680 5244 20686 5296
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 13044 5188 13093 5216
rect 13044 5176 13050 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5216 13231 5219
rect 13262 5216 13268 5228
rect 13219 5188 13268 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14424 5188 14473 5216
rect 14424 5176 14430 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 15194 5216 15200 5228
rect 14599 5188 15200 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 15838 5176 15844 5228
rect 15896 5216 15902 5228
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15896 5188 16037 5216
rect 15896 5176 15902 5188
rect 16025 5185 16037 5188
rect 16071 5216 16083 5219
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 16071 5188 17601 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 17589 5185 17601 5188
rect 17635 5185 17647 5219
rect 17589 5179 17647 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 18196 5188 18245 5216
rect 18196 5176 18202 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18506 5216 18512 5228
rect 18467 5188 18512 5216
rect 18233 5179 18291 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19392 5188 19441 5216
rect 19392 5176 19398 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 19576 5188 19621 5216
rect 19576 5176 19582 5188
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 14274 5148 14280 5160
rect 13495 5120 14280 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5148 14795 5151
rect 15010 5148 15016 5160
rect 14783 5120 15016 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15010 5108 15016 5120
rect 15068 5148 15074 5160
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 15068 5120 17417 5148
rect 15068 5108 15074 5120
rect 17405 5117 17417 5120
rect 17451 5148 17463 5151
rect 17678 5148 17684 5160
rect 17451 5120 17684 5148
rect 17451 5117 17463 5120
rect 17405 5111 17463 5117
rect 17678 5108 17684 5120
rect 17736 5148 17742 5160
rect 18782 5148 18788 5160
rect 17736 5120 18788 5148
rect 17736 5108 17742 5120
rect 18782 5108 18788 5120
rect 18840 5108 18846 5160
rect 18598 5080 18604 5092
rect 12406 5052 18604 5080
rect 3007 5049 3019 5052
rect 2961 5043 3019 5049
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 3142 4972 3148 5024
rect 3200 5012 3206 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3200 4984 3801 5012
rect 3200 4972 3206 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3789 4975 3847 4981
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 5166 5012 5172 5024
rect 4304 4984 5172 5012
rect 4304 4972 4310 4984
rect 5166 4972 5172 4984
rect 5224 5012 5230 5024
rect 5353 5015 5411 5021
rect 5353 5012 5365 5015
rect 5224 4984 5365 5012
rect 5224 4972 5230 4984
rect 5353 4981 5365 4984
rect 5399 4981 5411 5015
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 5353 4975 5411 4981
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 6972 4984 7297 5012
rect 6972 4972 6978 4984
rect 7285 4981 7297 4984
rect 7331 5012 7343 5015
rect 7558 5012 7564 5024
rect 7331 4984 7564 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 16945 5015 17003 5021
rect 16945 4981 16957 5015
rect 16991 5012 17003 5015
rect 17770 5012 17776 5024
rect 16991 4984 17776 5012
rect 16991 4981 17003 4984
rect 16945 4975 17003 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 18782 5012 18788 5024
rect 18555 4984 18788 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 18782 4972 18788 4984
rect 18840 5012 18846 5024
rect 19058 5012 19064 5024
rect 18840 4984 19064 5012
rect 18840 4972 18846 4984
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 1104 4922 22816 4944
rect 1104 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 9092 4922
rect 9144 4870 9156 4922
rect 9208 4870 9220 4922
rect 9272 4870 9284 4922
rect 9336 4870 9348 4922
rect 9400 4870 14520 4922
rect 14572 4870 14584 4922
rect 14636 4870 14648 4922
rect 14700 4870 14712 4922
rect 14764 4870 14776 4922
rect 14828 4870 19948 4922
rect 20000 4870 20012 4922
rect 20064 4870 20076 4922
rect 20128 4870 20140 4922
rect 20192 4870 20204 4922
rect 20256 4870 22816 4922
rect 1104 4848 22816 4870
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7340 4780 7389 4808
rect 7340 4768 7346 4780
rect 7377 4777 7389 4780
rect 7423 4808 7435 4811
rect 7466 4808 7472 4820
rect 7423 4780 7472 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 13538 4808 13544 4820
rect 13499 4780 13544 4808
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 14240 4780 14289 4808
rect 14240 4768 14246 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 14277 4771 14335 4777
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 16022 4808 16028 4820
rect 15983 4780 16028 4808
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 16666 4768 16672 4820
rect 16724 4808 16730 4820
rect 16761 4811 16819 4817
rect 16761 4808 16773 4811
rect 16724 4780 16773 4808
rect 16724 4768 16730 4780
rect 16761 4777 16773 4780
rect 16807 4777 16819 4811
rect 17954 4808 17960 4820
rect 17915 4780 17960 4808
rect 16761 4771 16819 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18693 4811 18751 4817
rect 18693 4808 18705 4811
rect 18472 4780 18705 4808
rect 18472 4768 18478 4780
rect 18693 4777 18705 4780
rect 18739 4777 18751 4811
rect 18693 4771 18751 4777
rect 19429 4811 19487 4817
rect 19429 4777 19441 4811
rect 19475 4808 19487 4811
rect 20438 4808 20444 4820
rect 19475 4780 20444 4808
rect 19475 4777 19487 4780
rect 19429 4771 19487 4777
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 3234 4700 3240 4752
rect 3292 4740 3298 4752
rect 3973 4743 4031 4749
rect 3973 4740 3985 4743
rect 3292 4712 3985 4740
rect 3292 4700 3298 4712
rect 3973 4709 3985 4712
rect 4019 4709 4031 4743
rect 15010 4740 15016 4752
rect 3973 4703 4031 4709
rect 14660 4712 15016 4740
rect 5994 4672 6000 4684
rect 5955 4644 6000 4672
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11698 4672 11704 4684
rect 11204 4644 11704 4672
rect 11204 4632 11210 4644
rect 11698 4632 11704 4644
rect 11756 4672 11762 4684
rect 14366 4672 14372 4684
rect 11756 4644 14372 4672
rect 11756 4632 11762 4644
rect 14366 4632 14372 4644
rect 14424 4672 14430 4684
rect 14424 4644 14596 4672
rect 14424 4632 14430 4644
rect 4246 4604 4252 4616
rect 4207 4576 4252 4604
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 6012 4604 6040 4632
rect 6822 4604 6828 4616
rect 6012 4576 6828 4604
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13814 4604 13820 4616
rect 13771 4576 13820 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14568 4613 14596 4644
rect 14660 4613 14688 4712
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 17862 4740 17868 4752
rect 17420 4712 17868 4740
rect 15194 4672 15200 4684
rect 14752 4644 15200 4672
rect 14752 4613 14780 4644
rect 15194 4632 15200 4644
rect 15252 4672 15258 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15252 4644 15485 4672
rect 15252 4632 15258 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 14553 4607 14611 4613
rect 14553 4573 14565 4607
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4573 14703 4607
rect 14645 4567 14703 4573
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4573 14795 4607
rect 14737 4567 14795 4573
rect 14826 4564 14832 4616
rect 14884 4604 14890 4616
rect 14921 4607 14979 4613
rect 14921 4604 14933 4607
rect 14884 4576 14933 4604
rect 14884 4564 14890 4576
rect 14921 4573 14933 4576
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16577 4607 16635 4613
rect 16577 4604 16589 4607
rect 16448 4576 16589 4604
rect 16448 4564 16454 4576
rect 16577 4573 16589 4576
rect 16623 4573 16635 4607
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 16577 4567 16635 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 17420 4613 17448 4712
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 18506 4632 18512 4684
rect 18564 4672 18570 4684
rect 18564 4644 18920 4672
rect 18564 4632 18570 4644
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17405 4567 17463 4573
rect 17678 4564 17684 4616
rect 17736 4604 17742 4616
rect 17865 4607 17923 4613
rect 17865 4604 17877 4607
rect 17736 4576 17877 4604
rect 17736 4564 17742 4576
rect 17865 4573 17877 4576
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4573 18107 4607
rect 18690 4604 18696 4616
rect 18651 4576 18696 4604
rect 18049 4567 18107 4573
rect 3510 4496 3516 4548
rect 3568 4536 3574 4548
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 3568 4508 3985 4536
rect 3568 4496 3574 4508
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 3973 4499 4031 4505
rect 6264 4539 6322 4545
rect 6264 4505 6276 4539
rect 6310 4536 6322 4539
rect 6546 4536 6552 4548
rect 6310 4508 6552 4536
rect 6310 4505 6322 4508
rect 6264 4499 6322 4505
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 15841 4539 15899 4545
rect 15841 4536 15853 4539
rect 11112 4508 15853 4536
rect 11112 4496 11118 4508
rect 15841 4505 15853 4508
rect 15887 4536 15899 4539
rect 17313 4539 17371 4545
rect 17313 4536 17325 4539
rect 15887 4508 17325 4536
rect 15887 4505 15899 4508
rect 15841 4499 15899 4505
rect 17313 4505 17325 4508
rect 17359 4505 17371 4539
rect 18064 4536 18092 4567
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 18892 4613 18920 4644
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19334 4536 19340 4548
rect 18064 4508 19340 4536
rect 17313 4499 17371 4505
rect 19334 4496 19340 4508
rect 19392 4496 19398 4548
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 5350 4468 5356 4480
rect 4203 4440 5356 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 5534 4468 5540 4480
rect 5495 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 14182 4468 14188 4480
rect 7616 4440 14188 4468
rect 7616 4428 7622 4440
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 19444 4468 19472 4567
rect 19518 4564 19524 4616
rect 19576 4604 19582 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 19576 4576 19625 4604
rect 19576 4564 19582 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 18380 4440 19472 4468
rect 18380 4428 18386 4440
rect 1104 4378 22976 4400
rect 1104 4326 6378 4378
rect 6430 4326 6442 4378
rect 6494 4326 6506 4378
rect 6558 4326 6570 4378
rect 6622 4326 6634 4378
rect 6686 4326 11806 4378
rect 11858 4326 11870 4378
rect 11922 4326 11934 4378
rect 11986 4326 11998 4378
rect 12050 4326 12062 4378
rect 12114 4326 17234 4378
rect 17286 4326 17298 4378
rect 17350 4326 17362 4378
rect 17414 4326 17426 4378
rect 17478 4326 17490 4378
rect 17542 4326 22662 4378
rect 22714 4326 22726 4378
rect 22778 4326 22790 4378
rect 22842 4326 22854 4378
rect 22906 4326 22918 4378
rect 22970 4326 22976 4378
rect 1104 4304 22976 4326
rect 15194 4224 15200 4276
rect 15252 4264 15258 4276
rect 15381 4267 15439 4273
rect 15381 4264 15393 4267
rect 15252 4236 15393 4264
rect 15252 4224 15258 4236
rect 15381 4233 15393 4236
rect 15427 4233 15439 4267
rect 15381 4227 15439 4233
rect 17681 4267 17739 4273
rect 17681 4233 17693 4267
rect 17727 4264 17739 4267
rect 18138 4264 18144 4276
rect 17727 4236 18144 4264
rect 17727 4233 17739 4236
rect 17681 4227 17739 4233
rect 18138 4224 18144 4236
rect 18196 4264 18202 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 18196 4236 18981 4264
rect 18196 4224 18202 4236
rect 18969 4233 18981 4236
rect 19015 4233 19027 4267
rect 18969 4227 19027 4233
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 14001 4199 14059 4205
rect 6972 4168 9260 4196
rect 6972 4156 6978 4168
rect 2676 4131 2734 4137
rect 2676 4097 2688 4131
rect 2722 4128 2734 4131
rect 3050 4128 3056 4140
rect 2722 4100 3056 4128
rect 2722 4097 2734 4100
rect 2676 4091 2734 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 4614 4128 4620 4140
rect 4575 4100 4620 4128
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4884 4131 4942 4137
rect 4884 4097 4896 4131
rect 4930 4128 4942 4131
rect 6086 4128 6092 4140
rect 4930 4100 6092 4128
rect 4930 4097 4942 4100
rect 4884 4091 4942 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7101 4131 7159 4137
rect 7101 4128 7113 4131
rect 7064 4100 7113 4128
rect 7064 4088 7070 4100
rect 7101 4097 7113 4100
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 8018 4128 8024 4140
rect 7423 4100 8024 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8938 4128 8944 4140
rect 8996 4137 9002 4140
rect 9232 4137 9260 4168
rect 14001 4165 14013 4199
rect 14047 4196 14059 4199
rect 14826 4196 14832 4208
rect 14047 4168 14832 4196
rect 14047 4165 14059 4168
rect 14001 4159 14059 4165
rect 8908 4100 8944 4128
rect 8938 4088 8944 4100
rect 8996 4091 9008 4137
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9490 4128 9496 4140
rect 9263 4100 9496 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 8996 4088 9002 4091
rect 9490 4088 9496 4100
rect 9548 4128 9554 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9548 4100 9689 4128
rect 9548 4088 9554 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9944 4131 10002 4137
rect 9944 4097 9956 4131
rect 9990 4128 10002 4131
rect 11054 4128 11060 4140
rect 9990 4100 11060 4128
rect 9990 4097 10002 4100
rect 9944 4091 10002 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4128 12127 4131
rect 12158 4128 12164 4140
rect 12115 4100 12164 4128
rect 12115 4097 12127 4100
rect 12069 4091 12127 4097
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12986 4128 12992 4140
rect 12947 4100 12992 4128
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 1636 4032 2421 4060
rect 1636 4020 1642 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 13078 4060 13084 4072
rect 13039 4032 13084 4060
rect 2409 4023 2467 4029
rect 2424 3924 2452 4023
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 7282 3992 7288 4004
rect 7243 3964 7288 3992
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 13170 3992 13176 4004
rect 12299 3964 13176 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 13357 3995 13415 4001
rect 13357 3961 13369 3995
rect 13403 3992 13415 3995
rect 14016 3992 14044 4159
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 18984 4196 19012 4227
rect 18984 4168 19196 4196
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 15562 4128 15568 4140
rect 14240 4100 14333 4128
rect 15523 4100 15568 4128
rect 14240 4088 14246 4100
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 15746 4128 15752 4140
rect 15707 4100 15752 4128
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 16482 4128 16488 4140
rect 15887 4100 16488 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 16482 4088 16488 4100
rect 16540 4128 16546 4140
rect 16942 4128 16948 4140
rect 16540 4100 16948 4128
rect 16540 4088 16546 4100
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17313 4131 17371 4137
rect 17313 4128 17325 4131
rect 17092 4100 17325 4128
rect 17092 4088 17098 4100
rect 17313 4097 17325 4100
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17770 4128 17776 4140
rect 17543 4100 17776 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 14200 4060 14228 4088
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14200 4032 14933 4060
rect 14921 4029 14933 4032
rect 14967 4060 14979 4063
rect 17512 4060 17540 4091
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18972 4131 19030 4137
rect 18972 4128 18984 4131
rect 17920 4100 18984 4128
rect 17920 4088 17926 4100
rect 18972 4097 18984 4100
rect 19018 4128 19030 4131
rect 19168 4128 19196 4168
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19018 4100 19104 4128
rect 19168 4100 19625 4128
rect 19018 4097 19030 4100
rect 18972 4091 19030 4097
rect 18506 4060 18512 4072
rect 14967 4032 17540 4060
rect 18467 4032 18512 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 13403 3964 14044 3992
rect 13403 3961 13415 3964
rect 13357 3955 13415 3961
rect 15746 3952 15752 4004
rect 15804 3992 15810 4004
rect 18414 3992 18420 4004
rect 15804 3964 18420 3992
rect 15804 3952 15810 3964
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 19076 3992 19104 4100
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 19797 4131 19855 4137
rect 19797 4097 19809 4131
rect 19843 4097 19855 4131
rect 19797 4091 19855 4097
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19705 4063 19763 4069
rect 19705 4060 19717 4063
rect 19392 4032 19717 4060
rect 19392 4020 19398 4032
rect 19705 4029 19717 4032
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 19812 3992 19840 4091
rect 19076 3964 19840 3992
rect 2682 3924 2688 3936
rect 2424 3896 2688 3924
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 3510 3884 3516 3936
rect 3568 3924 3574 3936
rect 3789 3927 3847 3933
rect 3789 3924 3801 3927
rect 3568 3896 3801 3924
rect 3568 3884 3574 3896
rect 3789 3893 3801 3896
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 5902 3924 5908 3936
rect 4120 3896 5908 3924
rect 4120 3884 4126 3896
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6546 3924 6552 3936
rect 6043 3896 6552 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 7156 3896 7205 3924
rect 7156 3884 7162 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7834 3924 7840 3936
rect 7795 3896 7840 3924
rect 7193 3887 7251 3893
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 11057 3927 11115 3933
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 12066 3924 12072 3936
rect 11103 3896 12072 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 12066 3884 12072 3896
rect 12124 3924 12130 3936
rect 13262 3924 13268 3936
rect 12124 3896 13268 3924
rect 12124 3884 12130 3896
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 13964 3896 14289 3924
rect 13964 3884 13970 3896
rect 14277 3893 14289 3896
rect 14323 3893 14335 3927
rect 14277 3887 14335 3893
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 17310 3924 17316 3936
rect 15160 3896 17316 3924
rect 15160 3884 15166 3896
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18601 3927 18659 3933
rect 18601 3924 18613 3927
rect 18380 3896 18613 3924
rect 18380 3884 18386 3896
rect 18601 3893 18613 3896
rect 18647 3893 18659 3927
rect 18601 3887 18659 3893
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3924 19211 3927
rect 20530 3924 20536 3936
rect 19199 3896 20536 3924
rect 19199 3893 19211 3896
rect 19153 3887 19211 3893
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 1104 3834 22816 3856
rect 1104 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 9092 3834
rect 9144 3782 9156 3834
rect 9208 3782 9220 3834
rect 9272 3782 9284 3834
rect 9336 3782 9348 3834
rect 9400 3782 14520 3834
rect 14572 3782 14584 3834
rect 14636 3782 14648 3834
rect 14700 3782 14712 3834
rect 14764 3782 14776 3834
rect 14828 3782 19948 3834
rect 20000 3782 20012 3834
rect 20064 3782 20076 3834
rect 20128 3782 20140 3834
rect 20192 3782 20204 3834
rect 20256 3782 22816 3834
rect 1104 3760 22816 3782
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3142 3720 3148 3732
rect 3099 3692 3148 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 4522 3720 4528 3732
rect 4172 3692 4528 3720
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 4172 3593 4200 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5408 3692 5549 3720
rect 5408 3680 5414 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 6086 3720 6092 3732
rect 6047 3692 6092 3720
rect 5537 3683 5595 3689
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 7282 3720 7288 3732
rect 6503 3692 7288 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 13078 3720 13084 3732
rect 12492 3692 13084 3720
rect 12492 3680 12498 3692
rect 13078 3680 13084 3692
rect 13136 3720 13142 3732
rect 14369 3723 14427 3729
rect 14369 3720 14381 3723
rect 13136 3692 14381 3720
rect 13136 3680 13142 3692
rect 14369 3689 14381 3692
rect 14415 3689 14427 3723
rect 14369 3683 14427 3689
rect 14737 3723 14795 3729
rect 14737 3689 14749 3723
rect 14783 3720 14795 3723
rect 14918 3720 14924 3732
rect 14783 3692 14924 3720
rect 14783 3689 14795 3692
rect 14737 3683 14795 3689
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 16577 3723 16635 3729
rect 16577 3689 16589 3723
rect 16623 3720 16635 3723
rect 17034 3720 17040 3732
rect 16623 3692 17040 3720
rect 16623 3689 16635 3692
rect 16577 3683 16635 3689
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 19613 3723 19671 3729
rect 17368 3692 19472 3720
rect 17368 3680 17374 3692
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 11885 3655 11943 3661
rect 11885 3652 11897 3655
rect 11756 3624 11897 3652
rect 11756 3612 11762 3624
rect 11885 3621 11897 3624
rect 11931 3652 11943 3655
rect 15286 3652 15292 3664
rect 11931 3624 12434 3652
rect 11931 3621 11943 3624
rect 11885 3615 11943 3621
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 2740 3556 4169 3584
rect 2740 3544 2746 3556
rect 4157 3553 4169 3556
rect 4203 3553 4215 3587
rect 6546 3584 6552 3596
rect 6507 3556 6552 3584
rect 4157 3547 4215 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6972 3556 7021 3584
rect 6972 3544 6978 3556
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9548 3556 9965 3584
rect 9548 3544 9554 3556
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 12406 3584 12434 3624
rect 13280 3624 15292 3652
rect 12989 3587 13047 3593
rect 12989 3584 13001 3587
rect 12406 3556 13001 3584
rect 9953 3547 10011 3553
rect 12989 3553 13001 3556
rect 13035 3553 13047 3587
rect 12989 3547 13047 3553
rect 13078 3544 13084 3596
rect 13136 3584 13142 3596
rect 13280 3593 13308 3624
rect 15286 3612 15292 3624
rect 15344 3612 15350 3664
rect 15838 3652 15844 3664
rect 15799 3624 15844 3652
rect 15838 3612 15844 3624
rect 15896 3652 15902 3664
rect 18322 3652 18328 3664
rect 15896 3624 18328 3652
rect 15896 3612 15902 3624
rect 18322 3612 18328 3624
rect 18380 3612 18386 3664
rect 18414 3612 18420 3664
rect 18472 3652 18478 3664
rect 18601 3655 18659 3661
rect 18601 3652 18613 3655
rect 18472 3624 18613 3652
rect 18472 3612 18478 3624
rect 18601 3621 18613 3624
rect 18647 3621 18659 3655
rect 18601 3615 18659 3621
rect 13265 3587 13323 3593
rect 13136 3556 13181 3584
rect 13136 3544 13142 3556
rect 13265 3553 13277 3587
rect 13311 3553 13323 3587
rect 13265 3547 13323 3553
rect 13449 3587 13507 3593
rect 13449 3553 13461 3587
rect 13495 3584 13507 3587
rect 13495 3556 13676 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3326 3516 3332 3528
rect 3283 3488 3332 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 5166 3516 5172 3528
rect 3467 3488 5172 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 6270 3516 6276 3528
rect 6231 3488 6276 3516
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7265 3519 7323 3525
rect 7265 3516 7277 3519
rect 7156 3488 7277 3516
rect 7156 3476 7162 3488
rect 7265 3485 7277 3488
rect 7311 3485 7323 3519
rect 7265 3479 7323 3485
rect 10220 3519 10278 3525
rect 10220 3485 10232 3519
rect 10266 3516 10278 3519
rect 12176 3516 12296 3518
rect 12342 3516 12348 3528
rect 10266 3488 11468 3516
rect 10266 3485 10278 3488
rect 10220 3479 10278 3485
rect 4424 3451 4482 3457
rect 4424 3417 4436 3451
rect 4470 3448 4482 3451
rect 4798 3448 4804 3460
rect 4470 3420 4804 3448
rect 4470 3417 4482 3420
rect 4424 3411 4482 3417
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 11054 3448 11060 3460
rect 5592 3420 11060 3448
rect 5592 3408 5598 3420
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 8110 3380 8116 3392
rect 7248 3352 8116 3380
rect 7248 3340 7254 3352
rect 8110 3340 8116 3352
rect 8168 3380 8174 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 8168 3352 8401 3380
rect 8168 3340 8174 3352
rect 8389 3349 8401 3352
rect 8435 3349 8447 3383
rect 8389 3343 8447 3349
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11333 3383 11391 3389
rect 11333 3380 11345 3383
rect 11204 3352 11345 3380
rect 11204 3340 11210 3352
rect 11333 3349 11345 3352
rect 11379 3349 11391 3383
rect 11440 3380 11468 3488
rect 12176 3490 12348 3516
rect 12066 3448 12072 3460
rect 12027 3420 12072 3448
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12176 3457 12204 3490
rect 12268 3488 12348 3490
rect 12342 3476 12348 3488
rect 12400 3516 12406 3528
rect 13173 3519 13231 3525
rect 13173 3516 13185 3519
rect 12400 3488 13185 3516
rect 12400 3476 12406 3488
rect 13173 3485 13185 3488
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 12161 3451 12219 3457
rect 12161 3417 12173 3451
rect 12207 3417 12219 3451
rect 12161 3411 12219 3417
rect 12253 3451 12311 3457
rect 12253 3417 12265 3451
rect 12299 3448 12311 3451
rect 12299 3420 12756 3448
rect 12299 3417 12311 3420
rect 12253 3411 12311 3417
rect 12618 3380 12624 3392
rect 11440 3352 12624 3380
rect 11333 3343 11391 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12728 3380 12756 3420
rect 13280 3380 13308 3547
rect 13648 3528 13676 3556
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 15194 3584 15200 3596
rect 13780 3556 15200 3584
rect 13780 3544 13786 3556
rect 15194 3544 15200 3556
rect 15252 3544 15258 3596
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3584 16543 3587
rect 16850 3584 16856 3596
rect 16531 3556 16856 3584
rect 16531 3553 16543 3556
rect 16485 3547 16543 3553
rect 16850 3544 16856 3556
rect 16908 3584 16914 3596
rect 16908 3556 17540 3584
rect 16908 3544 16914 3556
rect 13630 3516 13636 3528
rect 13543 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13688 3488 14289 3516
rect 13688 3476 13694 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 15102 3516 15108 3528
rect 14424 3488 15108 3516
rect 14424 3476 14430 3488
rect 15102 3476 15108 3488
rect 15160 3516 15166 3528
rect 15473 3519 15531 3525
rect 15473 3516 15485 3519
rect 15160 3488 15485 3516
rect 15160 3476 15166 3488
rect 15473 3485 15485 3488
rect 15519 3485 15531 3519
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 15473 3479 15531 3485
rect 15672 3488 16589 3516
rect 15672 3457 15700 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17512 3525 17540 3556
rect 17497 3519 17555 3525
rect 17000 3488 17448 3516
rect 17000 3476 17006 3488
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3417 15715 3451
rect 15657 3411 15715 3417
rect 12728 3352 13308 3380
rect 15672 3380 15700 3411
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 15988 3420 16313 3448
rect 15988 3408 15994 3420
rect 16301 3417 16313 3420
rect 16347 3448 16359 3451
rect 17313 3451 17371 3457
rect 17313 3448 17325 3451
rect 16347 3420 17325 3448
rect 16347 3417 16359 3420
rect 16301 3411 16359 3417
rect 17313 3417 17325 3420
rect 17359 3417 17371 3451
rect 17420 3448 17448 3488
rect 17497 3485 17509 3519
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18340 3525 18368 3612
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3584 18567 3587
rect 19334 3584 19340 3596
rect 18555 3556 19340 3584
rect 18555 3553 18567 3556
rect 18509 3547 18567 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17920 3488 18153 3516
rect 17920 3476 17926 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18524 3516 18736 3518
rect 18874 3516 18880 3528
rect 18463 3490 18880 3516
rect 18463 3488 18552 3490
rect 18708 3488 18880 3490
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 19444 3525 19472 3692
rect 19613 3689 19625 3723
rect 19659 3689 19671 3723
rect 19613 3683 19671 3689
rect 19518 3612 19524 3664
rect 19576 3612 19582 3664
rect 19628 3652 19656 3683
rect 19702 3680 19708 3732
rect 19760 3720 19766 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19760 3692 19809 3720
rect 19760 3680 19766 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19797 3683 19855 3689
rect 20254 3652 20260 3664
rect 19628 3624 19748 3652
rect 20215 3624 20260 3652
rect 19536 3584 19564 3612
rect 19720 3584 19748 3624
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 20993 3587 21051 3593
rect 20993 3584 21005 3587
rect 19536 3556 19656 3584
rect 19628 3525 19656 3556
rect 19720 3556 21005 3584
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 17681 3451 17739 3457
rect 17681 3448 17693 3451
rect 17420 3420 17693 3448
rect 17313 3411 17371 3417
rect 17681 3417 17693 3420
rect 17727 3417 17739 3451
rect 17681 3411 17739 3417
rect 17770 3408 17776 3460
rect 17828 3448 17834 3460
rect 19720 3448 19748 3556
rect 20993 3553 21005 3556
rect 21039 3553 21051 3587
rect 20993 3547 21051 3553
rect 20530 3516 20536 3528
rect 20491 3488 20536 3516
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 17828 3420 19748 3448
rect 17828 3408 17834 3420
rect 19978 3408 19984 3460
rect 20036 3448 20042 3460
rect 20257 3451 20315 3457
rect 20257 3448 20269 3451
rect 20036 3420 20269 3448
rect 20036 3408 20042 3420
rect 20257 3417 20269 3420
rect 20303 3417 20315 3451
rect 20257 3411 20315 3417
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 20441 3451 20499 3457
rect 20441 3448 20453 3451
rect 20404 3420 20453 3448
rect 20404 3408 20410 3420
rect 20441 3417 20453 3420
rect 20487 3417 20499 3451
rect 20441 3411 20499 3417
rect 16574 3380 16580 3392
rect 15672 3352 16580 3380
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 16758 3380 16764 3392
rect 16719 3352 16764 3380
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 18874 3380 18880 3392
rect 18835 3352 18880 3380
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 20364 3380 20392 3408
rect 19392 3352 20392 3380
rect 19392 3340 19398 3352
rect 1104 3290 22976 3312
rect 1104 3238 6378 3290
rect 6430 3238 6442 3290
rect 6494 3238 6506 3290
rect 6558 3238 6570 3290
rect 6622 3238 6634 3290
rect 6686 3238 11806 3290
rect 11858 3238 11870 3290
rect 11922 3238 11934 3290
rect 11986 3238 11998 3290
rect 12050 3238 12062 3290
rect 12114 3238 17234 3290
rect 17286 3238 17298 3290
rect 17350 3238 17362 3290
rect 17414 3238 17426 3290
rect 17478 3238 17490 3290
rect 17542 3238 22662 3290
rect 22714 3238 22726 3290
rect 22778 3238 22790 3290
rect 22842 3238 22854 3290
rect 22906 3238 22918 3290
rect 22970 3238 22976 3290
rect 1104 3216 22976 3238
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6788 3148 7113 3176
rect 6788 3136 6794 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7248 3148 7293 3176
rect 7248 3136 7254 3148
rect 8202 3136 8208 3188
rect 8260 3176 8266 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 8260 3148 10241 3176
rect 8260 3136 8266 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12400 3148 14780 3176
rect 12400 3136 12406 3148
rect 2682 3108 2688 3120
rect 2643 3080 2688 3108
rect 2682 3068 2688 3080
rect 2740 3068 2746 3120
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 7374 3108 7380 3120
rect 4387 3080 7380 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 7374 3068 7380 3080
rect 7432 3108 7438 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 7432 3080 7849 3108
rect 7432 3068 7438 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 9490 3108 9496 3120
rect 9451 3080 9496 3108
rect 7837 3071 7895 3077
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 11146 3108 11152 3120
rect 11107 3080 11152 3108
rect 11146 3068 11152 3080
rect 11204 3108 11210 3120
rect 11204 3080 12112 3108
rect 11204 3068 11210 3080
rect 4982 3040 4988 3052
rect 4943 3012 4988 3040
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 5350 3040 5356 3052
rect 5307 3012 5356 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 5951 3012 6837 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7055 3012 7144 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 5184 2972 5212 3000
rect 5721 2975 5779 2981
rect 5721 2972 5733 2975
rect 4856 2944 5733 2972
rect 4856 2932 4862 2944
rect 5721 2941 5733 2944
rect 5767 2941 5779 2975
rect 5721 2935 5779 2941
rect 7116 2916 7144 3012
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 12084 3049 12112 3080
rect 12176 3080 13124 3108
rect 12176 3049 12204 3080
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 7616 3012 10057 3040
rect 7616 3000 7622 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3040 11023 3043
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11011 3012 11989 3040
rect 11011 3009 11023 3012
rect 10965 3003 11023 3009
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12069 3003 12127 3009
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3009 12219 3043
rect 12986 3040 12992 3052
rect 12161 3003 12219 3009
rect 12406 3012 12992 3040
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 7248 2944 7389 2972
rect 7248 2932 7254 2944
rect 7377 2941 7389 2944
rect 7423 2972 7435 2975
rect 7466 2972 7472 2984
rect 7423 2944 7472 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 10336 2972 10364 3003
rect 9548 2944 10364 2972
rect 10888 2972 10916 3003
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 10888 2944 11897 2972
rect 9548 2932 9554 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11992 2972 12020 3003
rect 12406 2972 12434 3012
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13096 2984 13124 3080
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13630 3040 13636 3052
rect 13495 3012 13636 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 14752 3040 14780 3148
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15765 3179 15823 3185
rect 15765 3176 15777 3179
rect 15344 3148 15777 3176
rect 15344 3136 15350 3148
rect 15765 3145 15777 3148
rect 15811 3145 15823 3179
rect 15765 3139 15823 3145
rect 18230 3136 18236 3188
rect 18288 3176 18294 3188
rect 18417 3179 18475 3185
rect 18417 3176 18429 3179
rect 18288 3148 18429 3176
rect 18288 3136 18294 3148
rect 18417 3145 18429 3148
rect 18463 3145 18475 3179
rect 18417 3139 18475 3145
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 18564 3148 19625 3176
rect 18564 3136 18570 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 19613 3139 19671 3145
rect 19702 3136 19708 3188
rect 19760 3176 19766 3188
rect 19978 3176 19984 3188
rect 19760 3148 19984 3176
rect 19760 3136 19766 3148
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 15194 3068 15200 3120
rect 15252 3108 15258 3120
rect 15565 3111 15623 3117
rect 15565 3108 15577 3111
rect 15252 3080 15577 3108
rect 15252 3068 15258 3080
rect 15565 3077 15577 3080
rect 15611 3108 15623 3111
rect 15611 3080 19564 3108
rect 15611 3077 15623 3080
rect 15565 3071 15623 3077
rect 15856 3052 15884 3080
rect 19536 3052 19564 3080
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14752 3012 14933 3040
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 11992 2944 12434 2972
rect 11885 2935 11943 2941
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7834 2904 7840 2916
rect 7156 2876 7840 2904
rect 7156 2864 7162 2876
rect 7834 2864 7840 2876
rect 7892 2904 7898 2916
rect 9508 2904 9536 2932
rect 7892 2876 9536 2904
rect 11900 2904 11928 2935
rect 13078 2932 13084 2984
rect 13136 2972 13142 2984
rect 13173 2975 13231 2981
rect 13173 2972 13185 2975
rect 13136 2944 13185 2972
rect 13136 2932 13142 2944
rect 13173 2941 13185 2944
rect 13219 2941 13231 2975
rect 13173 2935 13231 2941
rect 12434 2904 12440 2916
rect 11900 2876 12440 2904
rect 7892 2864 7898 2876
rect 12434 2864 12440 2876
rect 12492 2904 12498 2916
rect 12492 2876 13124 2904
rect 12492 2864 12498 2876
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 7466 2836 7472 2848
rect 7064 2808 7472 2836
rect 7064 2796 7070 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11698 2836 11704 2848
rect 11659 2808 11704 2836
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 12894 2836 12900 2848
rect 12855 2808 12900 2836
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 13096 2845 13124 2876
rect 14274 2864 14280 2916
rect 14332 2904 14338 2916
rect 14553 2907 14611 2913
rect 14553 2904 14565 2907
rect 14332 2876 14565 2904
rect 14332 2864 14338 2876
rect 14553 2873 14565 2876
rect 14599 2873 14611 2907
rect 14553 2867 14611 2873
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2805 13139 2839
rect 14936 2836 14964 3003
rect 15838 3000 15844 3052
rect 15896 3000 15902 3052
rect 15930 3000 15936 3052
rect 15988 3040 15994 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 15988 3012 16865 3040
rect 15988 3000 15994 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 18690 3040 18696 3052
rect 18651 3012 18696 3040
rect 16853 3003 16911 3009
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2972 15071 2975
rect 15286 2972 15292 2984
rect 15059 2944 15292 2972
rect 15059 2941 15071 2944
rect 15013 2935 15071 2941
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 16942 2972 16948 2984
rect 16632 2944 16948 2972
rect 16632 2932 16638 2944
rect 16942 2932 16948 2944
rect 17000 2972 17006 2984
rect 17681 2975 17739 2981
rect 17681 2972 17693 2975
rect 17000 2944 17693 2972
rect 17000 2932 17006 2944
rect 17681 2941 17693 2944
rect 17727 2941 17739 2975
rect 18800 2972 18828 3003
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 18932 3012 18977 3040
rect 18932 3000 18938 3012
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19116 3012 19161 3040
rect 19116 3000 19122 3012
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19576 3012 19717 3040
rect 19576 3000 19582 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 20254 2972 20260 2984
rect 18800 2944 20260 2972
rect 17681 2935 17739 2941
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 15746 2836 15752 2848
rect 14936 2808 15752 2836
rect 13081 2799 13139 2805
rect 15746 2796 15752 2808
rect 15804 2796 15810 2848
rect 15933 2839 15991 2845
rect 15933 2805 15945 2839
rect 15979 2836 15991 2839
rect 16850 2836 16856 2848
rect 15979 2808 16856 2836
rect 15979 2805 15991 2808
rect 15933 2799 15991 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 17218 2836 17224 2848
rect 17179 2808 17224 2836
rect 17218 2796 17224 2808
rect 17276 2796 17282 2848
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 19334 2836 19340 2848
rect 18656 2808 19340 2836
rect 18656 2796 18662 2808
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 1104 2746 22816 2768
rect 1104 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 9092 2746
rect 9144 2694 9156 2746
rect 9208 2694 9220 2746
rect 9272 2694 9284 2746
rect 9336 2694 9348 2746
rect 9400 2694 14520 2746
rect 14572 2694 14584 2746
rect 14636 2694 14648 2746
rect 14700 2694 14712 2746
rect 14764 2694 14776 2746
rect 14828 2694 19948 2746
rect 20000 2694 20012 2746
rect 20064 2694 20076 2746
rect 20128 2694 20140 2746
rect 20192 2694 20204 2746
rect 20256 2694 22816 2746
rect 1104 2672 22816 2694
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3326 2592 3332 2644
rect 3384 2632 3390 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3384 2604 3985 2632
rect 3384 2592 3390 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 5040 2604 5089 2632
rect 5040 2592 5046 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6270 2632 6276 2644
rect 5767 2604 6276 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 7282 2632 7288 2644
rect 7239 2604 7288 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2601 7435 2635
rect 8018 2632 8024 2644
rect 7979 2604 8024 2632
rect 7377 2595 7435 2601
rect 3142 2564 3148 2576
rect 3103 2536 3148 2564
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 7392 2564 7420 2595
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 8938 2592 8944 2644
rect 8996 2632 9002 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8996 2604 9137 2632
rect 8996 2592 9002 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 9125 2595 9183 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 11054 2632 11060 2644
rect 11015 2604 11060 2632
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12158 2632 12164 2644
rect 12115 2604 12164 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 12713 2635 12771 2641
rect 12713 2601 12725 2635
rect 12759 2632 12771 2635
rect 13078 2632 13084 2644
rect 12759 2604 13084 2632
rect 12759 2601 12771 2604
rect 12713 2595 12771 2601
rect 8110 2564 8116 2576
rect 7392 2536 8116 2564
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 11072 2564 11100 2592
rect 12728 2564 12756 2595
rect 13078 2592 13084 2604
rect 13136 2632 13142 2644
rect 15197 2635 15255 2641
rect 15197 2632 15209 2635
rect 13136 2604 15209 2632
rect 13136 2592 13142 2604
rect 15197 2601 15209 2604
rect 15243 2632 15255 2635
rect 15930 2632 15936 2644
rect 15243 2604 15700 2632
rect 15891 2604 15936 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 11072 2536 12756 2564
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 5350 2496 5356 2508
rect 4387 2468 5356 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3292 2400 3337 2428
rect 3292 2388 3298 2400
rect 3510 2388 3516 2440
rect 3568 2428 3574 2440
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 3568 2400 4169 2428
rect 3568 2388 3574 2400
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4798 2428 4804 2440
rect 4759 2400 4804 2428
rect 4157 2391 4215 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 4908 2437 4936 2468
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 10042 2496 10048 2508
rect 9324 2468 10048 2496
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 4939 2400 4973 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5721 2431 5779 2437
rect 5721 2428 5733 2431
rect 5224 2400 5733 2428
rect 5224 2388 5230 2400
rect 5721 2397 5733 2400
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 7466 2428 7472 2440
rect 5951 2400 7472 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 5077 2363 5135 2369
rect 5077 2360 5089 2363
rect 3007 2332 5089 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 5077 2329 5089 2332
rect 5123 2360 5135 2363
rect 5920 2360 5948 2391
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8110 2428 8116 2440
rect 8067 2400 8116 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 9324 2437 9352 2468
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 15672 2496 15700 2604
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17862 2632 17868 2644
rect 16991 2604 17868 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18601 2635 18659 2641
rect 18601 2601 18613 2635
rect 18647 2632 18659 2635
rect 19702 2632 19708 2644
rect 18647 2604 19708 2632
rect 18647 2601 18659 2604
rect 18601 2595 18659 2601
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 15672 2468 15792 2496
rect 9309 2431 9367 2437
rect 8281 2409 8339 2415
rect 8281 2406 8293 2409
rect 8220 2378 8293 2406
rect 5123 2332 5948 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 7190 2320 7196 2372
rect 7248 2360 7254 2372
rect 7561 2363 7619 2369
rect 7561 2360 7573 2363
rect 7248 2332 7573 2360
rect 7248 2320 7254 2332
rect 7561 2329 7573 2332
rect 7607 2360 7619 2363
rect 7926 2360 7932 2372
rect 7607 2332 7932 2360
rect 7607 2329 7619 2332
rect 7561 2323 7619 2329
rect 7926 2320 7932 2332
rect 7984 2320 7990 2372
rect 8220 2360 8248 2378
rect 8281 2375 8293 2378
rect 8327 2375 8339 2409
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9309 2391 9367 2397
rect 9416 2400 9597 2428
rect 8281 2369 8339 2375
rect 8128 2332 8248 2360
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7361 2295 7419 2301
rect 7361 2292 7373 2295
rect 7156 2264 7373 2292
rect 7156 2252 7162 2264
rect 7361 2261 7373 2264
rect 7407 2292 7419 2295
rect 8128 2292 8156 2332
rect 7407 2264 8156 2292
rect 7407 2261 7419 2264
rect 7361 2255 7419 2261
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 9416 2292 9444 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 11698 2428 11704 2440
rect 11659 2400 11704 2428
rect 9585 2391 9643 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 12952 2400 13369 2428
rect 12952 2388 12958 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 15528 2400 15669 2428
rect 15528 2388 15534 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15764 2428 15792 2468
rect 16022 2456 16028 2508
rect 16080 2496 16086 2508
rect 18598 2496 18604 2508
rect 16080 2468 18604 2496
rect 16080 2456 16086 2468
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 16942 2428 16948 2440
rect 15764 2400 16948 2428
rect 15657 2391 15715 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17218 2428 17224 2440
rect 17083 2400 17224 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 17696 2400 18337 2428
rect 11146 2320 11152 2372
rect 11204 2360 11210 2372
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 11204 2332 11897 2360
rect 11204 2320 11210 2332
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 15746 2360 15752 2372
rect 15707 2332 15752 2360
rect 11885 2323 11943 2329
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 15838 2320 15844 2372
rect 15896 2360 15902 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 15896 2332 15945 2360
rect 15896 2320 15902 2332
rect 15933 2329 15945 2332
rect 15979 2329 15991 2363
rect 16960 2360 16988 2388
rect 17589 2363 17647 2369
rect 17589 2360 17601 2363
rect 16960 2332 17601 2360
rect 15933 2323 15991 2329
rect 17589 2329 17601 2332
rect 17635 2329 17647 2363
rect 17589 2323 17647 2329
rect 8260 2264 9444 2292
rect 13541 2295 13599 2301
rect 8260 2252 8266 2264
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 15562 2292 15568 2304
rect 13587 2264 15568 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 15562 2252 15568 2264
rect 15620 2292 15626 2304
rect 16022 2292 16028 2304
rect 15620 2264 16028 2292
rect 15620 2252 15626 2264
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17696 2292 17724 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 18616 2369 18644 2456
rect 18601 2363 18659 2369
rect 18601 2329 18613 2363
rect 18647 2329 18659 2363
rect 18601 2323 18659 2329
rect 16816 2264 17724 2292
rect 18417 2295 18475 2301
rect 16816 2252 16822 2264
rect 18417 2261 18429 2295
rect 18463 2292 18475 2295
rect 19794 2292 19800 2304
rect 18463 2264 19800 2292
rect 18463 2261 18475 2264
rect 18417 2255 18475 2261
rect 19794 2252 19800 2264
rect 19852 2252 19858 2304
rect 1104 2202 22976 2224
rect 1104 2150 6378 2202
rect 6430 2150 6442 2202
rect 6494 2150 6506 2202
rect 6558 2150 6570 2202
rect 6622 2150 6634 2202
rect 6686 2150 11806 2202
rect 11858 2150 11870 2202
rect 11922 2150 11934 2202
rect 11986 2150 11998 2202
rect 12050 2150 12062 2202
rect 12114 2150 17234 2202
rect 17286 2150 17298 2202
rect 17350 2150 17362 2202
rect 17414 2150 17426 2202
rect 17478 2150 17490 2202
rect 17542 2150 22662 2202
rect 22714 2150 22726 2202
rect 22778 2150 22790 2202
rect 22842 2150 22854 2202
rect 22906 2150 22918 2202
rect 22970 2150 22976 2202
rect 1104 2128 22976 2150
<< via1 >>
rect 6378 21734 6430 21786
rect 6442 21734 6494 21786
rect 6506 21734 6558 21786
rect 6570 21734 6622 21786
rect 6634 21734 6686 21786
rect 11806 21734 11858 21786
rect 11870 21734 11922 21786
rect 11934 21734 11986 21786
rect 11998 21734 12050 21786
rect 12062 21734 12114 21786
rect 17234 21734 17286 21786
rect 17298 21734 17350 21786
rect 17362 21734 17414 21786
rect 17426 21734 17478 21786
rect 17490 21734 17542 21786
rect 22662 21734 22714 21786
rect 22726 21734 22778 21786
rect 22790 21734 22842 21786
rect 22854 21734 22906 21786
rect 22918 21734 22970 21786
rect 3664 21190 3716 21242
rect 3728 21190 3780 21242
rect 3792 21190 3844 21242
rect 3856 21190 3908 21242
rect 3920 21190 3972 21242
rect 9092 21190 9144 21242
rect 9156 21190 9208 21242
rect 9220 21190 9272 21242
rect 9284 21190 9336 21242
rect 9348 21190 9400 21242
rect 14520 21190 14572 21242
rect 14584 21190 14636 21242
rect 14648 21190 14700 21242
rect 14712 21190 14764 21242
rect 14776 21190 14828 21242
rect 19948 21190 20000 21242
rect 20012 21190 20064 21242
rect 20076 21190 20128 21242
rect 20140 21190 20192 21242
rect 20204 21190 20256 21242
rect 6378 20646 6430 20698
rect 6442 20646 6494 20698
rect 6506 20646 6558 20698
rect 6570 20646 6622 20698
rect 6634 20646 6686 20698
rect 11806 20646 11858 20698
rect 11870 20646 11922 20698
rect 11934 20646 11986 20698
rect 11998 20646 12050 20698
rect 12062 20646 12114 20698
rect 17234 20646 17286 20698
rect 17298 20646 17350 20698
rect 17362 20646 17414 20698
rect 17426 20646 17478 20698
rect 17490 20646 17542 20698
rect 22662 20646 22714 20698
rect 22726 20646 22778 20698
rect 22790 20646 22842 20698
rect 22854 20646 22906 20698
rect 22918 20646 22970 20698
rect 3664 20102 3716 20154
rect 3728 20102 3780 20154
rect 3792 20102 3844 20154
rect 3856 20102 3908 20154
rect 3920 20102 3972 20154
rect 9092 20102 9144 20154
rect 9156 20102 9208 20154
rect 9220 20102 9272 20154
rect 9284 20102 9336 20154
rect 9348 20102 9400 20154
rect 14520 20102 14572 20154
rect 14584 20102 14636 20154
rect 14648 20102 14700 20154
rect 14712 20102 14764 20154
rect 14776 20102 14828 20154
rect 19948 20102 20000 20154
rect 20012 20102 20064 20154
rect 20076 20102 20128 20154
rect 20140 20102 20192 20154
rect 20204 20102 20256 20154
rect 6378 19558 6430 19610
rect 6442 19558 6494 19610
rect 6506 19558 6558 19610
rect 6570 19558 6622 19610
rect 6634 19558 6686 19610
rect 11806 19558 11858 19610
rect 11870 19558 11922 19610
rect 11934 19558 11986 19610
rect 11998 19558 12050 19610
rect 12062 19558 12114 19610
rect 17234 19558 17286 19610
rect 17298 19558 17350 19610
rect 17362 19558 17414 19610
rect 17426 19558 17478 19610
rect 17490 19558 17542 19610
rect 22662 19558 22714 19610
rect 22726 19558 22778 19610
rect 22790 19558 22842 19610
rect 22854 19558 22906 19610
rect 22918 19558 22970 19610
rect 2136 19499 2188 19508
rect 2136 19465 2145 19499
rect 2145 19465 2179 19499
rect 2179 19465 2188 19499
rect 2136 19456 2188 19465
rect 1860 19320 1912 19372
rect 3664 19014 3716 19066
rect 3728 19014 3780 19066
rect 3792 19014 3844 19066
rect 3856 19014 3908 19066
rect 3920 19014 3972 19066
rect 9092 19014 9144 19066
rect 9156 19014 9208 19066
rect 9220 19014 9272 19066
rect 9284 19014 9336 19066
rect 9348 19014 9400 19066
rect 14520 19014 14572 19066
rect 14584 19014 14636 19066
rect 14648 19014 14700 19066
rect 14712 19014 14764 19066
rect 14776 19014 14828 19066
rect 19948 19014 20000 19066
rect 20012 19014 20064 19066
rect 20076 19014 20128 19066
rect 20140 19014 20192 19066
rect 20204 19014 20256 19066
rect 6378 18470 6430 18522
rect 6442 18470 6494 18522
rect 6506 18470 6558 18522
rect 6570 18470 6622 18522
rect 6634 18470 6686 18522
rect 11806 18470 11858 18522
rect 11870 18470 11922 18522
rect 11934 18470 11986 18522
rect 11998 18470 12050 18522
rect 12062 18470 12114 18522
rect 17234 18470 17286 18522
rect 17298 18470 17350 18522
rect 17362 18470 17414 18522
rect 17426 18470 17478 18522
rect 17490 18470 17542 18522
rect 22662 18470 22714 18522
rect 22726 18470 22778 18522
rect 22790 18470 22842 18522
rect 22854 18470 22906 18522
rect 22918 18470 22970 18522
rect 3664 17926 3716 17978
rect 3728 17926 3780 17978
rect 3792 17926 3844 17978
rect 3856 17926 3908 17978
rect 3920 17926 3972 17978
rect 9092 17926 9144 17978
rect 9156 17926 9208 17978
rect 9220 17926 9272 17978
rect 9284 17926 9336 17978
rect 9348 17926 9400 17978
rect 14520 17926 14572 17978
rect 14584 17926 14636 17978
rect 14648 17926 14700 17978
rect 14712 17926 14764 17978
rect 14776 17926 14828 17978
rect 19948 17926 20000 17978
rect 20012 17926 20064 17978
rect 20076 17926 20128 17978
rect 20140 17926 20192 17978
rect 20204 17926 20256 17978
rect 6378 17382 6430 17434
rect 6442 17382 6494 17434
rect 6506 17382 6558 17434
rect 6570 17382 6622 17434
rect 6634 17382 6686 17434
rect 11806 17382 11858 17434
rect 11870 17382 11922 17434
rect 11934 17382 11986 17434
rect 11998 17382 12050 17434
rect 12062 17382 12114 17434
rect 17234 17382 17286 17434
rect 17298 17382 17350 17434
rect 17362 17382 17414 17434
rect 17426 17382 17478 17434
rect 17490 17382 17542 17434
rect 22662 17382 22714 17434
rect 22726 17382 22778 17434
rect 22790 17382 22842 17434
rect 22854 17382 22906 17434
rect 22918 17382 22970 17434
rect 3664 16838 3716 16890
rect 3728 16838 3780 16890
rect 3792 16838 3844 16890
rect 3856 16838 3908 16890
rect 3920 16838 3972 16890
rect 9092 16838 9144 16890
rect 9156 16838 9208 16890
rect 9220 16838 9272 16890
rect 9284 16838 9336 16890
rect 9348 16838 9400 16890
rect 14520 16838 14572 16890
rect 14584 16838 14636 16890
rect 14648 16838 14700 16890
rect 14712 16838 14764 16890
rect 14776 16838 14828 16890
rect 19948 16838 20000 16890
rect 20012 16838 20064 16890
rect 20076 16838 20128 16890
rect 20140 16838 20192 16890
rect 20204 16838 20256 16890
rect 6378 16294 6430 16346
rect 6442 16294 6494 16346
rect 6506 16294 6558 16346
rect 6570 16294 6622 16346
rect 6634 16294 6686 16346
rect 11806 16294 11858 16346
rect 11870 16294 11922 16346
rect 11934 16294 11986 16346
rect 11998 16294 12050 16346
rect 12062 16294 12114 16346
rect 17234 16294 17286 16346
rect 17298 16294 17350 16346
rect 17362 16294 17414 16346
rect 17426 16294 17478 16346
rect 17490 16294 17542 16346
rect 22662 16294 22714 16346
rect 22726 16294 22778 16346
rect 22790 16294 22842 16346
rect 22854 16294 22906 16346
rect 22918 16294 22970 16346
rect 5540 16124 5592 16176
rect 5172 16056 5224 16108
rect 5264 15988 5316 16040
rect 6092 16056 6144 16108
rect 8208 16056 8260 16108
rect 6276 15988 6328 16040
rect 4068 15852 4120 15904
rect 5540 15852 5592 15904
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 3664 15750 3716 15802
rect 3728 15750 3780 15802
rect 3792 15750 3844 15802
rect 3856 15750 3908 15802
rect 3920 15750 3972 15802
rect 9092 15750 9144 15802
rect 9156 15750 9208 15802
rect 9220 15750 9272 15802
rect 9284 15750 9336 15802
rect 9348 15750 9400 15802
rect 14520 15750 14572 15802
rect 14584 15750 14636 15802
rect 14648 15750 14700 15802
rect 14712 15750 14764 15802
rect 14776 15750 14828 15802
rect 19948 15750 20000 15802
rect 20012 15750 20064 15802
rect 20076 15750 20128 15802
rect 20140 15750 20192 15802
rect 20204 15750 20256 15802
rect 8208 15648 8260 15700
rect 6092 15580 6144 15632
rect 8116 15580 8168 15632
rect 5264 15487 5316 15496
rect 4896 15351 4948 15360
rect 4896 15317 4905 15351
rect 4905 15317 4939 15351
rect 4939 15317 4948 15351
rect 4896 15308 4948 15317
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 5540 15444 5592 15496
rect 6828 15512 6880 15564
rect 6920 15487 6972 15496
rect 5172 15419 5224 15428
rect 5172 15385 5181 15419
rect 5181 15385 5215 15419
rect 5215 15385 5224 15419
rect 6920 15453 6929 15487
rect 6929 15453 6963 15487
rect 6963 15453 6972 15487
rect 6920 15444 6972 15453
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 6092 15419 6144 15428
rect 5172 15376 5224 15385
rect 6092 15385 6101 15419
rect 6101 15385 6135 15419
rect 6135 15385 6144 15419
rect 6092 15376 6144 15385
rect 6276 15419 6328 15428
rect 6276 15385 6285 15419
rect 6285 15385 6319 15419
rect 6319 15385 6328 15419
rect 8760 15580 8812 15632
rect 7564 15419 7616 15428
rect 6276 15376 6328 15385
rect 7564 15385 7573 15419
rect 7573 15385 7607 15419
rect 7607 15385 7616 15419
rect 7564 15376 7616 15385
rect 7748 15419 7800 15428
rect 7748 15385 7757 15419
rect 7757 15385 7791 15419
rect 7791 15385 7800 15419
rect 7748 15376 7800 15385
rect 8760 15444 8812 15496
rect 9588 15376 9640 15428
rect 10600 15376 10652 15428
rect 6736 15351 6788 15360
rect 6736 15317 6745 15351
rect 6745 15317 6779 15351
rect 6779 15317 6788 15351
rect 6736 15308 6788 15317
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 9404 15351 9456 15360
rect 9404 15317 9413 15351
rect 9413 15317 9447 15351
rect 9447 15317 9456 15351
rect 9404 15308 9456 15317
rect 6378 15206 6430 15258
rect 6442 15206 6494 15258
rect 6506 15206 6558 15258
rect 6570 15206 6622 15258
rect 6634 15206 6686 15258
rect 11806 15206 11858 15258
rect 11870 15206 11922 15258
rect 11934 15206 11986 15258
rect 11998 15206 12050 15258
rect 12062 15206 12114 15258
rect 17234 15206 17286 15258
rect 17298 15206 17350 15258
rect 17362 15206 17414 15258
rect 17426 15206 17478 15258
rect 17490 15206 17542 15258
rect 22662 15206 22714 15258
rect 22726 15206 22778 15258
rect 22790 15206 22842 15258
rect 22854 15206 22906 15258
rect 22918 15206 22970 15258
rect 4896 15104 4948 15156
rect 6920 15104 6972 15156
rect 7104 15104 7156 15156
rect 8116 15104 8168 15156
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 5724 15036 5776 15088
rect 6276 15036 6328 15088
rect 2504 14968 2556 15020
rect 4252 14968 4304 15020
rect 5172 14968 5224 15020
rect 6828 14968 6880 15020
rect 9128 15036 9180 15088
rect 9864 15079 9916 15088
rect 9864 15045 9873 15079
rect 9873 15045 9907 15079
rect 9907 15045 9916 15079
rect 9864 15036 9916 15045
rect 8208 14968 8260 15020
rect 8760 15011 8812 15020
rect 8760 14977 8769 15011
rect 8769 14977 8803 15011
rect 8803 14977 8812 15011
rect 8760 14968 8812 14977
rect 9588 14968 9640 15020
rect 10048 15011 10100 15020
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 2780 14900 2832 14952
rect 3516 14943 3568 14952
rect 3516 14909 3525 14943
rect 3525 14909 3559 14943
rect 3559 14909 3568 14943
rect 3516 14900 3568 14909
rect 5080 14900 5132 14952
rect 3424 14832 3476 14884
rect 2136 14764 2188 14816
rect 2964 14764 3016 14816
rect 3240 14764 3292 14816
rect 4896 14764 4948 14816
rect 6828 14764 6880 14816
rect 7748 14900 7800 14952
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 9496 14900 9548 14952
rect 8944 14875 8996 14884
rect 8944 14841 8953 14875
rect 8953 14841 8987 14875
rect 8987 14841 8996 14875
rect 8944 14832 8996 14841
rect 7012 14764 7064 14816
rect 7564 14764 7616 14816
rect 9404 14764 9456 14816
rect 3664 14662 3716 14714
rect 3728 14662 3780 14714
rect 3792 14662 3844 14714
rect 3856 14662 3908 14714
rect 3920 14662 3972 14714
rect 9092 14662 9144 14714
rect 9156 14662 9208 14714
rect 9220 14662 9272 14714
rect 9284 14662 9336 14714
rect 9348 14662 9400 14714
rect 14520 14662 14572 14714
rect 14584 14662 14636 14714
rect 14648 14662 14700 14714
rect 14712 14662 14764 14714
rect 14776 14662 14828 14714
rect 19948 14662 20000 14714
rect 20012 14662 20064 14714
rect 20076 14662 20128 14714
rect 20140 14662 20192 14714
rect 20204 14662 20256 14714
rect 2320 14560 2372 14612
rect 7748 14560 7800 14612
rect 8760 14560 8812 14612
rect 9496 14560 9548 14612
rect 9588 14560 9640 14612
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2964 14467 3016 14476
rect 2780 14424 2832 14433
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 6736 14424 6788 14476
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 5540 14356 5592 14408
rect 7564 14424 7616 14476
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 5080 14331 5132 14340
rect 5080 14297 5089 14331
rect 5089 14297 5123 14331
rect 5123 14297 5132 14331
rect 5080 14288 5132 14297
rect 4896 14220 4948 14272
rect 7012 14288 7064 14340
rect 8300 14356 8352 14408
rect 10692 14424 10744 14476
rect 8668 14356 8720 14408
rect 8852 14356 8904 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 10048 14399 10100 14408
rect 10048 14365 10057 14399
rect 10057 14365 10091 14399
rect 10091 14365 10100 14399
rect 10048 14356 10100 14365
rect 6736 14220 6788 14272
rect 6378 14118 6430 14170
rect 6442 14118 6494 14170
rect 6506 14118 6558 14170
rect 6570 14118 6622 14170
rect 6634 14118 6686 14170
rect 11806 14118 11858 14170
rect 11870 14118 11922 14170
rect 11934 14118 11986 14170
rect 11998 14118 12050 14170
rect 12062 14118 12114 14170
rect 17234 14118 17286 14170
rect 17298 14118 17350 14170
rect 17362 14118 17414 14170
rect 17426 14118 17478 14170
rect 17490 14118 17542 14170
rect 22662 14118 22714 14170
rect 22726 14118 22778 14170
rect 22790 14118 22842 14170
rect 22854 14118 22906 14170
rect 22918 14118 22970 14170
rect 2044 14016 2096 14068
rect 3240 14059 3292 14068
rect 3240 14025 3249 14059
rect 3249 14025 3283 14059
rect 3283 14025 3292 14059
rect 3240 14016 3292 14025
rect 7012 13948 7064 14000
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 4252 13880 4304 13932
rect 4620 13880 4672 13932
rect 7104 13880 7156 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 9864 13880 9916 13932
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 6736 13812 6788 13864
rect 8852 13812 8904 13864
rect 9680 13812 9732 13864
rect 14280 13880 14332 13932
rect 7104 13744 7156 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 6736 13719 6788 13728
rect 6736 13685 6745 13719
rect 6745 13685 6779 13719
rect 6779 13685 6788 13719
rect 6736 13676 6788 13685
rect 10784 13676 10836 13728
rect 11152 13676 11204 13728
rect 3664 13574 3716 13626
rect 3728 13574 3780 13626
rect 3792 13574 3844 13626
rect 3856 13574 3908 13626
rect 3920 13574 3972 13626
rect 9092 13574 9144 13626
rect 9156 13574 9208 13626
rect 9220 13574 9272 13626
rect 9284 13574 9336 13626
rect 9348 13574 9400 13626
rect 14520 13574 14572 13626
rect 14584 13574 14636 13626
rect 14648 13574 14700 13626
rect 14712 13574 14764 13626
rect 14776 13574 14828 13626
rect 19948 13574 20000 13626
rect 20012 13574 20064 13626
rect 20076 13574 20128 13626
rect 20140 13574 20192 13626
rect 20204 13574 20256 13626
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 12256 13472 12308 13524
rect 2688 13379 2740 13388
rect 2688 13345 2697 13379
rect 2697 13345 2731 13379
rect 2731 13345 2740 13379
rect 2688 13336 2740 13345
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 3240 13268 3292 13320
rect 3608 13268 3660 13320
rect 5448 13404 5500 13456
rect 7656 13336 7708 13388
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 6828 13268 6880 13320
rect 6736 13200 6788 13252
rect 8944 13404 8996 13456
rect 8852 13336 8904 13388
rect 11060 13404 11112 13456
rect 12164 13336 12216 13388
rect 8300 13268 8352 13320
rect 8484 13268 8536 13320
rect 10784 13268 10836 13320
rect 10968 13268 11020 13320
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 11152 13200 11204 13252
rect 12348 13268 12400 13320
rect 12440 13200 12492 13252
rect 13268 13268 13320 13320
rect 14188 13268 14240 13320
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 2780 13132 2832 13184
rect 3424 13132 3476 13184
rect 3976 13132 4028 13184
rect 7472 13132 7524 13184
rect 8392 13132 8444 13184
rect 9588 13132 9640 13184
rect 10784 13132 10836 13184
rect 11520 13175 11572 13184
rect 11520 13141 11529 13175
rect 11529 13141 11563 13175
rect 11563 13141 11572 13175
rect 11520 13132 11572 13141
rect 6378 13030 6430 13082
rect 6442 13030 6494 13082
rect 6506 13030 6558 13082
rect 6570 13030 6622 13082
rect 6634 13030 6686 13082
rect 11806 13030 11858 13082
rect 11870 13030 11922 13082
rect 11934 13030 11986 13082
rect 11998 13030 12050 13082
rect 12062 13030 12114 13082
rect 17234 13030 17286 13082
rect 17298 13030 17350 13082
rect 17362 13030 17414 13082
rect 17426 13030 17478 13082
rect 17490 13030 17542 13082
rect 22662 13030 22714 13082
rect 22726 13030 22778 13082
rect 22790 13030 22842 13082
rect 22854 13030 22906 13082
rect 22918 13030 22970 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 5080 12928 5132 12980
rect 6828 12928 6880 12980
rect 7104 12928 7156 12980
rect 7748 12928 7800 12980
rect 9680 12928 9732 12980
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 2320 12724 2372 12776
rect 2688 12724 2740 12776
rect 3608 12835 3660 12844
rect 3608 12801 3617 12835
rect 3617 12801 3651 12835
rect 3651 12801 3660 12835
rect 3608 12792 3660 12801
rect 6736 12860 6788 12912
rect 2044 12656 2096 12708
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 5540 12792 5592 12844
rect 5724 12792 5776 12844
rect 4436 12724 4488 12776
rect 3976 12656 4028 12708
rect 9772 12860 9824 12912
rect 5080 12656 5132 12708
rect 6736 12656 6788 12708
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 4528 12588 4580 12640
rect 5172 12588 5224 12640
rect 6184 12588 6236 12640
rect 11060 12928 11112 12980
rect 10508 12860 10560 12912
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 10876 12792 10928 12844
rect 11060 12792 11112 12844
rect 11704 12792 11756 12844
rect 12624 12928 12676 12980
rect 12440 12903 12492 12912
rect 12440 12869 12449 12903
rect 12449 12869 12483 12903
rect 12483 12869 12492 12903
rect 12440 12860 12492 12869
rect 16948 12860 17000 12912
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12348 12835 12400 12844
rect 12164 12792 12216 12801
rect 12348 12801 12357 12835
rect 12357 12801 12391 12835
rect 12391 12801 12400 12835
rect 12348 12792 12400 12801
rect 14188 12835 14240 12844
rect 8300 12724 8352 12776
rect 11520 12724 11572 12776
rect 9864 12656 9916 12708
rect 11152 12656 11204 12708
rect 13452 12656 13504 12708
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 14280 12792 14332 12844
rect 9496 12588 9548 12640
rect 9680 12588 9732 12640
rect 14372 12588 14424 12640
rect 3664 12486 3716 12538
rect 3728 12486 3780 12538
rect 3792 12486 3844 12538
rect 3856 12486 3908 12538
rect 3920 12486 3972 12538
rect 9092 12486 9144 12538
rect 9156 12486 9208 12538
rect 9220 12486 9272 12538
rect 9284 12486 9336 12538
rect 9348 12486 9400 12538
rect 14520 12486 14572 12538
rect 14584 12486 14636 12538
rect 14648 12486 14700 12538
rect 14712 12486 14764 12538
rect 14776 12486 14828 12538
rect 19948 12486 20000 12538
rect 20012 12486 20064 12538
rect 20076 12486 20128 12538
rect 20140 12486 20192 12538
rect 20204 12486 20256 12538
rect 2964 12384 3016 12436
rect 4436 12384 4488 12436
rect 5172 12427 5224 12436
rect 5172 12393 5181 12427
rect 5181 12393 5215 12427
rect 5215 12393 5224 12427
rect 5172 12384 5224 12393
rect 5356 12384 5408 12436
rect 7748 12384 7800 12436
rect 8852 12384 8904 12436
rect 9680 12384 9732 12436
rect 10508 12427 10560 12436
rect 10508 12393 10517 12427
rect 10517 12393 10551 12427
rect 10551 12393 10560 12427
rect 10508 12384 10560 12393
rect 12348 12384 12400 12436
rect 10968 12316 11020 12368
rect 2136 12291 2188 12300
rect 2136 12257 2145 12291
rect 2145 12257 2179 12291
rect 2179 12257 2188 12291
rect 2136 12248 2188 12257
rect 4620 12248 4672 12300
rect 4896 12248 4948 12300
rect 11152 12291 11204 12300
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 16212 12316 16264 12368
rect 2964 12180 3016 12232
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 4712 12180 4764 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 2136 12112 2188 12164
rect 2688 12112 2740 12164
rect 4344 12112 4396 12164
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 5632 12180 5684 12232
rect 5908 12180 5960 12232
rect 6092 12180 6144 12232
rect 6920 12180 6972 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 7012 12112 7064 12164
rect 8300 12180 8352 12232
rect 8576 12180 8628 12232
rect 8944 12180 8996 12232
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 8024 12112 8076 12164
rect 9864 12180 9916 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 12348 12180 12400 12232
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 12440 12112 12492 12164
rect 14280 12291 14332 12300
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 14280 12257 14289 12291
rect 14289 12257 14323 12291
rect 14323 12257 14332 12291
rect 14280 12248 14332 12257
rect 14372 12248 14424 12300
rect 15016 12248 15068 12300
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 13912 12112 13964 12164
rect 5724 12044 5776 12096
rect 7748 12044 7800 12096
rect 8760 12044 8812 12096
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 11336 12087 11388 12096
rect 11336 12053 11345 12087
rect 11345 12053 11379 12087
rect 11379 12053 11388 12087
rect 11704 12087 11756 12096
rect 11336 12044 11388 12053
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 14280 12044 14332 12096
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 6378 11942 6430 11994
rect 6442 11942 6494 11994
rect 6506 11942 6558 11994
rect 6570 11942 6622 11994
rect 6634 11942 6686 11994
rect 11806 11942 11858 11994
rect 11870 11942 11922 11994
rect 11934 11942 11986 11994
rect 11998 11942 12050 11994
rect 12062 11942 12114 11994
rect 17234 11942 17286 11994
rect 17298 11942 17350 11994
rect 17362 11942 17414 11994
rect 17426 11942 17478 11994
rect 17490 11942 17542 11994
rect 22662 11942 22714 11994
rect 22726 11942 22778 11994
rect 22790 11942 22842 11994
rect 22854 11942 22906 11994
rect 22918 11942 22970 11994
rect 2136 11840 2188 11892
rect 4252 11883 4304 11892
rect 2044 11704 2096 11756
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 7656 11840 7708 11892
rect 11060 11883 11112 11892
rect 7472 11772 7524 11824
rect 8024 11772 8076 11824
rect 11060 11849 11069 11883
rect 11069 11849 11103 11883
rect 11103 11849 11112 11883
rect 11060 11840 11112 11849
rect 11244 11840 11296 11892
rect 14188 11840 14240 11892
rect 14740 11840 14792 11892
rect 10324 11772 10376 11824
rect 2780 11704 2832 11756
rect 3332 11704 3384 11756
rect 4068 11704 4120 11756
rect 8208 11704 8260 11756
rect 8392 11704 8444 11756
rect 2320 11568 2372 11620
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 3516 11500 3568 11552
rect 4344 11568 4396 11620
rect 6276 11636 6328 11688
rect 6460 11636 6512 11688
rect 7012 11568 7064 11620
rect 8944 11636 8996 11688
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 8852 11568 8904 11620
rect 4252 11500 4304 11552
rect 4804 11500 4856 11552
rect 5816 11500 5868 11552
rect 8208 11500 8260 11552
rect 11612 11704 11664 11756
rect 12164 11704 12216 11756
rect 12440 11704 12492 11756
rect 13268 11704 13320 11756
rect 12072 11636 12124 11688
rect 14372 11704 14424 11756
rect 14188 11636 14240 11688
rect 15200 11704 15252 11756
rect 11336 11568 11388 11620
rect 11152 11500 11204 11552
rect 12072 11500 12124 11552
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 13912 11500 13964 11509
rect 3664 11398 3716 11450
rect 3728 11398 3780 11450
rect 3792 11398 3844 11450
rect 3856 11398 3908 11450
rect 3920 11398 3972 11450
rect 9092 11398 9144 11450
rect 9156 11398 9208 11450
rect 9220 11398 9272 11450
rect 9284 11398 9336 11450
rect 9348 11398 9400 11450
rect 14520 11398 14572 11450
rect 14584 11398 14636 11450
rect 14648 11398 14700 11450
rect 14712 11398 14764 11450
rect 14776 11398 14828 11450
rect 19948 11398 20000 11450
rect 20012 11398 20064 11450
rect 20076 11398 20128 11450
rect 20140 11398 20192 11450
rect 20204 11398 20256 11450
rect 2872 11296 2924 11348
rect 4252 11296 4304 11348
rect 5448 11296 5500 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 11336 11339 11388 11348
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 11704 11296 11756 11348
rect 1860 11228 1912 11280
rect 2136 11160 2188 11212
rect 2596 11160 2648 11212
rect 2320 11092 2372 11144
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 4528 11135 4580 11144
rect 2136 11024 2188 11076
rect 2688 11024 2740 11076
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 6276 11092 6328 11144
rect 7748 11203 7800 11212
rect 7748 11169 7757 11203
rect 7757 11169 7791 11203
rect 7791 11169 7800 11203
rect 7748 11160 7800 11169
rect 8392 11135 8444 11144
rect 6736 11024 6788 11076
rect 7472 11024 7524 11076
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 9680 11092 9732 11144
rect 14280 11296 14332 11348
rect 15200 11160 15252 11212
rect 8852 11024 8904 11076
rect 11612 11024 11664 11076
rect 14188 11024 14240 11076
rect 4344 10999 4396 11008
rect 4344 10965 4353 10999
rect 4353 10965 4387 10999
rect 4387 10965 4396 10999
rect 4344 10956 4396 10965
rect 4436 10956 4488 11008
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 6378 10854 6430 10906
rect 6442 10854 6494 10906
rect 6506 10854 6558 10906
rect 6570 10854 6622 10906
rect 6634 10854 6686 10906
rect 11806 10854 11858 10906
rect 11870 10854 11922 10906
rect 11934 10854 11986 10906
rect 11998 10854 12050 10906
rect 12062 10854 12114 10906
rect 17234 10854 17286 10906
rect 17298 10854 17350 10906
rect 17362 10854 17414 10906
rect 17426 10854 17478 10906
rect 17490 10854 17542 10906
rect 22662 10854 22714 10906
rect 22726 10854 22778 10906
rect 22790 10854 22842 10906
rect 22854 10854 22906 10906
rect 22918 10854 22970 10906
rect 2136 10752 2188 10804
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 8392 10752 8444 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 3516 10684 3568 10736
rect 7104 10684 7156 10736
rect 8208 10684 8260 10736
rect 1860 10659 1912 10668
rect 1860 10625 1894 10659
rect 1894 10625 1912 10659
rect 1860 10616 1912 10625
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 13820 10752 13872 10804
rect 14372 10752 14424 10804
rect 14924 10684 14976 10736
rect 15016 10684 15068 10736
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 6184 10548 6236 10600
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9680 10548 9732 10600
rect 13360 10548 13412 10600
rect 15200 10659 15252 10668
rect 13452 10480 13504 10532
rect 13820 10548 13872 10600
rect 15200 10625 15209 10659
rect 15209 10625 15243 10659
rect 15243 10625 15252 10659
rect 15200 10616 15252 10625
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 14924 10412 14976 10464
rect 3664 10310 3716 10362
rect 3728 10310 3780 10362
rect 3792 10310 3844 10362
rect 3856 10310 3908 10362
rect 3920 10310 3972 10362
rect 9092 10310 9144 10362
rect 9156 10310 9208 10362
rect 9220 10310 9272 10362
rect 9284 10310 9336 10362
rect 9348 10310 9400 10362
rect 14520 10310 14572 10362
rect 14584 10310 14636 10362
rect 14648 10310 14700 10362
rect 14712 10310 14764 10362
rect 14776 10310 14828 10362
rect 19948 10310 20000 10362
rect 20012 10310 20064 10362
rect 20076 10310 20128 10362
rect 20140 10310 20192 10362
rect 20204 10310 20256 10362
rect 2688 10208 2740 10260
rect 6092 10208 6144 10260
rect 8208 10208 8260 10260
rect 12072 10208 12124 10260
rect 13820 10140 13872 10192
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 14372 10115 14424 10124
rect 14372 10081 14381 10115
rect 14381 10081 14415 10115
rect 14415 10081 14424 10115
rect 14372 10072 14424 10081
rect 1584 10004 1636 10056
rect 3424 10004 3476 10056
rect 4068 10004 4120 10056
rect 5724 10004 5776 10056
rect 7196 10004 7248 10056
rect 9680 10004 9732 10056
rect 12532 10004 12584 10056
rect 14188 10004 14240 10056
rect 14924 10072 14976 10124
rect 4436 9936 4488 9988
rect 6000 9936 6052 9988
rect 11152 9936 11204 9988
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 15660 9868 15712 9877
rect 6378 9766 6430 9818
rect 6442 9766 6494 9818
rect 6506 9766 6558 9818
rect 6570 9766 6622 9818
rect 6634 9766 6686 9818
rect 11806 9766 11858 9818
rect 11870 9766 11922 9818
rect 11934 9766 11986 9818
rect 11998 9766 12050 9818
rect 12062 9766 12114 9818
rect 17234 9766 17286 9818
rect 17298 9766 17350 9818
rect 17362 9766 17414 9818
rect 17426 9766 17478 9818
rect 17490 9766 17542 9818
rect 22662 9766 22714 9818
rect 22726 9766 22778 9818
rect 22790 9766 22842 9818
rect 22854 9766 22906 9818
rect 22918 9766 22970 9818
rect 1952 9596 2004 9648
rect 4344 9596 4396 9648
rect 9404 9639 9456 9648
rect 9404 9605 9422 9639
rect 9422 9605 9456 9639
rect 9404 9596 9456 9605
rect 13360 9639 13412 9648
rect 13360 9605 13369 9639
rect 13369 9605 13403 9639
rect 13403 9605 13412 9639
rect 13360 9596 13412 9605
rect 16580 9596 16632 9648
rect 4068 9528 4120 9580
rect 14924 9528 14976 9580
rect 15292 9528 15344 9580
rect 16212 9528 16264 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 13820 9460 13872 9512
rect 2872 9392 2924 9444
rect 5908 9392 5960 9444
rect 15016 9392 15068 9444
rect 16948 9392 17000 9444
rect 9772 9324 9824 9376
rect 12900 9324 12952 9376
rect 17040 9324 17092 9376
rect 3664 9222 3716 9274
rect 3728 9222 3780 9274
rect 3792 9222 3844 9274
rect 3856 9222 3908 9274
rect 3920 9222 3972 9274
rect 9092 9222 9144 9274
rect 9156 9222 9208 9274
rect 9220 9222 9272 9274
rect 9284 9222 9336 9274
rect 9348 9222 9400 9274
rect 14520 9222 14572 9274
rect 14584 9222 14636 9274
rect 14648 9222 14700 9274
rect 14712 9222 14764 9274
rect 14776 9222 14828 9274
rect 19948 9222 20000 9274
rect 20012 9222 20064 9274
rect 20076 9222 20128 9274
rect 20140 9222 20192 9274
rect 20204 9222 20256 9274
rect 4620 9120 4672 9172
rect 8944 9120 8996 9172
rect 14280 9120 14332 9172
rect 14372 9120 14424 9172
rect 17684 9120 17736 9172
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 9680 8984 9732 9036
rect 18604 9052 18656 9104
rect 19616 9095 19668 9104
rect 13360 8984 13412 9036
rect 4068 8916 4120 8968
rect 4252 8959 4304 8968
rect 4252 8925 4286 8959
rect 4286 8925 4304 8959
rect 4252 8916 4304 8925
rect 8392 8916 8444 8968
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 15660 8984 15712 9036
rect 19616 9061 19625 9095
rect 19625 9061 19659 9095
rect 19659 9061 19668 9095
rect 19616 9052 19668 9061
rect 13268 8848 13320 8900
rect 13820 8848 13872 8900
rect 16120 8916 16172 8968
rect 16764 8916 16816 8968
rect 16396 8848 16448 8900
rect 16488 8848 16540 8900
rect 17776 8916 17828 8968
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 19708 8916 19760 8968
rect 16948 8848 17000 8900
rect 18972 8848 19024 8900
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 16304 8780 16356 8832
rect 6378 8678 6430 8730
rect 6442 8678 6494 8730
rect 6506 8678 6558 8730
rect 6570 8678 6622 8730
rect 6634 8678 6686 8730
rect 11806 8678 11858 8730
rect 11870 8678 11922 8730
rect 11934 8678 11986 8730
rect 11998 8678 12050 8730
rect 12062 8678 12114 8730
rect 17234 8678 17286 8730
rect 17298 8678 17350 8730
rect 17362 8678 17414 8730
rect 17426 8678 17478 8730
rect 17490 8678 17542 8730
rect 22662 8678 22714 8730
rect 22726 8678 22778 8730
rect 22790 8678 22842 8730
rect 22854 8678 22906 8730
rect 22918 8678 22970 8730
rect 4712 8576 4764 8628
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 11612 8576 11664 8628
rect 2228 8508 2280 8560
rect 7196 8508 7248 8560
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 8760 8440 8812 8492
rect 18052 8619 18104 8628
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 19616 8576 19668 8628
rect 13268 8508 13320 8560
rect 9680 8440 9732 8492
rect 1584 8372 1636 8424
rect 4436 8304 4488 8356
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 14096 8483 14148 8492
rect 13912 8440 13964 8449
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 14372 8440 14424 8492
rect 15660 8508 15712 8560
rect 15476 8440 15528 8492
rect 16396 8508 16448 8560
rect 14004 8372 14056 8424
rect 15660 8372 15712 8424
rect 16212 8440 16264 8492
rect 17684 8440 17736 8492
rect 19892 8508 19944 8560
rect 20076 8576 20128 8628
rect 16672 8372 16724 8424
rect 16948 8372 17000 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 19156 8440 19208 8492
rect 19524 8440 19576 8492
rect 19800 8483 19852 8492
rect 19800 8449 19810 8483
rect 19810 8449 19844 8483
rect 19844 8449 19852 8483
rect 19800 8440 19852 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20352 8440 20404 8492
rect 15200 8304 15252 8356
rect 18420 8304 18472 8356
rect 18880 8347 18932 8356
rect 18880 8313 18889 8347
rect 18889 8313 18923 8347
rect 18923 8313 18932 8347
rect 18880 8304 18932 8313
rect 19616 8304 19668 8356
rect 20076 8304 20128 8356
rect 20444 8372 20496 8424
rect 5448 8236 5500 8288
rect 13360 8236 13412 8288
rect 17684 8236 17736 8288
rect 19064 8236 19116 8288
rect 3664 8134 3716 8186
rect 3728 8134 3780 8186
rect 3792 8134 3844 8186
rect 3856 8134 3908 8186
rect 3920 8134 3972 8186
rect 9092 8134 9144 8186
rect 9156 8134 9208 8186
rect 9220 8134 9272 8186
rect 9284 8134 9336 8186
rect 9348 8134 9400 8186
rect 14520 8134 14572 8186
rect 14584 8134 14636 8186
rect 14648 8134 14700 8186
rect 14712 8134 14764 8186
rect 14776 8134 14828 8186
rect 19948 8134 20000 8186
rect 20012 8134 20064 8186
rect 20076 8134 20128 8186
rect 20140 8134 20192 8186
rect 20204 8134 20256 8186
rect 6276 8032 6328 8084
rect 8484 8032 8536 8084
rect 12716 8032 12768 8084
rect 15200 8075 15252 8084
rect 15200 8041 15209 8075
rect 15209 8041 15243 8075
rect 15243 8041 15252 8075
rect 15200 8032 15252 8041
rect 16488 8032 16540 8084
rect 18972 8032 19024 8084
rect 19800 8032 19852 8084
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 3332 7828 3384 7880
rect 4804 7896 4856 7948
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 9680 7896 9732 7948
rect 12992 7896 13044 7948
rect 1952 7760 2004 7812
rect 4068 7692 4120 7744
rect 4620 7828 4672 7880
rect 12900 7828 12952 7880
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 15752 7896 15804 7948
rect 16304 7896 16356 7948
rect 17500 7964 17552 8016
rect 17684 7896 17736 7948
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15200 7828 15252 7880
rect 15476 7828 15528 7880
rect 16672 7828 16724 7880
rect 4896 7760 4948 7812
rect 5448 7803 5500 7812
rect 5448 7769 5482 7803
rect 5482 7769 5500 7803
rect 5448 7760 5500 7769
rect 10232 7760 10284 7812
rect 14004 7760 14056 7812
rect 15660 7760 15712 7812
rect 19340 7828 19392 7880
rect 19800 7896 19852 7948
rect 20168 7828 20220 7880
rect 20536 7828 20588 7880
rect 17776 7803 17828 7812
rect 17776 7769 17801 7803
rect 17801 7769 17828 7803
rect 17776 7760 17828 7769
rect 4528 7692 4580 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 12624 7692 12676 7744
rect 13268 7692 13320 7744
rect 13544 7692 13596 7744
rect 15016 7692 15068 7744
rect 15476 7692 15528 7744
rect 15936 7692 15988 7744
rect 17500 7692 17552 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18420 7803 18472 7812
rect 18420 7769 18429 7803
rect 18429 7769 18463 7803
rect 18463 7769 18472 7803
rect 18420 7760 18472 7769
rect 19708 7692 19760 7744
rect 6378 7590 6430 7642
rect 6442 7590 6494 7642
rect 6506 7590 6558 7642
rect 6570 7590 6622 7642
rect 6634 7590 6686 7642
rect 11806 7590 11858 7642
rect 11870 7590 11922 7642
rect 11934 7590 11986 7642
rect 11998 7590 12050 7642
rect 12062 7590 12114 7642
rect 17234 7590 17286 7642
rect 17298 7590 17350 7642
rect 17362 7590 17414 7642
rect 17426 7590 17478 7642
rect 17490 7590 17542 7642
rect 22662 7590 22714 7642
rect 22726 7590 22778 7642
rect 22790 7590 22842 7642
rect 22854 7590 22906 7642
rect 22918 7590 22970 7642
rect 1952 7531 2004 7540
rect 1952 7497 1961 7531
rect 1961 7497 1995 7531
rect 1995 7497 2004 7531
rect 1952 7488 2004 7497
rect 4068 7488 4120 7540
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 17132 7488 17184 7540
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 1584 7420 1636 7472
rect 7380 7420 7432 7472
rect 9680 7420 9732 7472
rect 16028 7420 16080 7472
rect 17960 7420 18012 7472
rect 18512 7420 18564 7472
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5264 7352 5316 7404
rect 12624 7352 12676 7404
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 5356 7284 5408 7336
rect 13544 7284 13596 7336
rect 12348 7216 12400 7268
rect 15016 7352 15068 7404
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 4896 7148 4948 7200
rect 6920 7148 6972 7200
rect 11244 7148 11296 7200
rect 13636 7148 13688 7200
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 19340 7420 19392 7472
rect 20352 7420 20404 7472
rect 18696 7352 18748 7361
rect 19064 7352 19116 7404
rect 16028 7284 16080 7336
rect 17592 7327 17644 7336
rect 16764 7216 16816 7268
rect 17592 7293 17601 7327
rect 17601 7293 17635 7327
rect 17635 7293 17644 7327
rect 17592 7284 17644 7293
rect 17776 7327 17828 7336
rect 17776 7293 17785 7327
rect 17785 7293 17819 7327
rect 17819 7293 17828 7327
rect 17776 7284 17828 7293
rect 18236 7284 18288 7336
rect 18696 7216 18748 7268
rect 20168 7259 20220 7268
rect 20168 7225 20177 7259
rect 20177 7225 20211 7259
rect 20211 7225 20220 7259
rect 20168 7216 20220 7225
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 16948 7148 17000 7200
rect 17868 7148 17920 7200
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20352 7148 20404 7157
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 9092 7046 9144 7098
rect 9156 7046 9208 7098
rect 9220 7046 9272 7098
rect 9284 7046 9336 7098
rect 9348 7046 9400 7098
rect 14520 7046 14572 7098
rect 14584 7046 14636 7098
rect 14648 7046 14700 7098
rect 14712 7046 14764 7098
rect 14776 7046 14828 7098
rect 19948 7046 20000 7098
rect 20012 7046 20064 7098
rect 20076 7046 20128 7098
rect 20140 7046 20192 7098
rect 20204 7046 20256 7098
rect 15200 6944 15252 6996
rect 15752 6919 15804 6928
rect 15752 6885 15761 6919
rect 15761 6885 15795 6919
rect 15795 6885 15804 6919
rect 15752 6876 15804 6885
rect 16120 6876 16172 6928
rect 17776 6876 17828 6928
rect 19156 6876 19208 6928
rect 5264 6808 5316 6860
rect 9680 6808 9732 6860
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 4252 6740 4304 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4528 6740 4580 6792
rect 4160 6672 4212 6724
rect 4896 6740 4948 6792
rect 5908 6715 5960 6724
rect 5908 6681 5917 6715
rect 5917 6681 5951 6715
rect 5951 6681 5960 6715
rect 5908 6672 5960 6681
rect 11244 6740 11296 6792
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 10508 6672 10560 6724
rect 12624 6672 12676 6724
rect 13544 6672 13596 6724
rect 13912 6740 13964 6792
rect 18420 6808 18472 6860
rect 18696 6808 18748 6860
rect 19800 6851 19852 6860
rect 19800 6817 19809 6851
rect 19809 6817 19843 6851
rect 19843 6817 19852 6851
rect 19800 6808 19852 6817
rect 15936 6740 15988 6792
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 17776 6740 17828 6792
rect 18880 6740 18932 6792
rect 19708 6783 19760 6792
rect 19708 6749 19717 6783
rect 19717 6749 19751 6783
rect 19751 6749 19760 6783
rect 19708 6740 19760 6749
rect 14004 6672 14056 6724
rect 15660 6672 15712 6724
rect 16120 6672 16172 6724
rect 16948 6672 17000 6724
rect 20812 6672 20864 6724
rect 2872 6604 2924 6656
rect 4804 6604 4856 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 13084 6647 13136 6656
rect 13084 6613 13099 6647
rect 13099 6613 13133 6647
rect 13133 6613 13136 6647
rect 13084 6604 13136 6613
rect 15016 6604 15068 6656
rect 19340 6604 19392 6656
rect 6378 6502 6430 6554
rect 6442 6502 6494 6554
rect 6506 6502 6558 6554
rect 6570 6502 6622 6554
rect 6634 6502 6686 6554
rect 11806 6502 11858 6554
rect 11870 6502 11922 6554
rect 11934 6502 11986 6554
rect 11998 6502 12050 6554
rect 12062 6502 12114 6554
rect 17234 6502 17286 6554
rect 17298 6502 17350 6554
rect 17362 6502 17414 6554
rect 17426 6502 17478 6554
rect 17490 6502 17542 6554
rect 22662 6502 22714 6554
rect 22726 6502 22778 6554
rect 22790 6502 22842 6554
rect 22854 6502 22906 6554
rect 22918 6502 22970 6554
rect 3332 6400 3384 6452
rect 2688 6264 2740 6316
rect 4712 6332 4764 6384
rect 5172 6400 5224 6452
rect 8116 6400 8168 6452
rect 12348 6400 12400 6452
rect 7012 6375 7064 6384
rect 7012 6341 7021 6375
rect 7021 6341 7055 6375
rect 7055 6341 7064 6375
rect 7012 6332 7064 6341
rect 4252 6264 4304 6316
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 4160 6239 4212 6248
rect 4160 6205 4169 6239
rect 4169 6205 4203 6239
rect 4203 6205 4212 6239
rect 6828 6264 6880 6316
rect 16396 6400 16448 6452
rect 17592 6400 17644 6452
rect 17684 6400 17736 6452
rect 20076 6400 20128 6452
rect 20536 6400 20588 6452
rect 14004 6307 14056 6316
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 15752 6332 15804 6384
rect 17960 6332 18012 6384
rect 18880 6375 18932 6384
rect 18880 6341 18889 6375
rect 18889 6341 18923 6375
rect 18923 6341 18932 6375
rect 18880 6332 18932 6341
rect 4160 6196 4212 6205
rect 9496 6196 9548 6248
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 13084 6196 13136 6248
rect 13176 6196 13228 6248
rect 14004 6128 14056 6180
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 15936 6307 15988 6316
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 16856 6307 16908 6316
rect 15936 6264 15988 6273
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 16948 6307 17000 6316
rect 16948 6273 16958 6307
rect 16958 6273 16992 6307
rect 16992 6273 17000 6307
rect 16948 6264 17000 6273
rect 17316 6307 17368 6316
rect 17316 6273 17330 6307
rect 17330 6273 17364 6307
rect 17364 6273 17368 6307
rect 17316 6264 17368 6273
rect 3516 6060 3568 6112
rect 12624 6060 12676 6112
rect 13452 6060 13504 6112
rect 14372 6128 14424 6180
rect 18420 6196 18472 6248
rect 18696 6196 18748 6248
rect 18972 6307 19024 6316
rect 18972 6273 18981 6307
rect 18981 6273 19015 6307
rect 19015 6273 19024 6307
rect 18972 6264 19024 6273
rect 19432 6264 19484 6316
rect 19248 6196 19300 6248
rect 20076 6307 20128 6316
rect 20076 6273 20085 6307
rect 20085 6273 20119 6307
rect 20119 6273 20128 6307
rect 20076 6264 20128 6273
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 20352 6239 20404 6248
rect 20352 6205 20361 6239
rect 20361 6205 20395 6239
rect 20395 6205 20404 6239
rect 20352 6196 20404 6205
rect 19616 6128 19668 6180
rect 19800 6128 19852 6180
rect 16396 6060 16448 6112
rect 18052 6060 18104 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 20536 6060 20588 6112
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 9092 5958 9144 6010
rect 9156 5958 9208 6010
rect 9220 5958 9272 6010
rect 9284 5958 9336 6010
rect 9348 5958 9400 6010
rect 14520 5958 14572 6010
rect 14584 5958 14636 6010
rect 14648 5958 14700 6010
rect 14712 5958 14764 6010
rect 14776 5958 14828 6010
rect 19948 5958 20000 6010
rect 20012 5958 20064 6010
rect 20076 5958 20128 6010
rect 20140 5958 20192 6010
rect 20204 5958 20256 6010
rect 2688 5899 2740 5908
rect 2688 5865 2697 5899
rect 2697 5865 2731 5899
rect 2731 5865 2740 5899
rect 2688 5856 2740 5865
rect 4528 5856 4580 5908
rect 4344 5720 4396 5772
rect 4436 5720 4488 5772
rect 5172 5720 5224 5772
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 4068 5652 4120 5704
rect 4252 5652 4304 5704
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 6000 5652 6052 5704
rect 12808 5856 12860 5908
rect 13544 5856 13596 5908
rect 14096 5856 14148 5908
rect 14372 5856 14424 5908
rect 16764 5856 16816 5908
rect 17316 5856 17368 5908
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 19616 5856 19668 5908
rect 12992 5788 13044 5840
rect 13268 5788 13320 5840
rect 15936 5788 15988 5840
rect 9496 5652 9548 5704
rect 11704 5652 11756 5704
rect 13636 5720 13688 5772
rect 12716 5652 12768 5704
rect 13176 5652 13228 5704
rect 5172 5584 5224 5636
rect 5540 5584 5592 5636
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4344 5559 4396 5568
rect 4344 5525 4353 5559
rect 4353 5525 4387 5559
rect 4387 5525 4396 5559
rect 4344 5516 4396 5525
rect 6828 5516 6880 5568
rect 9588 5516 9640 5568
rect 12808 5516 12860 5568
rect 13084 5584 13136 5636
rect 14188 5652 14240 5704
rect 14372 5720 14424 5772
rect 14924 5720 14976 5772
rect 15016 5695 15068 5704
rect 14096 5584 14148 5636
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 15752 5652 15804 5704
rect 17868 5788 17920 5840
rect 16672 5720 16724 5772
rect 16396 5695 16448 5704
rect 16396 5661 16405 5695
rect 16405 5661 16439 5695
rect 16439 5661 16448 5695
rect 16396 5652 16448 5661
rect 16764 5652 16816 5704
rect 16948 5652 17000 5704
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 17776 5652 17828 5704
rect 18144 5720 18196 5772
rect 18880 5720 18932 5772
rect 19156 5720 19208 5772
rect 20352 5788 20404 5840
rect 20536 5720 20588 5772
rect 18052 5695 18104 5704
rect 18052 5661 18061 5695
rect 18061 5661 18095 5695
rect 18095 5661 18104 5695
rect 18052 5652 18104 5661
rect 19616 5652 19668 5704
rect 18420 5584 18472 5636
rect 20444 5652 20496 5704
rect 20628 5652 20680 5704
rect 20352 5584 20404 5636
rect 13452 5516 13504 5568
rect 16856 5516 16908 5568
rect 18144 5516 18196 5568
rect 19524 5516 19576 5568
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 6378 5414 6430 5466
rect 6442 5414 6494 5466
rect 6506 5414 6558 5466
rect 6570 5414 6622 5466
rect 6634 5414 6686 5466
rect 11806 5414 11858 5466
rect 11870 5414 11922 5466
rect 11934 5414 11986 5466
rect 11998 5414 12050 5466
rect 12062 5414 12114 5466
rect 17234 5414 17286 5466
rect 17298 5414 17350 5466
rect 17362 5414 17414 5466
rect 17426 5414 17478 5466
rect 17490 5414 17542 5466
rect 22662 5414 22714 5466
rect 22726 5414 22778 5466
rect 22790 5414 22842 5466
rect 22854 5414 22906 5466
rect 22918 5414 22970 5466
rect 4436 5312 4488 5364
rect 4804 5312 4856 5364
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 8668 5312 8720 5364
rect 12716 5312 12768 5364
rect 14004 5312 14056 5364
rect 18972 5312 19024 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 3516 5176 3568 5228
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 3332 5108 3384 5160
rect 4068 5176 4120 5228
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 4528 5108 4580 5160
rect 7012 5244 7064 5296
rect 7288 5176 7340 5228
rect 11704 5176 11756 5228
rect 9496 5108 9548 5160
rect 13820 5244 13872 5296
rect 15016 5244 15068 5296
rect 16396 5244 16448 5296
rect 16764 5244 16816 5296
rect 17684 5244 17736 5296
rect 19800 5287 19852 5296
rect 19800 5253 19809 5287
rect 19809 5253 19843 5287
rect 19843 5253 19852 5287
rect 19800 5244 19852 5253
rect 20628 5244 20680 5296
rect 12992 5176 13044 5228
rect 13268 5176 13320 5228
rect 14372 5176 14424 5228
rect 15200 5176 15252 5228
rect 15844 5176 15896 5228
rect 18144 5176 18196 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 19340 5176 19392 5228
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 14280 5108 14332 5160
rect 15016 5108 15068 5160
rect 17684 5108 17736 5160
rect 18788 5108 18840 5160
rect 18604 5040 18656 5092
rect 3148 4972 3200 5024
rect 4252 4972 4304 5024
rect 5172 4972 5224 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 6920 4972 6972 5024
rect 7564 4972 7616 5024
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 17776 4972 17828 5024
rect 18788 4972 18840 5024
rect 19064 4972 19116 5024
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 9092 4870 9144 4922
rect 9156 4870 9208 4922
rect 9220 4870 9272 4922
rect 9284 4870 9336 4922
rect 9348 4870 9400 4922
rect 14520 4870 14572 4922
rect 14584 4870 14636 4922
rect 14648 4870 14700 4922
rect 14712 4870 14764 4922
rect 14776 4870 14828 4922
rect 19948 4870 20000 4922
rect 20012 4870 20064 4922
rect 20076 4870 20128 4922
rect 20140 4870 20192 4922
rect 20204 4870 20256 4922
rect 7288 4768 7340 4820
rect 7472 4768 7524 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14188 4768 14240 4820
rect 15844 4811 15896 4820
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 16028 4811 16080 4820
rect 16028 4777 16037 4811
rect 16037 4777 16071 4811
rect 16071 4777 16080 4811
rect 16028 4768 16080 4777
rect 16672 4768 16724 4820
rect 17960 4811 18012 4820
rect 17960 4777 17969 4811
rect 17969 4777 18003 4811
rect 18003 4777 18012 4811
rect 17960 4768 18012 4777
rect 18420 4768 18472 4820
rect 20444 4768 20496 4820
rect 3240 4700 3292 4752
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 11152 4632 11204 4684
rect 11704 4632 11756 4684
rect 14372 4632 14424 4684
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 6828 4564 6880 4616
rect 13820 4564 13872 4616
rect 15016 4700 15068 4752
rect 15200 4632 15252 4684
rect 14832 4564 14884 4616
rect 16396 4564 16448 4616
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 17868 4700 17920 4752
rect 18512 4632 18564 4684
rect 17684 4564 17736 4616
rect 18696 4607 18748 4616
rect 3516 4496 3568 4548
rect 6552 4496 6604 4548
rect 11060 4496 11112 4548
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 19340 4496 19392 4548
rect 5356 4428 5408 4480
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 7564 4428 7616 4480
rect 14188 4428 14240 4480
rect 18328 4428 18380 4480
rect 19524 4564 19576 4616
rect 6378 4326 6430 4378
rect 6442 4326 6494 4378
rect 6506 4326 6558 4378
rect 6570 4326 6622 4378
rect 6634 4326 6686 4378
rect 11806 4326 11858 4378
rect 11870 4326 11922 4378
rect 11934 4326 11986 4378
rect 11998 4326 12050 4378
rect 12062 4326 12114 4378
rect 17234 4326 17286 4378
rect 17298 4326 17350 4378
rect 17362 4326 17414 4378
rect 17426 4326 17478 4378
rect 17490 4326 17542 4378
rect 22662 4326 22714 4378
rect 22726 4326 22778 4378
rect 22790 4326 22842 4378
rect 22854 4326 22906 4378
rect 22918 4326 22970 4378
rect 15200 4224 15252 4276
rect 18144 4224 18196 4276
rect 6920 4156 6972 4208
rect 3056 4088 3108 4140
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 6092 4088 6144 4140
rect 7012 4088 7064 4140
rect 8024 4088 8076 4140
rect 8944 4131 8996 4140
rect 8944 4097 8962 4131
rect 8962 4097 8996 4131
rect 8944 4088 8996 4097
rect 9496 4088 9548 4140
rect 11060 4088 11112 4140
rect 12164 4088 12216 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 1584 4020 1636 4072
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 7288 3995 7340 4004
rect 7288 3961 7297 3995
rect 7297 3961 7331 3995
rect 7331 3961 7340 3995
rect 7288 3952 7340 3961
rect 13176 3952 13228 4004
rect 14832 4156 14884 4208
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 15568 4131 15620 4140
rect 14188 4088 14240 4097
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 16488 4088 16540 4140
rect 16948 4088 17000 4140
rect 17040 4088 17092 4140
rect 17776 4088 17828 4140
rect 17868 4088 17920 4140
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 15752 3952 15804 4004
rect 18420 3952 18472 4004
rect 19340 4020 19392 4072
rect 2688 3884 2740 3936
rect 3516 3884 3568 3936
rect 4068 3884 4120 3936
rect 5908 3884 5960 3936
rect 6552 3884 6604 3936
rect 7104 3884 7156 3936
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 12072 3884 12124 3936
rect 13268 3884 13320 3936
rect 13912 3884 13964 3936
rect 15108 3884 15160 3936
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 18328 3884 18380 3936
rect 20536 3884 20588 3936
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 9092 3782 9144 3834
rect 9156 3782 9208 3834
rect 9220 3782 9272 3834
rect 9284 3782 9336 3834
rect 9348 3782 9400 3834
rect 14520 3782 14572 3834
rect 14584 3782 14636 3834
rect 14648 3782 14700 3834
rect 14712 3782 14764 3834
rect 14776 3782 14828 3834
rect 19948 3782 20000 3834
rect 20012 3782 20064 3834
rect 20076 3782 20128 3834
rect 20140 3782 20192 3834
rect 20204 3782 20256 3834
rect 3148 3680 3200 3732
rect 2688 3544 2740 3596
rect 4528 3680 4580 3732
rect 5356 3680 5408 3732
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 7288 3680 7340 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 13084 3680 13136 3732
rect 14924 3680 14976 3732
rect 17040 3680 17092 3732
rect 17316 3680 17368 3732
rect 11704 3612 11756 3664
rect 6552 3587 6604 3596
rect 6552 3553 6561 3587
rect 6561 3553 6595 3587
rect 6595 3553 6604 3587
rect 6552 3544 6604 3553
rect 6920 3544 6972 3596
rect 9496 3544 9548 3596
rect 13084 3587 13136 3596
rect 13084 3553 13093 3587
rect 13093 3553 13127 3587
rect 13127 3553 13136 3587
rect 15292 3612 15344 3664
rect 15844 3655 15896 3664
rect 15844 3621 15853 3655
rect 15853 3621 15887 3655
rect 15887 3621 15896 3655
rect 15844 3612 15896 3621
rect 18328 3612 18380 3664
rect 18420 3612 18472 3664
rect 13084 3544 13136 3553
rect 3332 3476 3384 3528
rect 5172 3476 5224 3528
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 7104 3476 7156 3528
rect 4804 3408 4856 3460
rect 5540 3408 5592 3460
rect 11060 3408 11112 3460
rect 7196 3340 7248 3392
rect 8116 3340 8168 3392
rect 11152 3340 11204 3392
rect 12072 3451 12124 3460
rect 12072 3417 12081 3451
rect 12081 3417 12115 3451
rect 12115 3417 12124 3451
rect 12072 3408 12124 3417
rect 12348 3476 12400 3528
rect 12624 3340 12676 3392
rect 13728 3544 13780 3596
rect 15200 3544 15252 3596
rect 16856 3544 16908 3596
rect 13636 3476 13688 3528
rect 14372 3476 14424 3528
rect 15108 3476 15160 3528
rect 16948 3476 17000 3528
rect 15936 3408 15988 3460
rect 17868 3476 17920 3528
rect 19340 3544 19392 3596
rect 18880 3476 18932 3528
rect 19524 3612 19576 3664
rect 19708 3680 19760 3732
rect 20260 3655 20312 3664
rect 20260 3621 20269 3655
rect 20269 3621 20303 3655
rect 20303 3621 20312 3655
rect 20260 3612 20312 3621
rect 17776 3408 17828 3460
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 19984 3408 20036 3460
rect 20352 3408 20404 3460
rect 16580 3340 16632 3392
rect 16764 3383 16816 3392
rect 16764 3349 16773 3383
rect 16773 3349 16807 3383
rect 16807 3349 16816 3383
rect 16764 3340 16816 3349
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 19340 3340 19392 3392
rect 6378 3238 6430 3290
rect 6442 3238 6494 3290
rect 6506 3238 6558 3290
rect 6570 3238 6622 3290
rect 6634 3238 6686 3290
rect 11806 3238 11858 3290
rect 11870 3238 11922 3290
rect 11934 3238 11986 3290
rect 11998 3238 12050 3290
rect 12062 3238 12114 3290
rect 17234 3238 17286 3290
rect 17298 3238 17350 3290
rect 17362 3238 17414 3290
rect 17426 3238 17478 3290
rect 17490 3238 17542 3290
rect 22662 3238 22714 3290
rect 22726 3238 22778 3290
rect 22790 3238 22842 3290
rect 22854 3238 22906 3290
rect 22918 3238 22970 3290
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 6736 3136 6788 3188
rect 7196 3179 7248 3188
rect 7196 3145 7205 3179
rect 7205 3145 7239 3179
rect 7239 3145 7248 3179
rect 7196 3136 7248 3145
rect 8208 3136 8260 3188
rect 12348 3136 12400 3188
rect 2688 3111 2740 3120
rect 2688 3077 2697 3111
rect 2697 3077 2731 3111
rect 2731 3077 2740 3111
rect 2688 3068 2740 3077
rect 7380 3068 7432 3120
rect 9496 3111 9548 3120
rect 9496 3077 9505 3111
rect 9505 3077 9539 3111
rect 9539 3077 9548 3111
rect 9496 3068 9548 3077
rect 11152 3111 11204 3120
rect 11152 3077 11161 3111
rect 11161 3077 11195 3111
rect 11195 3077 11204 3111
rect 11152 3068 11204 3077
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5356 3000 5408 3052
rect 4804 2932 4856 2984
rect 7564 3000 7616 3052
rect 7196 2932 7248 2984
rect 7472 2932 7524 2984
rect 9496 2932 9548 2984
rect 12992 3000 13044 3052
rect 13636 3000 13688 3052
rect 15292 3136 15344 3188
rect 18236 3136 18288 3188
rect 18512 3136 18564 3188
rect 19708 3136 19760 3188
rect 19984 3136 20036 3188
rect 15200 3068 15252 3120
rect 7104 2864 7156 2916
rect 7840 2864 7892 2916
rect 13084 2932 13136 2984
rect 12440 2864 12492 2916
rect 7012 2796 7064 2848
rect 7472 2796 7524 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 11704 2839 11756 2848
rect 11704 2805 11713 2839
rect 11713 2805 11747 2839
rect 11747 2805 11756 2839
rect 11704 2796 11756 2805
rect 12900 2839 12952 2848
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 14280 2864 14332 2916
rect 15844 3000 15896 3052
rect 15936 3000 15988 3052
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 15292 2932 15344 2984
rect 16580 2932 16632 2984
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 19524 3000 19576 3052
rect 20260 2932 20312 2984
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 15752 2796 15804 2805
rect 16856 2839 16908 2848
rect 16856 2805 16865 2839
rect 16865 2805 16899 2839
rect 16899 2805 16908 2839
rect 16856 2796 16908 2805
rect 17224 2839 17276 2848
rect 17224 2805 17233 2839
rect 17233 2805 17267 2839
rect 17267 2805 17276 2839
rect 17224 2796 17276 2805
rect 18604 2796 18656 2848
rect 19340 2796 19392 2848
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 9092 2694 9144 2746
rect 9156 2694 9208 2746
rect 9220 2694 9272 2746
rect 9284 2694 9336 2746
rect 9348 2694 9400 2746
rect 14520 2694 14572 2746
rect 14584 2694 14636 2746
rect 14648 2694 14700 2746
rect 14712 2694 14764 2746
rect 14776 2694 14828 2746
rect 19948 2694 20000 2746
rect 20012 2694 20064 2746
rect 20076 2694 20128 2746
rect 20140 2694 20192 2746
rect 20204 2694 20256 2746
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 3332 2592 3384 2644
rect 4988 2592 5040 2644
rect 6276 2592 6328 2644
rect 7288 2592 7340 2644
rect 8024 2635 8076 2644
rect 3148 2567 3200 2576
rect 3148 2533 3157 2567
rect 3157 2533 3191 2567
rect 3191 2533 3200 2567
rect 3148 2524 3200 2533
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 8944 2592 8996 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 12164 2592 12216 2644
rect 8116 2524 8168 2576
rect 13084 2592 13136 2644
rect 15936 2635 15988 2644
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 3516 2388 3568 2440
rect 4804 2431 4856 2440
rect 4804 2397 4813 2431
rect 4813 2397 4847 2431
rect 4847 2397 4856 2431
rect 4804 2388 4856 2397
rect 5356 2456 5408 2508
rect 5172 2388 5224 2440
rect 7472 2388 7524 2440
rect 8116 2388 8168 2440
rect 10048 2456 10100 2508
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 17868 2592 17920 2644
rect 19708 2592 19760 2644
rect 7196 2320 7248 2372
rect 7932 2320 7984 2372
rect 7104 2252 7156 2304
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 12900 2388 12952 2440
rect 15476 2388 15528 2440
rect 16028 2456 16080 2508
rect 18604 2456 18656 2508
rect 16948 2388 17000 2440
rect 17224 2388 17276 2440
rect 11152 2320 11204 2372
rect 15752 2363 15804 2372
rect 15752 2329 15761 2363
rect 15761 2329 15795 2363
rect 15795 2329 15804 2363
rect 15752 2320 15804 2329
rect 15844 2320 15896 2372
rect 8208 2252 8260 2261
rect 15568 2252 15620 2304
rect 16028 2252 16080 2304
rect 16764 2252 16816 2304
rect 19800 2252 19852 2304
rect 6378 2150 6430 2202
rect 6442 2150 6494 2202
rect 6506 2150 6558 2202
rect 6570 2150 6622 2202
rect 6634 2150 6686 2202
rect 11806 2150 11858 2202
rect 11870 2150 11922 2202
rect 11934 2150 11986 2202
rect 11998 2150 12050 2202
rect 12062 2150 12114 2202
rect 17234 2150 17286 2202
rect 17298 2150 17350 2202
rect 17362 2150 17414 2202
rect 17426 2150 17478 2202
rect 17490 2150 17542 2202
rect 22662 2150 22714 2202
rect 22726 2150 22778 2202
rect 22790 2150 22842 2202
rect 22854 2150 22906 2202
rect 22918 2150 22970 2202
<< metal2 >>
rect 6378 21788 6686 21797
rect 6378 21786 6384 21788
rect 6440 21786 6464 21788
rect 6520 21786 6544 21788
rect 6600 21786 6624 21788
rect 6680 21786 6686 21788
rect 6440 21734 6442 21786
rect 6622 21734 6624 21786
rect 6378 21732 6384 21734
rect 6440 21732 6464 21734
rect 6520 21732 6544 21734
rect 6600 21732 6624 21734
rect 6680 21732 6686 21734
rect 6378 21723 6686 21732
rect 11806 21788 12114 21797
rect 11806 21786 11812 21788
rect 11868 21786 11892 21788
rect 11948 21786 11972 21788
rect 12028 21786 12052 21788
rect 12108 21786 12114 21788
rect 11868 21734 11870 21786
rect 12050 21734 12052 21786
rect 11806 21732 11812 21734
rect 11868 21732 11892 21734
rect 11948 21732 11972 21734
rect 12028 21732 12052 21734
rect 12108 21732 12114 21734
rect 11806 21723 12114 21732
rect 17234 21788 17542 21797
rect 17234 21786 17240 21788
rect 17296 21786 17320 21788
rect 17376 21786 17400 21788
rect 17456 21786 17480 21788
rect 17536 21786 17542 21788
rect 17296 21734 17298 21786
rect 17478 21734 17480 21786
rect 17234 21732 17240 21734
rect 17296 21732 17320 21734
rect 17376 21732 17400 21734
rect 17456 21732 17480 21734
rect 17536 21732 17542 21734
rect 17234 21723 17542 21732
rect 22662 21788 22970 21797
rect 22662 21786 22668 21788
rect 22724 21786 22748 21788
rect 22804 21786 22828 21788
rect 22884 21786 22908 21788
rect 22964 21786 22970 21788
rect 22724 21734 22726 21786
rect 22906 21734 22908 21786
rect 22662 21732 22668 21734
rect 22724 21732 22748 21734
rect 22804 21732 22828 21734
rect 22884 21732 22908 21734
rect 22964 21732 22970 21734
rect 22662 21723 22970 21732
rect 3664 21244 3972 21253
rect 3664 21242 3670 21244
rect 3726 21242 3750 21244
rect 3806 21242 3830 21244
rect 3886 21242 3910 21244
rect 3966 21242 3972 21244
rect 3726 21190 3728 21242
rect 3908 21190 3910 21242
rect 3664 21188 3670 21190
rect 3726 21188 3750 21190
rect 3806 21188 3830 21190
rect 3886 21188 3910 21190
rect 3966 21188 3972 21190
rect 3664 21179 3972 21188
rect 9092 21244 9400 21253
rect 9092 21242 9098 21244
rect 9154 21242 9178 21244
rect 9234 21242 9258 21244
rect 9314 21242 9338 21244
rect 9394 21242 9400 21244
rect 9154 21190 9156 21242
rect 9336 21190 9338 21242
rect 9092 21188 9098 21190
rect 9154 21188 9178 21190
rect 9234 21188 9258 21190
rect 9314 21188 9338 21190
rect 9394 21188 9400 21190
rect 9092 21179 9400 21188
rect 14520 21244 14828 21253
rect 14520 21242 14526 21244
rect 14582 21242 14606 21244
rect 14662 21242 14686 21244
rect 14742 21242 14766 21244
rect 14822 21242 14828 21244
rect 14582 21190 14584 21242
rect 14764 21190 14766 21242
rect 14520 21188 14526 21190
rect 14582 21188 14606 21190
rect 14662 21188 14686 21190
rect 14742 21188 14766 21190
rect 14822 21188 14828 21190
rect 14520 21179 14828 21188
rect 19948 21244 20256 21253
rect 19948 21242 19954 21244
rect 20010 21242 20034 21244
rect 20090 21242 20114 21244
rect 20170 21242 20194 21244
rect 20250 21242 20256 21244
rect 20010 21190 20012 21242
rect 20192 21190 20194 21242
rect 19948 21188 19954 21190
rect 20010 21188 20034 21190
rect 20090 21188 20114 21190
rect 20170 21188 20194 21190
rect 20250 21188 20256 21190
rect 19948 21179 20256 21188
rect 6378 20700 6686 20709
rect 6378 20698 6384 20700
rect 6440 20698 6464 20700
rect 6520 20698 6544 20700
rect 6600 20698 6624 20700
rect 6680 20698 6686 20700
rect 6440 20646 6442 20698
rect 6622 20646 6624 20698
rect 6378 20644 6384 20646
rect 6440 20644 6464 20646
rect 6520 20644 6544 20646
rect 6600 20644 6624 20646
rect 6680 20644 6686 20646
rect 6378 20635 6686 20644
rect 11806 20700 12114 20709
rect 11806 20698 11812 20700
rect 11868 20698 11892 20700
rect 11948 20698 11972 20700
rect 12028 20698 12052 20700
rect 12108 20698 12114 20700
rect 11868 20646 11870 20698
rect 12050 20646 12052 20698
rect 11806 20644 11812 20646
rect 11868 20644 11892 20646
rect 11948 20644 11972 20646
rect 12028 20644 12052 20646
rect 12108 20644 12114 20646
rect 11806 20635 12114 20644
rect 17234 20700 17542 20709
rect 17234 20698 17240 20700
rect 17296 20698 17320 20700
rect 17376 20698 17400 20700
rect 17456 20698 17480 20700
rect 17536 20698 17542 20700
rect 17296 20646 17298 20698
rect 17478 20646 17480 20698
rect 17234 20644 17240 20646
rect 17296 20644 17320 20646
rect 17376 20644 17400 20646
rect 17456 20644 17480 20646
rect 17536 20644 17542 20646
rect 17234 20635 17542 20644
rect 22662 20700 22970 20709
rect 22662 20698 22668 20700
rect 22724 20698 22748 20700
rect 22804 20698 22828 20700
rect 22884 20698 22908 20700
rect 22964 20698 22970 20700
rect 22724 20646 22726 20698
rect 22906 20646 22908 20698
rect 22662 20644 22668 20646
rect 22724 20644 22748 20646
rect 22804 20644 22828 20646
rect 22884 20644 22908 20646
rect 22964 20644 22970 20646
rect 22662 20635 22970 20644
rect 3664 20156 3972 20165
rect 3664 20154 3670 20156
rect 3726 20154 3750 20156
rect 3806 20154 3830 20156
rect 3886 20154 3910 20156
rect 3966 20154 3972 20156
rect 3726 20102 3728 20154
rect 3908 20102 3910 20154
rect 3664 20100 3670 20102
rect 3726 20100 3750 20102
rect 3806 20100 3830 20102
rect 3886 20100 3910 20102
rect 3966 20100 3972 20102
rect 3664 20091 3972 20100
rect 9092 20156 9400 20165
rect 9092 20154 9098 20156
rect 9154 20154 9178 20156
rect 9234 20154 9258 20156
rect 9314 20154 9338 20156
rect 9394 20154 9400 20156
rect 9154 20102 9156 20154
rect 9336 20102 9338 20154
rect 9092 20100 9098 20102
rect 9154 20100 9178 20102
rect 9234 20100 9258 20102
rect 9314 20100 9338 20102
rect 9394 20100 9400 20102
rect 9092 20091 9400 20100
rect 14520 20156 14828 20165
rect 14520 20154 14526 20156
rect 14582 20154 14606 20156
rect 14662 20154 14686 20156
rect 14742 20154 14766 20156
rect 14822 20154 14828 20156
rect 14582 20102 14584 20154
rect 14764 20102 14766 20154
rect 14520 20100 14526 20102
rect 14582 20100 14606 20102
rect 14662 20100 14686 20102
rect 14742 20100 14766 20102
rect 14822 20100 14828 20102
rect 14520 20091 14828 20100
rect 19948 20156 20256 20165
rect 19948 20154 19954 20156
rect 20010 20154 20034 20156
rect 20090 20154 20114 20156
rect 20170 20154 20194 20156
rect 20250 20154 20256 20156
rect 20010 20102 20012 20154
rect 20192 20102 20194 20154
rect 19948 20100 19954 20102
rect 20010 20100 20034 20102
rect 20090 20100 20114 20102
rect 20170 20100 20194 20102
rect 20250 20100 20256 20102
rect 19948 20091 20256 20100
rect 2134 19816 2190 19825
rect 2134 19751 2190 19760
rect 2148 19514 2176 19751
rect 6378 19612 6686 19621
rect 6378 19610 6384 19612
rect 6440 19610 6464 19612
rect 6520 19610 6544 19612
rect 6600 19610 6624 19612
rect 6680 19610 6686 19612
rect 6440 19558 6442 19610
rect 6622 19558 6624 19610
rect 6378 19556 6384 19558
rect 6440 19556 6464 19558
rect 6520 19556 6544 19558
rect 6600 19556 6624 19558
rect 6680 19556 6686 19558
rect 6378 19547 6686 19556
rect 11806 19612 12114 19621
rect 11806 19610 11812 19612
rect 11868 19610 11892 19612
rect 11948 19610 11972 19612
rect 12028 19610 12052 19612
rect 12108 19610 12114 19612
rect 11868 19558 11870 19610
rect 12050 19558 12052 19610
rect 11806 19556 11812 19558
rect 11868 19556 11892 19558
rect 11948 19556 11972 19558
rect 12028 19556 12052 19558
rect 12108 19556 12114 19558
rect 11806 19547 12114 19556
rect 17234 19612 17542 19621
rect 17234 19610 17240 19612
rect 17296 19610 17320 19612
rect 17376 19610 17400 19612
rect 17456 19610 17480 19612
rect 17536 19610 17542 19612
rect 17296 19558 17298 19610
rect 17478 19558 17480 19610
rect 17234 19556 17240 19558
rect 17296 19556 17320 19558
rect 17376 19556 17400 19558
rect 17456 19556 17480 19558
rect 17536 19556 17542 19558
rect 17234 19547 17542 19556
rect 22662 19612 22970 19621
rect 22662 19610 22668 19612
rect 22724 19610 22748 19612
rect 22804 19610 22828 19612
rect 22884 19610 22908 19612
rect 22964 19610 22970 19612
rect 22724 19558 22726 19610
rect 22906 19558 22908 19610
rect 22662 19556 22668 19558
rect 22724 19556 22748 19558
rect 22804 19556 22828 19558
rect 22884 19556 22908 19558
rect 22964 19556 22970 19558
rect 22662 19547 22970 19556
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1872 12986 1900 19314
rect 3664 19068 3972 19077
rect 3664 19066 3670 19068
rect 3726 19066 3750 19068
rect 3806 19066 3830 19068
rect 3886 19066 3910 19068
rect 3966 19066 3972 19068
rect 3726 19014 3728 19066
rect 3908 19014 3910 19066
rect 3664 19012 3670 19014
rect 3726 19012 3750 19014
rect 3806 19012 3830 19014
rect 3886 19012 3910 19014
rect 3966 19012 3972 19014
rect 3664 19003 3972 19012
rect 9092 19068 9400 19077
rect 9092 19066 9098 19068
rect 9154 19066 9178 19068
rect 9234 19066 9258 19068
rect 9314 19066 9338 19068
rect 9394 19066 9400 19068
rect 9154 19014 9156 19066
rect 9336 19014 9338 19066
rect 9092 19012 9098 19014
rect 9154 19012 9178 19014
rect 9234 19012 9258 19014
rect 9314 19012 9338 19014
rect 9394 19012 9400 19014
rect 9092 19003 9400 19012
rect 14520 19068 14828 19077
rect 14520 19066 14526 19068
rect 14582 19066 14606 19068
rect 14662 19066 14686 19068
rect 14742 19066 14766 19068
rect 14822 19066 14828 19068
rect 14582 19014 14584 19066
rect 14764 19014 14766 19066
rect 14520 19012 14526 19014
rect 14582 19012 14606 19014
rect 14662 19012 14686 19014
rect 14742 19012 14766 19014
rect 14822 19012 14828 19014
rect 14520 19003 14828 19012
rect 19948 19068 20256 19077
rect 19948 19066 19954 19068
rect 20010 19066 20034 19068
rect 20090 19066 20114 19068
rect 20170 19066 20194 19068
rect 20250 19066 20256 19068
rect 20010 19014 20012 19066
rect 20192 19014 20194 19066
rect 19948 19012 19954 19014
rect 20010 19012 20034 19014
rect 20090 19012 20114 19014
rect 20170 19012 20194 19014
rect 20250 19012 20256 19014
rect 19948 19003 20256 19012
rect 6378 18524 6686 18533
rect 6378 18522 6384 18524
rect 6440 18522 6464 18524
rect 6520 18522 6544 18524
rect 6600 18522 6624 18524
rect 6680 18522 6686 18524
rect 6440 18470 6442 18522
rect 6622 18470 6624 18522
rect 6378 18468 6384 18470
rect 6440 18468 6464 18470
rect 6520 18468 6544 18470
rect 6600 18468 6624 18470
rect 6680 18468 6686 18470
rect 6378 18459 6686 18468
rect 11806 18524 12114 18533
rect 11806 18522 11812 18524
rect 11868 18522 11892 18524
rect 11948 18522 11972 18524
rect 12028 18522 12052 18524
rect 12108 18522 12114 18524
rect 11868 18470 11870 18522
rect 12050 18470 12052 18522
rect 11806 18468 11812 18470
rect 11868 18468 11892 18470
rect 11948 18468 11972 18470
rect 12028 18468 12052 18470
rect 12108 18468 12114 18470
rect 11806 18459 12114 18468
rect 17234 18524 17542 18533
rect 17234 18522 17240 18524
rect 17296 18522 17320 18524
rect 17376 18522 17400 18524
rect 17456 18522 17480 18524
rect 17536 18522 17542 18524
rect 17296 18470 17298 18522
rect 17478 18470 17480 18522
rect 17234 18468 17240 18470
rect 17296 18468 17320 18470
rect 17376 18468 17400 18470
rect 17456 18468 17480 18470
rect 17536 18468 17542 18470
rect 17234 18459 17542 18468
rect 22662 18524 22970 18533
rect 22662 18522 22668 18524
rect 22724 18522 22748 18524
rect 22804 18522 22828 18524
rect 22884 18522 22908 18524
rect 22964 18522 22970 18524
rect 22724 18470 22726 18522
rect 22906 18470 22908 18522
rect 22662 18468 22668 18470
rect 22724 18468 22748 18470
rect 22804 18468 22828 18470
rect 22884 18468 22908 18470
rect 22964 18468 22970 18470
rect 22662 18459 22970 18468
rect 3664 17980 3972 17989
rect 3664 17978 3670 17980
rect 3726 17978 3750 17980
rect 3806 17978 3830 17980
rect 3886 17978 3910 17980
rect 3966 17978 3972 17980
rect 3726 17926 3728 17978
rect 3908 17926 3910 17978
rect 3664 17924 3670 17926
rect 3726 17924 3750 17926
rect 3806 17924 3830 17926
rect 3886 17924 3910 17926
rect 3966 17924 3972 17926
rect 3664 17915 3972 17924
rect 9092 17980 9400 17989
rect 9092 17978 9098 17980
rect 9154 17978 9178 17980
rect 9234 17978 9258 17980
rect 9314 17978 9338 17980
rect 9394 17978 9400 17980
rect 9154 17926 9156 17978
rect 9336 17926 9338 17978
rect 9092 17924 9098 17926
rect 9154 17924 9178 17926
rect 9234 17924 9258 17926
rect 9314 17924 9338 17926
rect 9394 17924 9400 17926
rect 9092 17915 9400 17924
rect 14520 17980 14828 17989
rect 14520 17978 14526 17980
rect 14582 17978 14606 17980
rect 14662 17978 14686 17980
rect 14742 17978 14766 17980
rect 14822 17978 14828 17980
rect 14582 17926 14584 17978
rect 14764 17926 14766 17978
rect 14520 17924 14526 17926
rect 14582 17924 14606 17926
rect 14662 17924 14686 17926
rect 14742 17924 14766 17926
rect 14822 17924 14828 17926
rect 14520 17915 14828 17924
rect 19948 17980 20256 17989
rect 19948 17978 19954 17980
rect 20010 17978 20034 17980
rect 20090 17978 20114 17980
rect 20170 17978 20194 17980
rect 20250 17978 20256 17980
rect 20010 17926 20012 17978
rect 20192 17926 20194 17978
rect 19948 17924 19954 17926
rect 20010 17924 20034 17926
rect 20090 17924 20114 17926
rect 20170 17924 20194 17926
rect 20250 17924 20256 17926
rect 19948 17915 20256 17924
rect 6378 17436 6686 17445
rect 6378 17434 6384 17436
rect 6440 17434 6464 17436
rect 6520 17434 6544 17436
rect 6600 17434 6624 17436
rect 6680 17434 6686 17436
rect 6440 17382 6442 17434
rect 6622 17382 6624 17434
rect 6378 17380 6384 17382
rect 6440 17380 6464 17382
rect 6520 17380 6544 17382
rect 6600 17380 6624 17382
rect 6680 17380 6686 17382
rect 6378 17371 6686 17380
rect 11806 17436 12114 17445
rect 11806 17434 11812 17436
rect 11868 17434 11892 17436
rect 11948 17434 11972 17436
rect 12028 17434 12052 17436
rect 12108 17434 12114 17436
rect 11868 17382 11870 17434
rect 12050 17382 12052 17434
rect 11806 17380 11812 17382
rect 11868 17380 11892 17382
rect 11948 17380 11972 17382
rect 12028 17380 12052 17382
rect 12108 17380 12114 17382
rect 11806 17371 12114 17380
rect 17234 17436 17542 17445
rect 17234 17434 17240 17436
rect 17296 17434 17320 17436
rect 17376 17434 17400 17436
rect 17456 17434 17480 17436
rect 17536 17434 17542 17436
rect 17296 17382 17298 17434
rect 17478 17382 17480 17434
rect 17234 17380 17240 17382
rect 17296 17380 17320 17382
rect 17376 17380 17400 17382
rect 17456 17380 17480 17382
rect 17536 17380 17542 17382
rect 17234 17371 17542 17380
rect 22662 17436 22970 17445
rect 22662 17434 22668 17436
rect 22724 17434 22748 17436
rect 22804 17434 22828 17436
rect 22884 17434 22908 17436
rect 22964 17434 22970 17436
rect 22724 17382 22726 17434
rect 22906 17382 22908 17434
rect 22662 17380 22668 17382
rect 22724 17380 22748 17382
rect 22804 17380 22828 17382
rect 22884 17380 22908 17382
rect 22964 17380 22970 17382
rect 22662 17371 22970 17380
rect 3664 16892 3972 16901
rect 3664 16890 3670 16892
rect 3726 16890 3750 16892
rect 3806 16890 3830 16892
rect 3886 16890 3910 16892
rect 3966 16890 3972 16892
rect 3726 16838 3728 16890
rect 3908 16838 3910 16890
rect 3664 16836 3670 16838
rect 3726 16836 3750 16838
rect 3806 16836 3830 16838
rect 3886 16836 3910 16838
rect 3966 16836 3972 16838
rect 3664 16827 3972 16836
rect 9092 16892 9400 16901
rect 9092 16890 9098 16892
rect 9154 16890 9178 16892
rect 9234 16890 9258 16892
rect 9314 16890 9338 16892
rect 9394 16890 9400 16892
rect 9154 16838 9156 16890
rect 9336 16838 9338 16890
rect 9092 16836 9098 16838
rect 9154 16836 9178 16838
rect 9234 16836 9258 16838
rect 9314 16836 9338 16838
rect 9394 16836 9400 16838
rect 9092 16827 9400 16836
rect 14520 16892 14828 16901
rect 14520 16890 14526 16892
rect 14582 16890 14606 16892
rect 14662 16890 14686 16892
rect 14742 16890 14766 16892
rect 14822 16890 14828 16892
rect 14582 16838 14584 16890
rect 14764 16838 14766 16890
rect 14520 16836 14526 16838
rect 14582 16836 14606 16838
rect 14662 16836 14686 16838
rect 14742 16836 14766 16838
rect 14822 16836 14828 16838
rect 14520 16827 14828 16836
rect 19948 16892 20256 16901
rect 19948 16890 19954 16892
rect 20010 16890 20034 16892
rect 20090 16890 20114 16892
rect 20170 16890 20194 16892
rect 20250 16890 20256 16892
rect 20010 16838 20012 16890
rect 20192 16838 20194 16890
rect 19948 16836 19954 16838
rect 20010 16836 20034 16838
rect 20090 16836 20114 16838
rect 20170 16836 20194 16838
rect 20250 16836 20256 16838
rect 19948 16827 20256 16836
rect 6378 16348 6686 16357
rect 6378 16346 6384 16348
rect 6440 16346 6464 16348
rect 6520 16346 6544 16348
rect 6600 16346 6624 16348
rect 6680 16346 6686 16348
rect 6440 16294 6442 16346
rect 6622 16294 6624 16346
rect 6378 16292 6384 16294
rect 6440 16292 6464 16294
rect 6520 16292 6544 16294
rect 6600 16292 6624 16294
rect 6680 16292 6686 16294
rect 6378 16283 6686 16292
rect 11806 16348 12114 16357
rect 11806 16346 11812 16348
rect 11868 16346 11892 16348
rect 11948 16346 11972 16348
rect 12028 16346 12052 16348
rect 12108 16346 12114 16348
rect 11868 16294 11870 16346
rect 12050 16294 12052 16346
rect 11806 16292 11812 16294
rect 11868 16292 11892 16294
rect 11948 16292 11972 16294
rect 12028 16292 12052 16294
rect 12108 16292 12114 16294
rect 11806 16283 12114 16292
rect 17234 16348 17542 16357
rect 17234 16346 17240 16348
rect 17296 16346 17320 16348
rect 17376 16346 17400 16348
rect 17456 16346 17480 16348
rect 17536 16346 17542 16348
rect 17296 16294 17298 16346
rect 17478 16294 17480 16346
rect 17234 16292 17240 16294
rect 17296 16292 17320 16294
rect 17376 16292 17400 16294
rect 17456 16292 17480 16294
rect 17536 16292 17542 16294
rect 17234 16283 17542 16292
rect 22662 16348 22970 16357
rect 22662 16346 22668 16348
rect 22724 16346 22748 16348
rect 22804 16346 22828 16348
rect 22884 16346 22908 16348
rect 22964 16346 22970 16348
rect 22724 16294 22726 16346
rect 22906 16294 22908 16346
rect 22662 16292 22668 16294
rect 22724 16292 22748 16294
rect 22804 16292 22828 16294
rect 22884 16292 22908 16294
rect 22964 16292 22970 16294
rect 22662 16283 22970 16292
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3664 15804 3972 15813
rect 3664 15802 3670 15804
rect 3726 15802 3750 15804
rect 3806 15802 3830 15804
rect 3886 15802 3910 15804
rect 3966 15802 3972 15804
rect 3726 15750 3728 15802
rect 3908 15750 3910 15802
rect 3664 15748 3670 15750
rect 3726 15748 3750 15750
rect 3806 15748 3830 15750
rect 3886 15748 3910 15750
rect 3966 15748 3972 15750
rect 3664 15739 3972 15748
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 14074 2084 14350
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2148 13938 2176 14758
rect 2332 14618 2360 14894
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1872 10674 1900 11222
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 10062 1624 10542
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9518 1624 9998
rect 1964 9654 1992 13670
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 2056 11762 2084 12650
rect 2148 12306 2176 13126
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2148 11898 2176 12106
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 11098 2084 11698
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11218 2176 11494
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2056 11082 2176 11098
rect 2056 11076 2188 11082
rect 2056 11070 2136 11076
rect 2136 11018 2188 11024
rect 2148 10810 2176 11018
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 8430 1624 9454
rect 2240 8566 2268 14214
rect 2516 13326 2544 14962
rect 2780 14952 2832 14958
rect 3516 14952 3568 14958
rect 2780 14894 2832 14900
rect 3514 14920 3516 14929
rect 3568 14920 3570 14929
rect 2792 14482 2820 14894
rect 3424 14884 3476 14890
rect 3514 14855 3570 14864
rect 3424 14826 3476 14832
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 2976 14482 3004 14758
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 3252 14074 3280 14758
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3436 13870 3464 14826
rect 3664 14716 3972 14725
rect 3664 14714 3670 14716
rect 3726 14714 3750 14716
rect 3806 14714 3830 14716
rect 3886 14714 3910 14716
rect 3966 14714 3972 14716
rect 3726 14662 3728 14714
rect 3908 14662 3910 14714
rect 3664 14660 3670 14662
rect 3726 14660 3750 14662
rect 3806 14660 3830 14662
rect 3886 14660 3910 14662
rect 3966 14660 3972 14662
rect 3664 14651 3972 14660
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2700 12782 2728 13330
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2332 11626 2360 12718
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2332 11150 2360 11562
rect 2608 11218 2636 12038
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2700 11082 2728 12106
rect 2792 11937 2820 13126
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2778 11928 2834 11937
rect 2778 11863 2834 11872
rect 2792 11762 2820 11863
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2884 11354 2912 12786
rect 2976 12442 3004 12786
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3252 12238 3280 13262
rect 3436 13190 3464 13806
rect 3664 13628 3972 13637
rect 3664 13626 3670 13628
rect 3726 13626 3750 13628
rect 3806 13626 3830 13628
rect 3886 13626 3910 13628
rect 3966 13626 3972 13628
rect 3726 13574 3728 13626
rect 3908 13574 3910 13626
rect 3664 13572 3670 13574
rect 3726 13572 3750 13574
rect 3806 13572 3830 13574
rect 3886 13572 3910 13574
rect 3966 13572 3972 13574
rect 3664 13563 3972 13572
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3620 12850 3648 13262
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3988 12730 4016 13126
rect 4080 12850 4108 15846
rect 5184 15434 5212 16050
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5276 15502 5304 15982
rect 5552 15910 5580 16118
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15502 5580 15846
rect 6104 15638 6132 16050
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4908 15162 4936 15302
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 5184 15026 5212 15370
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3988 12714 4108 12730
rect 3976 12708 4108 12714
rect 4028 12702 4108 12708
rect 3976 12650 4028 12656
rect 3664 12540 3972 12549
rect 3664 12538 3670 12540
rect 3726 12538 3750 12540
rect 3806 12538 3830 12540
rect 3886 12538 3910 12540
rect 3966 12538 3972 12540
rect 3726 12486 3728 12538
rect 3908 12486 3910 12538
rect 3664 12484 3670 12486
rect 3726 12484 3750 12486
rect 3806 12484 3830 12486
rect 3886 12484 3910 12486
rect 3966 12484 3972 12486
rect 3664 12475 3972 12484
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2872 11144 2924 11150
rect 2976 11132 3004 12174
rect 4080 11762 4108 12702
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 2924 11104 3004 11132
rect 2872 11086 2924 11092
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2700 10266 2728 11018
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2884 9450 2912 11086
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 7954 1624 8366
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1596 7478 1624 7890
rect 3344 7886 3372 11698
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 10742 3556 11494
rect 3664 11452 3972 11461
rect 3664 11450 3670 11452
rect 3726 11450 3750 11452
rect 3806 11450 3830 11452
rect 3886 11450 3910 11452
rect 3966 11450 3972 11452
rect 3726 11398 3728 11450
rect 3908 11398 3910 11450
rect 3664 11396 3670 11398
rect 3726 11396 3750 11398
rect 3806 11396 3830 11398
rect 3886 11396 3910 11398
rect 3966 11396 3972 11398
rect 3664 11387 3972 11396
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 4172 10690 4200 14214
rect 4264 13938 4292 14962
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14414 4936 14758
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 5092 14346 5120 14894
rect 5552 14414 5580 15438
rect 6104 15434 6132 15574
rect 6288 15434 6316 15982
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6288 15094 6316 15370
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6378 15260 6686 15269
rect 6378 15258 6384 15260
rect 6440 15258 6464 15260
rect 6520 15258 6544 15260
rect 6600 15258 6624 15260
rect 6680 15258 6686 15260
rect 6440 15206 6442 15258
rect 6622 15206 6624 15258
rect 6378 15204 6384 15206
rect 6440 15204 6464 15206
rect 6520 15204 6544 15206
rect 6600 15204 6624 15206
rect 6680 15204 6686 15206
rect 6378 15195 6686 15204
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 11898 4292 12582
rect 4448 12442 4476 12718
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4356 11626 4384 12106
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11354 4292 11494
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4540 11150 4568 12582
rect 4632 12434 4660 13874
rect 4632 12406 4752 12434
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4172 10662 4292 10690
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3436 10062 3464 10542
rect 3664 10364 3972 10373
rect 3664 10362 3670 10364
rect 3726 10362 3750 10364
rect 3806 10362 3830 10364
rect 3886 10362 3910 10364
rect 3966 10362 3972 10364
rect 3726 10310 3728 10362
rect 3908 10310 3910 10362
rect 3664 10308 3670 10310
rect 3726 10308 3750 10310
rect 3806 10308 3830 10310
rect 3886 10308 3910 10310
rect 3966 10308 3972 10310
rect 3664 10299 3972 10308
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9586 4108 9998
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3664 9276 3972 9285
rect 3664 9274 3670 9276
rect 3726 9274 3750 9276
rect 3806 9274 3830 9276
rect 3886 9274 3910 9276
rect 3966 9274 3972 9276
rect 3726 9222 3728 9274
rect 3908 9222 3910 9274
rect 3664 9220 3670 9222
rect 3726 9220 3750 9222
rect 3806 9220 3830 9222
rect 3886 9220 3910 9222
rect 3966 9220 3972 9222
rect 3664 9211 3972 9220
rect 4080 8974 4108 9522
rect 4264 8974 4292 10662
rect 4356 9654 4384 10950
rect 4448 9994 4476 10950
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4632 9178 4660 12242
rect 4724 12238 4752 12406
rect 4908 12306 4936 14214
rect 5092 13818 5120 14282
rect 5092 13790 5212 13818
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5092 12714 5120 12922
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 5184 12646 5212 13790
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12442 5212 12582
rect 5368 12442 5396 14350
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 5368 12238 5396 12378
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4724 8634 4752 12174
rect 4804 11552 4856 11558
rect 5460 11506 5488 13398
rect 5736 12850 5764 15030
rect 6748 14482 6776 15302
rect 6840 15026 6868 15506
rect 7024 15502 7052 15846
rect 8220 15706 8248 16050
rect 9092 15804 9400 15813
rect 9092 15802 9098 15804
rect 9154 15802 9178 15804
rect 9234 15802 9258 15804
rect 9314 15802 9338 15804
rect 9394 15802 9400 15804
rect 9154 15750 9156 15802
rect 9336 15750 9338 15802
rect 9092 15748 9098 15750
rect 9154 15748 9178 15750
rect 9234 15748 9258 15750
rect 9314 15748 9338 15750
rect 9394 15748 9400 15750
rect 9092 15739 9400 15748
rect 14520 15804 14828 15813
rect 14520 15802 14526 15804
rect 14582 15802 14606 15804
rect 14662 15802 14686 15804
rect 14742 15802 14766 15804
rect 14822 15802 14828 15804
rect 14582 15750 14584 15802
rect 14764 15750 14766 15802
rect 14520 15748 14526 15750
rect 14582 15748 14606 15750
rect 14662 15748 14686 15750
rect 14742 15748 14766 15750
rect 14822 15748 14828 15750
rect 14520 15739 14828 15748
rect 19948 15804 20256 15813
rect 19948 15802 19954 15804
rect 20010 15802 20034 15804
rect 20090 15802 20114 15804
rect 20170 15802 20194 15804
rect 20250 15802 20256 15804
rect 20010 15750 20012 15802
rect 20192 15750 20194 15802
rect 19948 15748 19954 15750
rect 20010 15748 20034 15750
rect 20090 15748 20114 15750
rect 20170 15748 20194 15750
rect 20250 15748 20256 15750
rect 19948 15739 20256 15748
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6932 15162 6960 15438
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6828 15020 6880 15026
rect 6880 14980 6960 15008
rect 6828 14962 6880 14968
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6378 14172 6686 14181
rect 6378 14170 6384 14172
rect 6440 14170 6464 14172
rect 6520 14170 6544 14172
rect 6600 14170 6624 14172
rect 6680 14170 6686 14172
rect 6440 14118 6442 14170
rect 6622 14118 6624 14170
rect 6378 14116 6384 14118
rect 6440 14116 6464 14118
rect 6520 14116 6544 14118
rect 6600 14116 6624 14118
rect 6680 14116 6686 14118
rect 6378 14107 6686 14116
rect 6748 13870 6776 14214
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5552 12434 5580 12786
rect 6196 12646 6224 13262
rect 6748 13258 6776 13670
rect 6840 13326 6868 14758
rect 6932 14328 6960 14980
rect 7024 14822 7052 15438
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7116 14414 7144 15098
rect 7576 14822 7604 15370
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7576 14482 7604 14758
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 14340 7064 14346
rect 6932 14300 7012 14328
rect 7012 14282 7064 14288
rect 7024 14006 7052 14282
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7116 13938 7144 14350
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6378 13084 6686 13093
rect 6378 13082 6384 13084
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6680 13082 6686 13084
rect 6440 13030 6442 13082
rect 6622 13030 6624 13082
rect 6378 13028 6384 13030
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6680 13028 6686 13030
rect 6378 13019 6686 13028
rect 6748 12918 6776 13194
rect 7116 12986 7144 13738
rect 7668 13394 7696 15302
rect 7760 14958 7788 15370
rect 8128 15162 8156 15574
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8128 14958 8156 15098
rect 8220 15026 8248 15642
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8772 15502 8800 15574
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8772 15026 8800 15438
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9140 15094 9168 15302
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7760 14618 7788 14894
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 6828 12980 6880 12986
rect 7104 12980 7156 12986
rect 6880 12940 6960 12968
rect 6828 12922 6880 12928
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 5552 12406 5672 12434
rect 5644 12238 5672 12406
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 4804 11494 4856 11500
rect 4816 10810 4844 11494
rect 5368 11478 5488 11506
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3664 8188 3972 8197
rect 3664 8186 3670 8188
rect 3726 8186 3750 8188
rect 3806 8186 3830 8188
rect 3886 8186 3910 8188
rect 3966 8186 3972 8188
rect 3726 8134 3728 8186
rect 3908 8134 3910 8186
rect 3664 8132 3670 8134
rect 3726 8132 3750 8134
rect 3806 8132 3830 8134
rect 3886 8132 3910 8134
rect 3966 8132 3972 8134
rect 3664 8123 3972 8132
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7546 1992 7754
rect 4080 7750 4108 8434
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7546 4108 7686
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 3664 7100 3972 7109
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7035 3972 7044
rect 4448 6798 4476 8298
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4540 6798 4568 7686
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5166 1624 6190
rect 2700 5914 2728 6258
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2884 5710 2912 6598
rect 3344 6458 3372 6734
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3344 5710 3372 6394
rect 4172 6254 4200 6666
rect 4264 6322 4292 6734
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3528 5234 3556 6054
rect 3664 6012 3972 6021
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5947 3972 5956
rect 4264 5710 4292 6258
rect 4540 5914 4568 6734
rect 4632 6322 4660 7822
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 6390 4752 7686
rect 4816 6662 4844 7890
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4908 7206 4936 7754
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 6798 4936 7142
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4080 5234 4108 5646
rect 4356 5574 4384 5714
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4264 5250 4292 5510
rect 4448 5370 4476 5714
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4264 5234 4476 5250
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4264 5228 4488 5234
rect 4264 5222 4436 5228
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 1596 4078 1624 5102
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3602 2728 3878
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2700 3126 2728 3538
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 3068 2650 3096 4082
rect 3160 3738 3188 4966
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3160 2582 3188 3674
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3252 2446 3280 4694
rect 3344 3534 3372 5102
rect 4264 5030 4292 5222
rect 4436 5170 4488 5176
rect 4540 5166 4568 5646
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3664 4924 3972 4933
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4859 3972 4868
rect 4264 4622 4292 4966
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3528 3942 3556 4490
rect 4632 4146 4660 6258
rect 4816 5370 4844 6598
rect 5184 6458 5212 7346
rect 5276 6866 5304 7346
rect 5368 7342 5396 11478
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5460 8294 5488 11290
rect 5736 10062 5764 12038
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11150 5856 11494
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5920 9450 5948 12174
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6012 9994 6040 10950
rect 6104 10266 6132 12174
rect 6378 11996 6686 12005
rect 6378 11994 6384 11996
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6680 11994 6686 11996
rect 6440 11942 6442 11994
rect 6622 11942 6624 11994
rect 6378 11940 6384 11942
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6680 11940 6686 11942
rect 6378 11931 6686 11940
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6288 11150 6316 11630
rect 6472 11354 6500 11630
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6196 10130 6224 10542
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 7818 5488 8230
rect 6288 8090 6316 11086
rect 6748 11082 6776 12650
rect 6932 12238 6960 12940
rect 7104 12922 7156 12928
rect 7484 12238 7512 13126
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7760 12442 7788 12922
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7024 11626 7052 12106
rect 7668 11898 7696 12174
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6378 10908 6686 10917
rect 6378 10906 6384 10908
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6680 10906 6686 10908
rect 6440 10854 6442 10906
rect 6622 10854 6624 10906
rect 6378 10852 6384 10854
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6680 10852 6686 10854
rect 6378 10843 6686 10852
rect 6378 9820 6686 9829
rect 6378 9818 6384 9820
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6680 9818 6686 9820
rect 6440 9766 6442 9818
rect 6622 9766 6624 9818
rect 6378 9764 6384 9766
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6680 9764 6686 9766
rect 6378 9755 6686 9764
rect 6378 8732 6686 8741
rect 6378 8730 6384 8732
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6680 8730 6686 8732
rect 6440 8678 6442 8730
rect 6622 8678 6624 8730
rect 6378 8676 6384 8678
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6680 8676 6686 8678
rect 6378 8667 6686 8676
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5460 6882 5488 7754
rect 6378 7644 6686 7653
rect 6378 7642 6384 7644
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6680 7642 6686 7644
rect 6440 7590 6442 7642
rect 6622 7590 6624 7642
rect 6378 7588 6384 7590
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6680 7588 6686 7590
rect 6378 7579 6686 7588
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 5264 6860 5316 6866
rect 5460 6854 5580 6882
rect 5264 6802 5316 6808
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5184 5778 5212 6394
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5552 5642 5580 6854
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5184 5370 5212 5578
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 4080 3942 4108 3975
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3344 2650 3372 3470
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3528 2446 3556 3878
rect 3664 3836 3972 3845
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 3664 3771 3972 3780
rect 4528 3732 4580 3738
rect 4632 3720 4660 4082
rect 4580 3692 4660 3720
rect 4528 3674 4580 3680
rect 5184 3534 5212 4966
rect 5552 4486 5580 5578
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5368 3738 5396 4422
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4816 3194 4844 3402
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5184 3058 5212 3470
rect 5368 3058 5396 3674
rect 5552 3466 5580 4422
rect 5920 3942 5948 6666
rect 6378 6556 6686 6565
rect 6378 6554 6384 6556
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6680 6554 6686 6556
rect 6440 6502 6442 6554
rect 6622 6502 6624 6554
rect 6378 6500 6384 6502
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6680 6500 6686 6502
rect 6378 6491 6686 6500
rect 6828 6316 6880 6322
rect 6932 6304 6960 7142
rect 7024 6390 7052 11562
rect 7484 11082 7512 11766
rect 7760 11218 7788 12038
rect 8036 11830 8064 12106
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10742 7144 10950
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9042 7236 9998
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7208 8566 7236 8978
rect 7484 8634 7512 11018
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7208 7954 7236 8502
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7392 6662 7420 7414
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6880 6276 6960 6304
rect 6828 6258 6880 6264
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 4690 6040 5646
rect 6828 5568 6880 5574
rect 6932 5556 6960 6276
rect 6880 5528 6960 5556
rect 6828 5510 6880 5516
rect 6378 5468 6686 5477
rect 6378 5466 6384 5468
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6680 5466 6686 5468
rect 6440 5414 6442 5466
rect 6622 5414 6624 5466
rect 6378 5412 6384 5414
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6680 5412 6686 5414
rect 6378 5403 6686 5412
rect 6932 5030 6960 5528
rect 7024 5302 7052 6326
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6564 4554 6592 4966
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6378 4380 6686 4389
rect 6378 4378 6384 4380
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6680 4378 6686 4380
rect 6440 4326 6442 4378
rect 6622 4326 6624 4378
rect 6378 4324 6384 4326
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6680 4324 6686 4326
rect 6378 4315 6686 4324
rect 6840 4162 6868 4558
rect 6932 4214 6960 4245
rect 6920 4208 6972 4214
rect 6840 4156 6920 4162
rect 6840 4150 6972 4156
rect 6092 4140 6144 4146
rect 6840 4134 6960 4150
rect 7024 4146 7052 5238
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 4826 7328 5170
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 6092 4082 6144 4088
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 6104 3738 6132 4082
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6564 3602 6592 3878
rect 6932 3602 6960 4134
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6552 3596 6604 3602
rect 6920 3596 6972 3602
rect 6604 3556 6776 3584
rect 6552 3538 6604 3544
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 3664 2748 3972 2757
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2683 3972 2692
rect 4816 2446 4844 2926
rect 5000 2650 5028 2994
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5184 2446 5212 2994
rect 5368 2514 5396 2994
rect 6288 2650 6316 3470
rect 6378 3292 6686 3301
rect 6378 3290 6384 3292
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6680 3290 6686 3292
rect 6440 3238 6442 3290
rect 6622 3238 6624 3290
rect 6378 3236 6384 3238
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6680 3236 6686 3238
rect 6378 3227 6686 3236
rect 6748 3194 6776 3556
rect 6920 3538 6972 3544
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 7024 2854 7052 4082
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 3534 7144 3878
rect 7300 3738 7328 3946
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 3194 7236 3334
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 7116 2310 7144 2858
rect 7208 2378 7236 2926
rect 7300 2650 7328 3674
rect 7392 3126 7420 6598
rect 8128 6458 8156 14894
rect 8772 14618 8800 14962
rect 8942 14920 8998 14929
rect 8942 14855 8944 14864
rect 8996 14855 8998 14864
rect 8944 14826 8996 14832
rect 9416 14822 9444 15302
rect 9600 15026 9628 15370
rect 10612 15162 10640 15370
rect 11806 15260 12114 15269
rect 11806 15258 11812 15260
rect 11868 15258 11892 15260
rect 11948 15258 11972 15260
rect 12028 15258 12052 15260
rect 12108 15258 12114 15260
rect 11868 15206 11870 15258
rect 12050 15206 12052 15258
rect 11806 15204 11812 15206
rect 11868 15204 11892 15206
rect 11948 15204 11972 15206
rect 12028 15204 12052 15206
rect 12108 15204 12114 15206
rect 11806 15195 12114 15204
rect 17234 15260 17542 15269
rect 17234 15258 17240 15260
rect 17296 15258 17320 15260
rect 17376 15258 17400 15260
rect 17456 15258 17480 15260
rect 17536 15258 17542 15260
rect 17296 15206 17298 15258
rect 17478 15206 17480 15258
rect 17234 15204 17240 15206
rect 17296 15204 17320 15206
rect 17376 15204 17400 15206
rect 17456 15204 17480 15206
rect 17536 15204 17542 15206
rect 17234 15195 17542 15204
rect 22662 15260 22970 15269
rect 22662 15258 22668 15260
rect 22724 15258 22748 15260
rect 22804 15258 22828 15260
rect 22884 15258 22908 15260
rect 22964 15258 22970 15260
rect 22724 15206 22726 15258
rect 22906 15206 22908 15258
rect 22662 15204 22668 15206
rect 22724 15204 22748 15206
rect 22804 15204 22828 15206
rect 22884 15204 22908 15206
rect 22964 15204 22970 15206
rect 22662 15195 22970 15204
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9092 14716 9400 14725
rect 9092 14714 9098 14716
rect 9154 14714 9178 14716
rect 9234 14714 9258 14716
rect 9314 14714 9338 14716
rect 9394 14714 9400 14716
rect 9154 14662 9156 14714
rect 9336 14662 9338 14714
rect 9092 14660 9098 14662
rect 9154 14660 9178 14662
rect 9234 14660 9258 14662
rect 9314 14660 9338 14662
rect 9394 14660 9400 14662
rect 9092 14651 9400 14660
rect 9508 14618 9536 14894
rect 9600 14618 9628 14962
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9876 14414 9904 15030
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10060 14414 10088 14962
rect 10704 14482 10732 14962
rect 14520 14716 14828 14725
rect 14520 14714 14526 14716
rect 14582 14714 14606 14716
rect 14662 14714 14686 14716
rect 14742 14714 14766 14716
rect 14822 14714 14828 14716
rect 14582 14662 14584 14714
rect 14764 14662 14766 14714
rect 14520 14660 14526 14662
rect 14582 14660 14606 14662
rect 14662 14660 14686 14662
rect 14742 14660 14766 14662
rect 14822 14660 14828 14662
rect 14520 14651 14828 14660
rect 19948 14716 20256 14725
rect 19948 14714 19954 14716
rect 20010 14714 20034 14716
rect 20090 14714 20114 14716
rect 20170 14714 20194 14716
rect 20250 14714 20256 14716
rect 20010 14662 20012 14714
rect 20192 14662 20194 14714
rect 19948 14660 19954 14662
rect 20010 14660 20034 14662
rect 20090 14660 20114 14662
rect 20170 14660 20194 14662
rect 20250 14660 20256 14662
rect 19948 14651 20256 14660
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 8312 13326 8340 14350
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8404 13190 8432 13874
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12238 8340 12718
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8220 11558 8248 11698
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 10742 8248 11494
rect 8404 11150 8432 11698
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8404 10810 8432 11086
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8220 10266 8248 10678
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8404 8974 8432 10406
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8496 8090 8524 13262
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 10674 8616 12174
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8680 5370 8708 14350
rect 8864 13870 8892 14350
rect 9876 13938 9904 14350
rect 11806 14172 12114 14181
rect 11806 14170 11812 14172
rect 11868 14170 11892 14172
rect 11948 14170 11972 14172
rect 12028 14170 12052 14172
rect 12108 14170 12114 14172
rect 11868 14118 11870 14170
rect 12050 14118 12052 14170
rect 11806 14116 11812 14118
rect 11868 14116 11892 14118
rect 11948 14116 11972 14118
rect 12028 14116 12052 14118
rect 12108 14116 12114 14118
rect 11806 14107 12114 14116
rect 17234 14172 17542 14181
rect 17234 14170 17240 14172
rect 17296 14170 17320 14172
rect 17376 14170 17400 14172
rect 17456 14170 17480 14172
rect 17536 14170 17542 14172
rect 17296 14118 17298 14170
rect 17478 14118 17480 14170
rect 17234 14116 17240 14118
rect 17296 14116 17320 14118
rect 17376 14116 17400 14118
rect 17456 14116 17480 14118
rect 17536 14116 17542 14118
rect 17234 14107 17542 14116
rect 22662 14172 22970 14181
rect 22662 14170 22668 14172
rect 22724 14170 22748 14172
rect 22804 14170 22828 14172
rect 22884 14170 22908 14172
rect 22964 14170 22970 14172
rect 22724 14118 22726 14170
rect 22906 14118 22908 14170
rect 22662 14116 22668 14118
rect 22724 14116 22748 14118
rect 22804 14116 22828 14118
rect 22884 14116 22908 14118
rect 22964 14116 22970 14118
rect 22662 14107 22970 14116
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 8864 13394 8892 13806
rect 9092 13628 9400 13637
rect 9092 13626 9098 13628
rect 9154 13626 9178 13628
rect 9234 13626 9258 13628
rect 9314 13626 9338 13628
rect 9394 13626 9400 13628
rect 9154 13574 9156 13626
rect 9336 13574 9338 13626
rect 9092 13572 9098 13574
rect 9154 13572 9178 13574
rect 9234 13572 9258 13574
rect 9314 13572 9338 13574
rect 9394 13572 9400 13574
rect 9092 13563 9400 13572
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 8498 8800 12038
rect 8864 11626 8892 12378
rect 8956 12238 8984 13398
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9092 12540 9400 12549
rect 9092 12538 9098 12540
rect 9154 12538 9178 12540
rect 9234 12538 9258 12540
rect 9314 12538 9338 12540
rect 9394 12538 9400 12540
rect 9154 12486 9156 12538
rect 9336 12486 9338 12538
rect 9092 12484 9098 12486
rect 9154 12484 9178 12486
rect 9234 12484 9258 12486
rect 9314 12484 9338 12486
rect 9394 12484 9400 12486
rect 9092 12475 9400 12484
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11694 9444 12174
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11082 8892 11562
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8864 10606 8892 11018
rect 8956 10674 8984 11630
rect 9092 11452 9400 11461
rect 9092 11450 9098 11452
rect 9154 11450 9178 11452
rect 9234 11450 9258 11452
rect 9314 11450 9338 11452
rect 9394 11450 9400 11452
rect 9154 11398 9156 11450
rect 9336 11398 9338 11450
rect 9092 11396 9098 11398
rect 9154 11396 9178 11398
rect 9234 11396 9258 11398
rect 9314 11396 9338 11398
rect 9394 11396 9400 11398
rect 9092 11387 9400 11396
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8956 9178 8984 10610
rect 9092 10364 9400 10373
rect 9092 10362 9098 10364
rect 9154 10362 9178 10364
rect 9234 10362 9258 10364
rect 9314 10362 9338 10364
rect 9394 10362 9400 10364
rect 9154 10310 9156 10362
rect 9336 10310 9338 10362
rect 9092 10308 9098 10310
rect 9154 10308 9178 10310
rect 9234 10308 9258 10310
rect 9314 10308 9338 10310
rect 9394 10308 9400 10310
rect 9092 10299 9400 10308
rect 9508 10248 9536 12582
rect 9416 10220 9536 10248
rect 9416 9654 9444 10220
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9092 9276 9400 9285
rect 9092 9274 9098 9276
rect 9154 9274 9178 9276
rect 9234 9274 9258 9276
rect 9314 9274 9338 9276
rect 9394 9274 9400 9276
rect 9154 9222 9156 9274
rect 9336 9222 9338 9274
rect 9092 9220 9098 9222
rect 9154 9220 9178 9222
rect 9234 9220 9258 9222
rect 9314 9220 9338 9222
rect 9394 9220 9400 9222
rect 9092 9211 9400 9220
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 9092 8188 9400 8197
rect 9092 8186 9098 8188
rect 9154 8186 9178 8188
rect 9234 8186 9258 8188
rect 9314 8186 9338 8188
rect 9394 8186 9400 8188
rect 9154 8134 9156 8186
rect 9336 8134 9338 8186
rect 9092 8132 9098 8134
rect 9154 8132 9178 8134
rect 9234 8132 9258 8134
rect 9314 8132 9338 8134
rect 9394 8132 9400 8134
rect 9092 8123 9400 8132
rect 9092 7100 9400 7109
rect 9092 7098 9098 7100
rect 9154 7098 9178 7100
rect 9234 7098 9258 7100
rect 9314 7098 9338 7100
rect 9394 7098 9400 7100
rect 9154 7046 9156 7098
rect 9336 7046 9338 7098
rect 9092 7044 9098 7046
rect 9154 7044 9178 7046
rect 9234 7044 9258 7046
rect 9314 7044 9338 7046
rect 9394 7044 9400 7046
rect 9092 7035 9400 7044
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9092 6012 9400 6021
rect 9092 6010 9098 6012
rect 9154 6010 9178 6012
rect 9234 6010 9258 6012
rect 9314 6010 9338 6012
rect 9394 6010 9400 6012
rect 9154 5958 9156 6010
rect 9336 5958 9338 6010
rect 9092 5956 9098 5958
rect 9154 5956 9178 5958
rect 9234 5956 9258 5958
rect 9314 5956 9338 5958
rect 9394 5956 9400 5958
rect 9092 5947 9400 5956
rect 9508 5710 9536 6190
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 9508 5166 9536 5646
rect 9600 5574 9628 13126
rect 9692 12986 9720 13806
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12442 9720 12582
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10606 9720 11086
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9692 10062 9720 10542
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9518 9720 9998
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9042 9720 9454
rect 9784 9382 9812 12854
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9876 12238 9904 12650
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 10336 11830 10364 13874
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10796 13326 10824 13670
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10520 12442 10548 12854
rect 10796 12850 10824 13126
rect 10888 12850 10916 13466
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10980 12374 11008 13262
rect 11072 12986 11100 13398
rect 11164 13258 11192 13670
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8498 9720 8978
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9692 7954 9720 8434
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7478 9720 7890
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9680 7472 9732 7478
rect 10244 7449 10272 7754
rect 9680 7414 9732 7420
rect 10230 7440 10286 7449
rect 9692 6866 9720 7414
rect 10230 7375 10286 7384
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 10520 6730 10548 12174
rect 11072 11898 11100 12786
rect 11532 12782 11560 13126
rect 11716 12850 11744 13262
rect 11806 13084 12114 13093
rect 11806 13082 11812 13084
rect 11868 13082 11892 13084
rect 11948 13082 11972 13084
rect 12028 13082 12052 13084
rect 12108 13082 12114 13084
rect 11868 13030 11870 13082
rect 12050 13030 12052 13082
rect 11806 13028 11812 13030
rect 11868 13028 11892 13030
rect 11948 13028 11972 13030
rect 12028 13028 12052 13030
rect 12108 13028 12114 13030
rect 11806 13019 12114 13028
rect 12176 12850 12204 13330
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11164 12306 11192 12650
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11256 11898 11284 12038
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11348 11626 11376 12038
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 10810 11192 11494
rect 11348 11354 11376 11562
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11624 11082 11652 11698
rect 11716 11354 11744 12038
rect 11806 11996 12114 12005
rect 11806 11994 11812 11996
rect 11868 11994 11892 11996
rect 11948 11994 11972 11996
rect 12028 11994 12052 11996
rect 12108 11994 12114 11996
rect 11868 11942 11870 11994
rect 12050 11942 12052 11994
rect 11806 11940 11812 11942
rect 11868 11940 11892 11942
rect 11948 11940 11972 11942
rect 12028 11940 12052 11942
rect 12108 11940 12114 11942
rect 11806 11931 12114 11940
rect 12164 11756 12216 11762
rect 12268 11744 12296 13466
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 12360 12850 12388 13262
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12452 12918 12480 13194
rect 12636 12986 12756 13002
rect 12624 12980 12756 12986
rect 12676 12974 12756 12980
rect 12624 12922 12676 12928
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12442 12388 12786
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12360 12238 12388 12378
rect 12728 12238 12756 12974
rect 13280 12238 13308 13262
rect 14200 12850 14228 13262
rect 14292 12850 14320 13874
rect 14520 13628 14828 13637
rect 14520 13626 14526 13628
rect 14582 13626 14606 13628
rect 14662 13626 14686 13628
rect 14742 13626 14766 13628
rect 14822 13626 14828 13628
rect 14582 13574 14584 13626
rect 14764 13574 14766 13626
rect 14520 13572 14526 13574
rect 14582 13572 14606 13574
rect 14662 13572 14686 13574
rect 14742 13572 14766 13574
rect 14822 13572 14828 13574
rect 14520 13563 14828 13572
rect 19948 13628 20256 13637
rect 19948 13626 19954 13628
rect 20010 13626 20034 13628
rect 20090 13626 20114 13628
rect 20170 13626 20194 13628
rect 20250 13626 20256 13628
rect 20010 13574 20012 13626
rect 20192 13574 20194 13626
rect 19948 13572 19954 13574
rect 20010 13572 20034 13574
rect 20090 13572 20114 13574
rect 20170 13572 20194 13574
rect 20250 13572 20256 13574
rect 19948 13563 20256 13572
rect 17234 13084 17542 13093
rect 17234 13082 17240 13084
rect 17296 13082 17320 13084
rect 17376 13082 17400 13084
rect 17456 13082 17480 13084
rect 17536 13082 17542 13084
rect 17296 13030 17298 13082
rect 17478 13030 17480 13082
rect 17234 13028 17240 13030
rect 17296 13028 17320 13030
rect 17376 13028 17400 13030
rect 17456 13028 17480 13030
rect 17536 13028 17542 13030
rect 17234 13019 17542 13028
rect 22662 13084 22970 13093
rect 22662 13082 22668 13084
rect 22724 13082 22748 13084
rect 22804 13082 22828 13084
rect 22884 13082 22908 13084
rect 22964 13082 22970 13084
rect 22724 13030 22726 13082
rect 22906 13030 22908 13082
rect 22662 13028 22668 13030
rect 22724 13028 22748 13030
rect 22804 13028 22828 13030
rect 22884 13028 22908 13030
rect 22964 13028 22970 13030
rect 22662 13019 22970 13028
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12452 11762 12480 12106
rect 12216 11716 12296 11744
rect 12440 11756 12492 11762
rect 12164 11698 12216 11704
rect 12440 11698 12492 11704
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 11558 12112 11630
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11164 9994 11192 10746
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11624 8634 11652 11018
rect 11806 10908 12114 10917
rect 11806 10906 11812 10908
rect 11868 10906 11892 10908
rect 11948 10906 11972 10908
rect 12028 10906 12052 10908
rect 12108 10906 12114 10908
rect 11868 10854 11870 10906
rect 12050 10854 12052 10906
rect 11806 10852 11812 10854
rect 11868 10852 11892 10854
rect 11948 10852 11972 10854
rect 12028 10852 12052 10854
rect 12108 10852 12114 10854
rect 11806 10843 12114 10852
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10266 12112 10610
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12544 10062 12572 10406
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 11806 9820 12114 9829
rect 11806 9818 11812 9820
rect 11868 9818 11892 9820
rect 11948 9818 11972 9820
rect 12028 9818 12052 9820
rect 12108 9818 12114 9820
rect 11868 9766 11870 9818
rect 12050 9766 12052 9818
rect 11806 9764 11812 9766
rect 11868 9764 11892 9766
rect 11948 9764 11972 9766
rect 12028 9764 12052 9766
rect 12108 9764 12114 9766
rect 11806 9755 12114 9764
rect 11806 8732 12114 8741
rect 11806 8730 11812 8732
rect 11868 8730 11892 8732
rect 11948 8730 11972 8732
rect 12028 8730 12052 8732
rect 12108 8730 12114 8732
rect 11868 8678 11870 8730
rect 12050 8678 12052 8730
rect 11806 8676 11812 8678
rect 11868 8676 11892 8678
rect 11948 8676 11972 8678
rect 12028 8676 12052 8678
rect 12108 8676 12114 8678
rect 11806 8667 12114 8676
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 12728 8090 12756 12174
rect 13280 11762 13308 12174
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 8974 12940 9318
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 13280 8906 13308 11698
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 9654 13400 10542
rect 13464 10538 13492 12650
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13924 11558 13952 12106
rect 14200 11898 14228 12786
rect 14292 12306 14320 12786
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12306 14412 12582
rect 14520 12540 14828 12549
rect 14520 12538 14526 12540
rect 14582 12538 14606 12540
rect 14662 12538 14686 12540
rect 14742 12538 14766 12540
rect 14822 12538 14828 12540
rect 14582 12486 14584 12538
rect 14764 12486 14766 12538
rect 14520 12484 14526 12486
rect 14582 12484 14606 12486
rect 14662 12484 14686 12486
rect 14742 12484 14766 12486
rect 14822 12484 14828 12486
rect 14520 12475 14828 12484
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 14200 11082 14228 11630
rect 14292 11354 14320 12038
rect 14752 11898 14780 12174
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13832 10606 13860 10746
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13464 10130 13492 10474
rect 13832 10198 13860 10542
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13464 10010 13492 10066
rect 13464 9982 13584 10010
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13372 9042 13400 9590
rect 13556 9518 13584 9982
rect 13832 9518 13860 10134
rect 14200 10062 14228 11018
rect 14384 10810 14412 11698
rect 14520 11452 14828 11461
rect 14520 11450 14526 11452
rect 14582 11450 14606 11452
rect 14662 11450 14686 11452
rect 14742 11450 14766 11452
rect 14822 11450 14828 11452
rect 14582 11398 14584 11450
rect 14764 11398 14766 11450
rect 14520 11396 14526 11398
rect 14582 11396 14606 11398
rect 14662 11396 14686 11398
rect 14742 11396 14766 11398
rect 14822 11396 14828 11398
rect 14520 11387 14828 11396
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14384 10130 14412 10746
rect 14936 10742 14964 12038
rect 15028 10742 15056 12242
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15212 11218 15240 11698
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14520 10364 14828 10373
rect 14520 10362 14526 10364
rect 14582 10362 14606 10364
rect 14662 10362 14686 10364
rect 14742 10362 14766 10364
rect 14822 10362 14828 10364
rect 14582 10310 14584 10362
rect 14764 10310 14766 10362
rect 14520 10308 14526 10310
rect 14582 10308 14606 10310
rect 14662 10308 14686 10310
rect 14742 10308 14766 10310
rect 14822 10308 14828 10310
rect 14520 10299 14828 10308
rect 14936 10130 14964 10406
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13832 8906 13860 9454
rect 14292 9178 14320 9930
rect 14936 9586 14964 10066
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 15028 9450 15056 10678
rect 15212 10674 15240 11154
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 10577 15240 10610
rect 15198 10568 15254 10577
rect 15198 10503 15254 10512
rect 16224 10062 16252 12310
rect 16960 10062 16988 12854
rect 19948 12540 20256 12549
rect 19948 12538 19954 12540
rect 20010 12538 20034 12540
rect 20090 12538 20114 12540
rect 20170 12538 20194 12540
rect 20250 12538 20256 12540
rect 20010 12486 20012 12538
rect 20192 12486 20194 12538
rect 19948 12484 19954 12486
rect 20010 12484 20034 12486
rect 20090 12484 20114 12486
rect 20170 12484 20194 12486
rect 20250 12484 20256 12486
rect 19948 12475 20256 12484
rect 17234 11996 17542 12005
rect 17234 11994 17240 11996
rect 17296 11994 17320 11996
rect 17376 11994 17400 11996
rect 17456 11994 17480 11996
rect 17536 11994 17542 11996
rect 17296 11942 17298 11994
rect 17478 11942 17480 11994
rect 17234 11940 17240 11942
rect 17296 11940 17320 11942
rect 17376 11940 17400 11942
rect 17456 11940 17480 11942
rect 17536 11940 17542 11942
rect 17234 11931 17542 11940
rect 22662 11996 22970 12005
rect 22662 11994 22668 11996
rect 22724 11994 22748 11996
rect 22804 11994 22828 11996
rect 22884 11994 22908 11996
rect 22964 11994 22970 11996
rect 22724 11942 22726 11994
rect 22906 11942 22908 11994
rect 22662 11940 22668 11942
rect 22724 11940 22748 11942
rect 22804 11940 22828 11942
rect 22884 11940 22908 11942
rect 22964 11940 22970 11942
rect 22662 11931 22970 11940
rect 19948 11452 20256 11461
rect 19948 11450 19954 11452
rect 20010 11450 20034 11452
rect 20090 11450 20114 11452
rect 20170 11450 20194 11452
rect 20250 11450 20256 11452
rect 20010 11398 20012 11450
rect 20192 11398 20194 11450
rect 19948 11396 19954 11398
rect 20010 11396 20034 11398
rect 20090 11396 20114 11398
rect 20170 11396 20194 11398
rect 20250 11396 20256 11398
rect 19948 11387 20256 11396
rect 17234 10908 17542 10917
rect 17234 10906 17240 10908
rect 17296 10906 17320 10908
rect 17376 10906 17400 10908
rect 17456 10906 17480 10908
rect 17536 10906 17542 10908
rect 17296 10854 17298 10906
rect 17478 10854 17480 10906
rect 17234 10852 17240 10854
rect 17296 10852 17320 10854
rect 17376 10852 17400 10854
rect 17456 10852 17480 10854
rect 17536 10852 17542 10854
rect 17234 10843 17542 10852
rect 22662 10908 22970 10917
rect 22662 10906 22668 10908
rect 22724 10906 22748 10908
rect 22804 10906 22828 10908
rect 22884 10906 22908 10908
rect 22964 10906 22970 10908
rect 22724 10854 22726 10906
rect 22906 10854 22908 10906
rect 22662 10852 22668 10854
rect 22724 10852 22748 10854
rect 22804 10852 22828 10854
rect 22884 10852 22908 10854
rect 22964 10852 22970 10854
rect 22662 10843 22970 10852
rect 19948 10364 20256 10373
rect 19948 10362 19954 10364
rect 20010 10362 20034 10364
rect 20090 10362 20114 10364
rect 20170 10362 20194 10364
rect 20250 10362 20256 10364
rect 20010 10310 20012 10362
rect 20192 10310 20194 10362
rect 19948 10308 19954 10310
rect 20010 10308 20034 10310
rect 20090 10308 20114 10310
rect 20170 10308 20194 10310
rect 20250 10308 20256 10310
rect 19948 10299 20256 10308
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14520 9276 14828 9285
rect 14520 9274 14526 9276
rect 14582 9274 14606 9276
rect 14662 9274 14686 9276
rect 14742 9274 14766 9276
rect 14822 9274 14828 9276
rect 14582 9222 14584 9274
rect 14764 9222 14766 9274
rect 14520 9220 14526 9222
rect 14582 9220 14606 9222
rect 14662 9220 14686 9222
rect 14742 9220 14766 9222
rect 14822 9220 14828 9222
rect 14520 9211 14828 9220
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 11806 7644 12114 7653
rect 11806 7642 11812 7644
rect 11868 7642 11892 7644
rect 11948 7642 11972 7644
rect 12028 7642 12052 7644
rect 12108 7642 12114 7644
rect 11868 7590 11870 7642
rect 12050 7590 12052 7642
rect 11806 7588 11812 7590
rect 11868 7588 11892 7590
rect 11948 7588 11972 7590
rect 12028 7588 12052 7590
rect 12108 7588 12114 7590
rect 11806 7579 12114 7588
rect 12636 7410 12664 7686
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 6798 11284 7142
rect 11244 6792 11296 6798
rect 11150 6760 11206 6769
rect 10508 6724 10560 6730
rect 11244 6734 11296 6740
rect 11150 6695 11206 6704
rect 10508 6666 10560 6672
rect 11164 6662 11192 6695
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11806 6556 12114 6565
rect 11806 6554 11812 6556
rect 11868 6554 11892 6556
rect 11948 6554 11972 6556
rect 12028 6554 12052 6556
rect 12108 6554 12114 6556
rect 11868 6502 11870 6554
rect 12050 6502 12052 6554
rect 11806 6500 11812 6502
rect 11868 6500 11892 6502
rect 11948 6500 11972 6502
rect 12028 6500 12052 6502
rect 12108 6500 12114 6502
rect 11806 6491 12114 6500
rect 12360 6458 12388 7210
rect 12636 6730 12664 7346
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 11716 5234 11744 5646
rect 11806 5468 12114 5477
rect 11806 5466 11812 5468
rect 11868 5466 11892 5468
rect 11948 5466 11972 5468
rect 12028 5466 12052 5468
rect 12108 5466 12114 5468
rect 11868 5414 11870 5466
rect 12050 5414 12052 5466
rect 11806 5412 11812 5414
rect 11868 5412 11892 5414
rect 11948 5412 11972 5414
rect 12028 5412 12052 5414
rect 12108 5412 12114 5414
rect 11806 5403 12114 5412
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7484 2990 7512 4762
rect 7576 4486 7604 4966
rect 9092 4924 9400 4933
rect 9092 4922 9098 4924
rect 9154 4922 9178 4924
rect 9234 4922 9258 4924
rect 9314 4922 9338 4924
rect 9394 4922 9400 4924
rect 9154 4870 9156 4922
rect 9336 4870 9338 4922
rect 9092 4868 9098 4870
rect 9154 4868 9178 4870
rect 9234 4868 9258 4870
rect 9314 4868 9338 4870
rect 9394 4868 9400 4870
rect 9092 4859 9400 4868
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 9508 4146 9536 5102
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4690 11192 4966
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 4146 11100 4490
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7472 2848 7524 2854
rect 7576 2802 7604 2994
rect 7852 2922 7880 3878
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 7524 2796 7604 2802
rect 7472 2790 7604 2796
rect 7484 2774 7604 2790
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7484 2446 7512 2774
rect 8036 2650 8064 4082
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8128 2582 8156 3334
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8128 2446 8156 2518
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7944 2258 7972 2314
rect 8220 2310 8248 3130
rect 8956 2650 8984 4082
rect 9092 3836 9400 3845
rect 9092 3834 9098 3836
rect 9154 3834 9178 3836
rect 9234 3834 9258 3836
rect 9314 3834 9338 3836
rect 9394 3834 9400 3836
rect 9154 3782 9156 3834
rect 9336 3782 9338 3834
rect 9092 3780 9098 3782
rect 9154 3780 9178 3782
rect 9234 3780 9258 3782
rect 9314 3780 9338 3782
rect 9394 3780 9400 3782
rect 9092 3771 9400 3780
rect 9508 3602 9536 4082
rect 11716 3670 11744 4626
rect 11806 4380 12114 4389
rect 11806 4378 11812 4380
rect 11868 4378 11892 4380
rect 11948 4378 11972 4380
rect 12028 4378 12052 4380
rect 12108 4378 12114 4380
rect 11868 4326 11870 4378
rect 12050 4326 12052 4378
rect 11806 4324 11812 4326
rect 11868 4324 11892 4326
rect 11948 4324 11972 4326
rect 12028 4324 12052 4326
rect 12108 4324 12114 4326
rect 11806 4315 12114 4324
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9508 3126 9536 3538
rect 12084 3466 12112 3878
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9092 2748 9400 2757
rect 9092 2746 9098 2748
rect 9154 2746 9178 2748
rect 9234 2746 9258 2748
rect 9314 2746 9338 2748
rect 9394 2746 9400 2748
rect 9154 2694 9156 2746
rect 9336 2694 9338 2746
rect 9092 2692 9098 2694
rect 9154 2692 9178 2694
rect 9234 2692 9258 2694
rect 9314 2692 9338 2694
rect 9394 2692 9400 2694
rect 9092 2683 9400 2692
rect 9508 2650 9536 2926
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 10060 2514 10088 2790
rect 11072 2650 11100 3402
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3126 11192 3334
rect 11806 3292 12114 3301
rect 11806 3290 11812 3292
rect 11868 3290 11892 3292
rect 11948 3290 11972 3292
rect 12028 3290 12052 3292
rect 12108 3290 12114 3292
rect 11868 3238 11870 3290
rect 12050 3238 12052 3290
rect 11806 3236 11812 3238
rect 11868 3236 11892 3238
rect 11948 3236 11972 3238
rect 12028 3236 12052 3238
rect 12108 3236 12114 3238
rect 11806 3227 12114 3236
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 11164 2378 11192 2790
rect 11716 2446 11744 2790
rect 12176 2650 12204 4082
rect 12360 3534 12388 6394
rect 12636 6118 12664 6666
rect 12912 6254 12940 7822
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12360 3194 12388 3470
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12452 2922 12480 3674
rect 12636 3398 12664 6054
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5370 12756 5646
rect 12820 5574 12848 5850
rect 13004 5846 13032 7890
rect 13280 7886 13308 8502
rect 14384 8498 14412 9114
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7410 13308 7686
rect 13372 7410 13400 8230
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13556 7342 13584 7686
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13648 7206 13676 7822
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13084 6656 13136 6662
rect 13136 6604 13216 6610
rect 13084 6598 13216 6604
rect 13096 6582 13216 6598
rect 13188 6254 13216 6582
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 13004 5234 13032 5782
rect 13096 5642 13124 6190
rect 13188 5710 13216 6190
rect 13280 5846 13308 6734
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 4146 13032 5170
rect 13096 4162 13124 5578
rect 13280 5234 13308 5782
rect 13464 5574 13492 6054
rect 13556 5914 13584 6666
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13556 4826 13584 5850
rect 13648 5778 13676 7142
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 12992 4140 13044 4146
rect 13096 4134 13216 4162
rect 12992 4082 13044 4088
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 13004 3058 13032 4082
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3738 13124 4014
rect 13188 4010 13216 4134
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13280 3618 13308 3878
rect 13740 3618 13768 7822
rect 13924 6798 13952 8434
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14016 7818 14044 8366
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 7546 14044 7754
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13832 4622 13860 5238
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13924 4049 13952 6734
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6322 14044 6666
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14016 5370 14044 6122
rect 14108 5914 14136 8434
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5794 14228 8434
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 14520 8188 14828 8197
rect 14520 8186 14526 8188
rect 14582 8186 14606 8188
rect 14662 8186 14686 8188
rect 14742 8186 14766 8188
rect 14822 8186 14828 8188
rect 14582 8134 14584 8186
rect 14764 8134 14766 8186
rect 14520 8132 14526 8134
rect 14582 8132 14606 8134
rect 14662 8132 14686 8134
rect 14742 8132 14766 8134
rect 14822 8132 14828 8134
rect 14520 8123 14828 8132
rect 15212 8090 15240 8298
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7410 15056 7686
rect 15212 7410 15240 7822
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 14520 7100 14828 7109
rect 14520 7098 14526 7100
rect 14582 7098 14606 7100
rect 14662 7098 14686 7100
rect 14742 7098 14766 7100
rect 14822 7098 14828 7100
rect 14582 7046 14584 7098
rect 14764 7046 14766 7098
rect 14520 7044 14526 7046
rect 14582 7044 14606 7046
rect 14662 7044 14686 7046
rect 14742 7044 14766 7046
rect 14822 7044 14828 7046
rect 14520 7035 14828 7044
rect 15212 7002 15240 7346
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14384 5914 14412 6122
rect 14520 6012 14828 6021
rect 14520 6010 14526 6012
rect 14582 6010 14606 6012
rect 14662 6010 14686 6012
rect 14742 6010 14766 6012
rect 14822 6010 14828 6012
rect 14582 5958 14584 6010
rect 14764 5958 14766 6010
rect 14520 5956 14526 5958
rect 14582 5956 14606 5958
rect 14662 5956 14686 5958
rect 14742 5956 14766 5958
rect 14822 5956 14828 5958
rect 14520 5947 14828 5956
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14108 5766 14228 5794
rect 14384 5778 14412 5850
rect 14372 5772 14424 5778
rect 14108 5642 14136 5766
rect 14372 5714 14424 5720
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14200 4826 14228 5646
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4146 14228 4422
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13910 4040 13966 4049
rect 13910 3975 13966 3984
rect 13924 3942 13952 3975
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13096 3602 13768 3618
rect 13084 3596 13780 3602
rect 13136 3590 13728 3596
rect 13084 3538 13136 3544
rect 13728 3538 13780 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 14292 3516 14320 5102
rect 14384 4690 14412 5170
rect 14520 4924 14828 4933
rect 14520 4922 14526 4924
rect 14582 4922 14606 4924
rect 14662 4922 14686 4924
rect 14742 4922 14766 4924
rect 14822 4922 14828 4924
rect 14582 4870 14584 4922
rect 14764 4870 14766 4922
rect 14520 4868 14526 4870
rect 14582 4868 14606 4870
rect 14662 4868 14686 4870
rect 14742 4868 14766 4870
rect 14822 4868 14828 4870
rect 14520 4859 14828 4868
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14844 4214 14872 4558
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14520 3836 14828 3845
rect 14520 3834 14526 3836
rect 14582 3834 14606 3836
rect 14662 3834 14686 3836
rect 14742 3834 14766 3836
rect 14822 3834 14828 3836
rect 14582 3782 14584 3834
rect 14764 3782 14766 3834
rect 14520 3780 14526 3782
rect 14582 3780 14606 3782
rect 14662 3780 14686 3782
rect 14742 3780 14766 3782
rect 14822 3780 14828 3782
rect 14520 3771 14828 3780
rect 14936 3738 14964 5714
rect 15028 5710 15056 6598
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15028 5302 15056 5646
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 15028 4758 15056 5102
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15212 4690 15240 5170
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15212 4282 15240 4626
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15120 3534 15148 3878
rect 15304 3670 15332 9522
rect 15672 9042 15700 9862
rect 16224 9586 16252 9998
rect 16592 9654 16620 9998
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8566 15700 8978
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 7886 15516 8434
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 7954 15700 8366
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7750 15516 7822
rect 15672 7818 15700 7890
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15764 6934 15792 7890
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15672 6322 15700 6666
rect 15764 6390 15792 6870
rect 15948 6798 15976 7686
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 16040 7342 16068 7414
rect 16132 7410 16160 8910
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16224 8498 16252 8774
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16316 7954 16344 8774
rect 16408 8566 16436 8842
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15936 6792 15988 6798
rect 15856 6740 15936 6746
rect 15856 6734 15988 6740
rect 15856 6718 15976 6734
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15856 6202 15884 6718
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15764 6174 15884 6202
rect 15764 5710 15792 6174
rect 15948 5846 15976 6258
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15764 4146 15792 5646
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15856 4826 15884 5170
rect 16040 4826 16068 7142
rect 16132 6934 16160 7346
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16132 6730 16160 6870
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16408 6458 16436 8502
rect 16500 8090 16528 8842
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16500 6798 16528 8026
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16408 6118 16436 6394
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5710 16436 6054
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 5302 16436 5646
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 14372 3528 14424 3534
rect 14292 3488 14372 3516
rect 13648 3058 13676 3470
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12912 2446 12940 2790
rect 13096 2650 13124 2926
rect 14292 2922 14320 3488
rect 14372 3470 14424 3476
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15212 3126 15240 3538
rect 15304 3194 15332 3606
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15304 2990 15332 3130
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 15304 2774 15332 2926
rect 14520 2748 14828 2757
rect 14520 2746 14526 2748
rect 14582 2746 14606 2748
rect 14662 2746 14686 2748
rect 14742 2746 14766 2748
rect 14822 2746 14828 2748
rect 15304 2746 15516 2774
rect 14582 2694 14584 2746
rect 14764 2694 14766 2746
rect 14520 2692 14526 2694
rect 14582 2692 14606 2694
rect 14662 2692 14686 2694
rect 14742 2692 14766 2694
rect 14822 2692 14828 2694
rect 14520 2683 14828 2692
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 15488 2446 15516 2746
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 15580 2310 15608 4082
rect 15764 4010 15792 4082
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15856 3670 15884 4762
rect 16408 4622 16436 5238
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16500 4146 16528 6734
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15948 3058 15976 3402
rect 16592 3398 16620 9590
rect 16960 9450 16988 9998
rect 17234 9820 17542 9829
rect 17234 9818 17240 9820
rect 17296 9818 17320 9820
rect 17376 9818 17400 9820
rect 17456 9818 17480 9820
rect 17536 9818 17542 9820
rect 17296 9766 17298 9818
rect 17478 9766 17480 9818
rect 17234 9764 17240 9766
rect 17296 9764 17320 9766
rect 17376 9764 17400 9766
rect 17456 9764 17480 9766
rect 17536 9764 17542 9766
rect 17234 9755 17542 9764
rect 22662 9820 22970 9829
rect 22662 9818 22668 9820
rect 22724 9818 22748 9820
rect 22804 9818 22828 9820
rect 22884 9818 22908 9820
rect 22964 9818 22970 9820
rect 22724 9766 22726 9818
rect 22906 9766 22908 9818
rect 22662 9764 22668 9766
rect 22724 9764 22748 9766
rect 22804 9764 22828 9766
rect 22884 9764 22908 9766
rect 22964 9764 22970 9766
rect 22662 9755 22970 9764
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 7886 16712 8366
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 5778 16712 7822
rect 16776 7274 16804 8910
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16960 8430 16988 8842
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 6730 16988 7142
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16960 6322 16988 6666
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16776 5710 16804 5850
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16776 5522 16804 5646
rect 16868 5574 16896 6258
rect 16960 5710 16988 6258
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16684 5494 16804 5522
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16684 4826 16712 5494
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16776 4622 16804 5238
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16776 3398 16804 4558
rect 17052 4146 17080 9318
rect 19948 9276 20256 9285
rect 19948 9274 19954 9276
rect 20010 9274 20034 9276
rect 20090 9274 20114 9276
rect 20170 9274 20194 9276
rect 20250 9274 20256 9276
rect 20010 9222 20012 9274
rect 20192 9222 20194 9274
rect 19948 9220 19954 9222
rect 20010 9220 20034 9222
rect 20090 9220 20114 9222
rect 20170 9220 20194 9222
rect 20250 9220 20256 9222
rect 19948 9211 20256 9220
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17234 8732 17542 8741
rect 17234 8730 17240 8732
rect 17296 8730 17320 8732
rect 17376 8730 17400 8732
rect 17456 8730 17480 8732
rect 17536 8730 17542 8732
rect 17296 8678 17298 8730
rect 17478 8678 17480 8730
rect 17234 8676 17240 8678
rect 17296 8676 17320 8678
rect 17376 8676 17400 8678
rect 17456 8676 17480 8678
rect 17536 8676 17542 8678
rect 17234 8667 17542 8676
rect 17696 8498 17724 9114
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17144 7546 17172 8366
rect 17696 8294 17724 8434
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17512 7750 17540 7958
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17234 7644 17542 7653
rect 17234 7642 17240 7644
rect 17296 7642 17320 7644
rect 17376 7642 17400 7644
rect 17456 7642 17480 7644
rect 17536 7642 17542 7644
rect 17296 7590 17298 7642
rect 17478 7590 17480 7642
rect 17234 7588 17240 7590
rect 17296 7588 17320 7590
rect 17376 7588 17400 7590
rect 17456 7588 17480 7590
rect 17536 7588 17542 7590
rect 17234 7579 17542 7588
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17420 7449 17448 7482
rect 17406 7440 17462 7449
rect 17406 7375 17462 7384
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17234 6556 17542 6565
rect 17234 6554 17240 6556
rect 17296 6554 17320 6556
rect 17376 6554 17400 6556
rect 17456 6554 17480 6556
rect 17536 6554 17542 6556
rect 17296 6502 17298 6554
rect 17478 6502 17480 6554
rect 17234 6500 17240 6502
rect 17296 6500 17320 6502
rect 17376 6500 17400 6502
rect 17456 6500 17480 6502
rect 17536 6500 17542 6502
rect 17234 6491 17542 6500
rect 17604 6458 17632 7278
rect 17696 6458 17724 7890
rect 17788 7818 17816 8910
rect 18064 8634 18092 8910
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18432 7818 18460 8298
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7478 18000 7686
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 17788 6934 17816 7278
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17788 6798 17816 6870
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17328 5914 17356 6258
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17696 5794 17724 6394
rect 17880 5846 17908 7142
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17868 5840 17920 5846
rect 17696 5766 17816 5794
rect 17868 5782 17920 5788
rect 17788 5710 17816 5766
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17234 5468 17542 5477
rect 17234 5466 17240 5468
rect 17296 5466 17320 5468
rect 17376 5466 17400 5468
rect 17456 5466 17480 5468
rect 17536 5466 17542 5468
rect 17296 5414 17298 5466
rect 17478 5414 17480 5466
rect 17234 5412 17240 5414
rect 17296 5412 17320 5414
rect 17376 5412 17400 5414
rect 17456 5412 17480 5414
rect 17536 5412 17542 5414
rect 17234 5403 17542 5412
rect 17696 5302 17724 5646
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17696 4622 17724 5102
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17234 4380 17542 4389
rect 17234 4378 17240 4380
rect 17296 4378 17320 4380
rect 17376 4378 17400 4380
rect 17456 4378 17480 4380
rect 17536 4378 17542 4380
rect 17296 4326 17298 4378
rect 17478 4326 17480 4378
rect 17234 4324 17240 4326
rect 17296 4324 17320 4326
rect 17376 4324 17400 4326
rect 17456 4324 17480 4326
rect 17536 4324 17542 4326
rect 17234 4315 17542 4324
rect 17788 4146 17816 4966
rect 17880 4758 17908 5782
rect 17972 4826 18000 6326
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 18064 5710 18092 6054
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18156 5574 18184 5714
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 17880 4146 17908 4694
rect 18156 4282 18184 5170
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15764 2378 15792 2790
rect 15856 2378 15884 2994
rect 15948 2650 15976 2994
rect 16592 2990 16620 3334
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 16040 2310 16068 2450
rect 16776 2310 16804 3334
rect 16868 2854 16896 3538
rect 16960 3534 16988 4082
rect 17052 3738 17080 4082
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17328 3738 17356 3878
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17788 3466 17816 4082
rect 17880 3534 17908 4082
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17234 3292 17542 3301
rect 17234 3290 17240 3292
rect 17296 3290 17320 3292
rect 17376 3290 17400 3292
rect 17456 3290 17480 3292
rect 17536 3290 17542 3292
rect 17296 3238 17298 3290
rect 17478 3238 17480 3290
rect 17234 3236 17240 3238
rect 17296 3236 17320 3238
rect 17376 3236 17400 3238
rect 17456 3236 17480 3238
rect 17536 3236 17542 3238
rect 17234 3227 17542 3236
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16960 2446 16988 2926
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17236 2446 17264 2790
rect 17880 2650 17908 3470
rect 18248 3194 18276 7278
rect 18432 6866 18460 7754
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18432 6254 18460 6802
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18432 4826 18460 5578
rect 18524 5234 18552 7414
rect 18616 7410 18644 9046
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18984 8498 19012 8842
rect 19628 8634 19656 9046
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18708 7274 18736 7346
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18708 6866 18736 7210
rect 18696 6860 18748 6866
rect 18748 6820 18828 6848
rect 18696 6802 18748 6808
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18616 5098 18644 6054
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 3942 18368 4422
rect 18524 4078 18552 4626
rect 18708 4622 18736 6190
rect 18800 5166 18828 6820
rect 18892 6798 18920 8298
rect 18984 8090 19012 8434
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 19076 7410 19104 8230
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18892 6390 18920 6734
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18800 4434 18828 4966
rect 18708 4406 18828 4434
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 3670 18368 3878
rect 18432 3670 18460 3946
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18524 3194 18552 4014
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18708 3058 18736 4406
rect 18892 3534 18920 5714
rect 18984 5370 19012 6258
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 19076 5030 19104 7346
rect 19168 6934 19196 8434
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 7478 19380 7822
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19168 5778 19196 6870
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19260 5370 19288 6190
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19352 5234 19380 6598
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19444 5914 19472 6258
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19430 5808 19486 5817
rect 19536 5794 19564 8434
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19628 6361 19656 8298
rect 19720 7750 19748 8910
rect 22662 8732 22970 8741
rect 22662 8730 22668 8732
rect 22724 8730 22748 8732
rect 22804 8730 22828 8732
rect 22884 8730 22908 8732
rect 22964 8730 22970 8732
rect 22724 8678 22726 8730
rect 22906 8678 22908 8730
rect 22662 8676 22668 8678
rect 22724 8676 22748 8678
rect 22804 8676 22828 8678
rect 22884 8676 22908 8678
rect 22964 8676 22970 8678
rect 22662 8667 22970 8676
rect 19904 8634 20116 8650
rect 19904 8628 20128 8634
rect 19904 8622 20076 8628
rect 19904 8566 19932 8622
rect 20076 8570 20128 8576
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 19812 8090 19840 8434
rect 20088 8362 20116 8434
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19948 8188 20256 8197
rect 19948 8186 19954 8188
rect 20010 8186 20034 8188
rect 20090 8186 20114 8188
rect 20170 8186 20194 8188
rect 20250 8186 20256 8188
rect 20010 8134 20012 8186
rect 20192 8134 20194 8186
rect 19948 8132 19954 8134
rect 20010 8132 20034 8134
rect 20090 8132 20114 8134
rect 20170 8132 20194 8134
rect 20250 8132 20256 8134
rect 19948 8123 20256 8132
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 6798 19748 7686
rect 19812 6866 19840 7890
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 7274 20208 7822
rect 20364 7478 20392 8434
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19948 7100 20256 7109
rect 19948 7098 19954 7100
rect 20010 7098 20034 7100
rect 20090 7098 20114 7100
rect 20170 7098 20194 7100
rect 20250 7098 20256 7100
rect 20010 7046 20012 7098
rect 20192 7046 20194 7098
rect 19948 7044 19954 7046
rect 20010 7044 20034 7046
rect 20090 7044 20114 7046
rect 20170 7044 20194 7046
rect 20250 7044 20256 7046
rect 19948 7035 20256 7044
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19614 6352 19670 6361
rect 19812 6338 19840 6802
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19614 6287 19670 6296
rect 19720 6310 19840 6338
rect 20088 6322 20116 6394
rect 20076 6316 20128 6322
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 19628 5914 19656 6122
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19536 5766 19656 5794
rect 19430 5743 19486 5752
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19444 4706 19472 5743
rect 19628 5710 19656 5766
rect 19616 5704 19668 5710
rect 19614 5672 19616 5681
rect 19668 5672 19670 5681
rect 19614 5607 19670 5616
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19536 5234 19564 5510
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19444 4678 19564 4706
rect 19536 4622 19564 4678
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 4078 19380 4490
rect 19340 4072 19392 4078
rect 19062 4040 19118 4049
rect 19340 4014 19392 4020
rect 19062 3975 19118 3984
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3058 18920 3334
rect 19076 3058 19104 3975
rect 19536 3670 19564 4558
rect 19720 3738 19748 6310
rect 20076 6258 20128 6264
rect 20364 6254 20392 7142
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19812 5302 19840 6122
rect 19948 6012 20256 6021
rect 19948 6010 19954 6012
rect 20010 6010 20034 6012
rect 20090 6010 20114 6012
rect 20170 6010 20194 6012
rect 20250 6010 20256 6012
rect 20010 5958 20012 6010
rect 20192 5958 20194 6010
rect 19948 5956 19954 5958
rect 20010 5956 20034 5958
rect 20090 5956 20114 5958
rect 20170 5956 20194 5958
rect 20250 5956 20256 5958
rect 19948 5947 20256 5956
rect 20364 5846 20392 6190
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20456 5710 20484 8366
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20548 6458 20576 7822
rect 22662 7644 22970 7653
rect 22662 7642 22668 7644
rect 22724 7642 22748 7644
rect 22804 7642 22828 7644
rect 22884 7642 22908 7644
rect 22964 7642 22970 7644
rect 22724 7590 22726 7642
rect 22906 7590 22908 7642
rect 22662 7588 22668 7590
rect 22724 7588 22748 7590
rect 22804 7588 22828 7590
rect 22884 7588 22908 7590
rect 22964 7588 22970 7590
rect 22662 7579 22970 7588
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20536 6452 20588 6458
rect 20588 6412 20668 6440
rect 20536 6394 20588 6400
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5778 20576 6054
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20352 5636 20404 5642
rect 20352 5578 20404 5584
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19948 4924 20256 4933
rect 19948 4922 19954 4924
rect 20010 4922 20034 4924
rect 20090 4922 20114 4924
rect 20170 4922 20194 4924
rect 20250 4922 20256 4924
rect 20010 4870 20012 4922
rect 20192 4870 20194 4922
rect 19948 4868 19954 4870
rect 20010 4868 20034 4870
rect 20090 4868 20114 4870
rect 20170 4868 20194 4870
rect 20250 4868 20256 4870
rect 19948 4859 20256 4868
rect 19948 3836 20256 3845
rect 19948 3834 19954 3836
rect 20010 3834 20034 3836
rect 20090 3834 20114 3836
rect 20170 3834 20194 3836
rect 20250 3834 20256 3836
rect 20010 3782 20012 3834
rect 20192 3782 20194 3834
rect 19948 3780 19954 3782
rect 20010 3780 20034 3782
rect 20090 3780 20114 3782
rect 20170 3780 20194 3782
rect 20250 3780 20256 3782
rect 19948 3771 20256 3780
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19720 3618 19748 3674
rect 20260 3664 20312 3670
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19352 3398 19380 3538
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19352 2854 19380 3334
rect 19536 3058 19564 3606
rect 19720 3590 19840 3618
rect 20260 3606 20312 3612
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 18616 2514 18644 2790
rect 19720 2650 19748 3130
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 19812 2310 19840 3590
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19996 3194 20024 3402
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20272 2990 20300 3606
rect 20364 3466 20392 5578
rect 20456 4826 20484 5646
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20548 3942 20576 5714
rect 20640 5710 20668 6412
rect 20824 6322 20852 6666
rect 22662 6556 22970 6565
rect 22662 6554 22668 6556
rect 22724 6554 22748 6556
rect 22804 6554 22828 6556
rect 22884 6554 22908 6556
rect 22964 6554 22970 6556
rect 22724 6502 22726 6554
rect 22906 6502 22908 6554
rect 22662 6500 22668 6502
rect 22724 6500 22748 6502
rect 22804 6500 22828 6502
rect 22884 6500 22908 6502
rect 22964 6500 22970 6502
rect 22662 6491 22970 6500
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20640 5302 20668 5510
rect 22662 5468 22970 5477
rect 22662 5466 22668 5468
rect 22724 5466 22748 5468
rect 22804 5466 22828 5468
rect 22884 5466 22908 5468
rect 22964 5466 22970 5468
rect 22724 5414 22726 5466
rect 22906 5414 22908 5466
rect 22662 5412 22668 5414
rect 22724 5412 22748 5414
rect 22804 5412 22828 5414
rect 22884 5412 22908 5414
rect 22964 5412 22970 5414
rect 22662 5403 22970 5412
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 22662 4380 22970 4389
rect 22662 4378 22668 4380
rect 22724 4378 22748 4380
rect 22804 4378 22828 4380
rect 22884 4378 22908 4380
rect 22964 4378 22970 4380
rect 22724 4326 22726 4378
rect 22906 4326 22908 4378
rect 22662 4324 22668 4326
rect 22724 4324 22748 4326
rect 22804 4324 22828 4326
rect 22884 4324 22908 4326
rect 22964 4324 22970 4326
rect 22662 4315 22970 4324
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20548 3534 20576 3878
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 22662 3292 22970 3301
rect 22662 3290 22668 3292
rect 22724 3290 22748 3292
rect 22804 3290 22828 3292
rect 22884 3290 22908 3292
rect 22964 3290 22970 3292
rect 22724 3238 22726 3290
rect 22906 3238 22908 3290
rect 22662 3236 22668 3238
rect 22724 3236 22748 3238
rect 22804 3236 22828 3238
rect 22884 3236 22908 3238
rect 22964 3236 22970 3238
rect 22662 3227 22970 3236
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 19948 2748 20256 2757
rect 19948 2746 19954 2748
rect 20010 2746 20034 2748
rect 20090 2746 20114 2748
rect 20170 2746 20194 2748
rect 20250 2746 20256 2748
rect 20010 2694 20012 2746
rect 20192 2694 20194 2746
rect 19948 2692 19954 2694
rect 20010 2692 20034 2694
rect 20090 2692 20114 2694
rect 20170 2692 20194 2694
rect 20250 2692 20256 2694
rect 19948 2683 20256 2692
rect 8208 2304 8260 2310
rect 7944 2252 8208 2258
rect 7944 2246 8260 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 19800 2304 19852 2310
rect 19800 2246 19852 2252
rect 7944 2230 8248 2246
rect 6378 2204 6686 2213
rect 6378 2202 6384 2204
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6680 2202 6686 2204
rect 6440 2150 6442 2202
rect 6622 2150 6624 2202
rect 6378 2148 6384 2150
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6680 2148 6686 2150
rect 6378 2139 6686 2148
rect 11806 2204 12114 2213
rect 11806 2202 11812 2204
rect 11868 2202 11892 2204
rect 11948 2202 11972 2204
rect 12028 2202 12052 2204
rect 12108 2202 12114 2204
rect 11868 2150 11870 2202
rect 12050 2150 12052 2202
rect 11806 2148 11812 2150
rect 11868 2148 11892 2150
rect 11948 2148 11972 2150
rect 12028 2148 12052 2150
rect 12108 2148 12114 2150
rect 11806 2139 12114 2148
rect 17234 2204 17542 2213
rect 17234 2202 17240 2204
rect 17296 2202 17320 2204
rect 17376 2202 17400 2204
rect 17456 2202 17480 2204
rect 17536 2202 17542 2204
rect 17296 2150 17298 2202
rect 17478 2150 17480 2202
rect 17234 2148 17240 2150
rect 17296 2148 17320 2150
rect 17376 2148 17400 2150
rect 17456 2148 17480 2150
rect 17536 2148 17542 2150
rect 17234 2139 17542 2148
rect 22662 2204 22970 2213
rect 22662 2202 22668 2204
rect 22724 2202 22748 2204
rect 22804 2202 22828 2204
rect 22884 2202 22908 2204
rect 22964 2202 22970 2204
rect 22724 2150 22726 2202
rect 22906 2150 22908 2202
rect 22662 2148 22668 2150
rect 22724 2148 22748 2150
rect 22804 2148 22828 2150
rect 22884 2148 22908 2150
rect 22964 2148 22970 2150
rect 22662 2139 22970 2148
<< via2 >>
rect 6384 21786 6440 21788
rect 6464 21786 6520 21788
rect 6544 21786 6600 21788
rect 6624 21786 6680 21788
rect 6384 21734 6430 21786
rect 6430 21734 6440 21786
rect 6464 21734 6494 21786
rect 6494 21734 6506 21786
rect 6506 21734 6520 21786
rect 6544 21734 6558 21786
rect 6558 21734 6570 21786
rect 6570 21734 6600 21786
rect 6624 21734 6634 21786
rect 6634 21734 6680 21786
rect 6384 21732 6440 21734
rect 6464 21732 6520 21734
rect 6544 21732 6600 21734
rect 6624 21732 6680 21734
rect 11812 21786 11868 21788
rect 11892 21786 11948 21788
rect 11972 21786 12028 21788
rect 12052 21786 12108 21788
rect 11812 21734 11858 21786
rect 11858 21734 11868 21786
rect 11892 21734 11922 21786
rect 11922 21734 11934 21786
rect 11934 21734 11948 21786
rect 11972 21734 11986 21786
rect 11986 21734 11998 21786
rect 11998 21734 12028 21786
rect 12052 21734 12062 21786
rect 12062 21734 12108 21786
rect 11812 21732 11868 21734
rect 11892 21732 11948 21734
rect 11972 21732 12028 21734
rect 12052 21732 12108 21734
rect 17240 21786 17296 21788
rect 17320 21786 17376 21788
rect 17400 21786 17456 21788
rect 17480 21786 17536 21788
rect 17240 21734 17286 21786
rect 17286 21734 17296 21786
rect 17320 21734 17350 21786
rect 17350 21734 17362 21786
rect 17362 21734 17376 21786
rect 17400 21734 17414 21786
rect 17414 21734 17426 21786
rect 17426 21734 17456 21786
rect 17480 21734 17490 21786
rect 17490 21734 17536 21786
rect 17240 21732 17296 21734
rect 17320 21732 17376 21734
rect 17400 21732 17456 21734
rect 17480 21732 17536 21734
rect 22668 21786 22724 21788
rect 22748 21786 22804 21788
rect 22828 21786 22884 21788
rect 22908 21786 22964 21788
rect 22668 21734 22714 21786
rect 22714 21734 22724 21786
rect 22748 21734 22778 21786
rect 22778 21734 22790 21786
rect 22790 21734 22804 21786
rect 22828 21734 22842 21786
rect 22842 21734 22854 21786
rect 22854 21734 22884 21786
rect 22908 21734 22918 21786
rect 22918 21734 22964 21786
rect 22668 21732 22724 21734
rect 22748 21732 22804 21734
rect 22828 21732 22884 21734
rect 22908 21732 22964 21734
rect 3670 21242 3726 21244
rect 3750 21242 3806 21244
rect 3830 21242 3886 21244
rect 3910 21242 3966 21244
rect 3670 21190 3716 21242
rect 3716 21190 3726 21242
rect 3750 21190 3780 21242
rect 3780 21190 3792 21242
rect 3792 21190 3806 21242
rect 3830 21190 3844 21242
rect 3844 21190 3856 21242
rect 3856 21190 3886 21242
rect 3910 21190 3920 21242
rect 3920 21190 3966 21242
rect 3670 21188 3726 21190
rect 3750 21188 3806 21190
rect 3830 21188 3886 21190
rect 3910 21188 3966 21190
rect 9098 21242 9154 21244
rect 9178 21242 9234 21244
rect 9258 21242 9314 21244
rect 9338 21242 9394 21244
rect 9098 21190 9144 21242
rect 9144 21190 9154 21242
rect 9178 21190 9208 21242
rect 9208 21190 9220 21242
rect 9220 21190 9234 21242
rect 9258 21190 9272 21242
rect 9272 21190 9284 21242
rect 9284 21190 9314 21242
rect 9338 21190 9348 21242
rect 9348 21190 9394 21242
rect 9098 21188 9154 21190
rect 9178 21188 9234 21190
rect 9258 21188 9314 21190
rect 9338 21188 9394 21190
rect 14526 21242 14582 21244
rect 14606 21242 14662 21244
rect 14686 21242 14742 21244
rect 14766 21242 14822 21244
rect 14526 21190 14572 21242
rect 14572 21190 14582 21242
rect 14606 21190 14636 21242
rect 14636 21190 14648 21242
rect 14648 21190 14662 21242
rect 14686 21190 14700 21242
rect 14700 21190 14712 21242
rect 14712 21190 14742 21242
rect 14766 21190 14776 21242
rect 14776 21190 14822 21242
rect 14526 21188 14582 21190
rect 14606 21188 14662 21190
rect 14686 21188 14742 21190
rect 14766 21188 14822 21190
rect 19954 21242 20010 21244
rect 20034 21242 20090 21244
rect 20114 21242 20170 21244
rect 20194 21242 20250 21244
rect 19954 21190 20000 21242
rect 20000 21190 20010 21242
rect 20034 21190 20064 21242
rect 20064 21190 20076 21242
rect 20076 21190 20090 21242
rect 20114 21190 20128 21242
rect 20128 21190 20140 21242
rect 20140 21190 20170 21242
rect 20194 21190 20204 21242
rect 20204 21190 20250 21242
rect 19954 21188 20010 21190
rect 20034 21188 20090 21190
rect 20114 21188 20170 21190
rect 20194 21188 20250 21190
rect 6384 20698 6440 20700
rect 6464 20698 6520 20700
rect 6544 20698 6600 20700
rect 6624 20698 6680 20700
rect 6384 20646 6430 20698
rect 6430 20646 6440 20698
rect 6464 20646 6494 20698
rect 6494 20646 6506 20698
rect 6506 20646 6520 20698
rect 6544 20646 6558 20698
rect 6558 20646 6570 20698
rect 6570 20646 6600 20698
rect 6624 20646 6634 20698
rect 6634 20646 6680 20698
rect 6384 20644 6440 20646
rect 6464 20644 6520 20646
rect 6544 20644 6600 20646
rect 6624 20644 6680 20646
rect 11812 20698 11868 20700
rect 11892 20698 11948 20700
rect 11972 20698 12028 20700
rect 12052 20698 12108 20700
rect 11812 20646 11858 20698
rect 11858 20646 11868 20698
rect 11892 20646 11922 20698
rect 11922 20646 11934 20698
rect 11934 20646 11948 20698
rect 11972 20646 11986 20698
rect 11986 20646 11998 20698
rect 11998 20646 12028 20698
rect 12052 20646 12062 20698
rect 12062 20646 12108 20698
rect 11812 20644 11868 20646
rect 11892 20644 11948 20646
rect 11972 20644 12028 20646
rect 12052 20644 12108 20646
rect 17240 20698 17296 20700
rect 17320 20698 17376 20700
rect 17400 20698 17456 20700
rect 17480 20698 17536 20700
rect 17240 20646 17286 20698
rect 17286 20646 17296 20698
rect 17320 20646 17350 20698
rect 17350 20646 17362 20698
rect 17362 20646 17376 20698
rect 17400 20646 17414 20698
rect 17414 20646 17426 20698
rect 17426 20646 17456 20698
rect 17480 20646 17490 20698
rect 17490 20646 17536 20698
rect 17240 20644 17296 20646
rect 17320 20644 17376 20646
rect 17400 20644 17456 20646
rect 17480 20644 17536 20646
rect 22668 20698 22724 20700
rect 22748 20698 22804 20700
rect 22828 20698 22884 20700
rect 22908 20698 22964 20700
rect 22668 20646 22714 20698
rect 22714 20646 22724 20698
rect 22748 20646 22778 20698
rect 22778 20646 22790 20698
rect 22790 20646 22804 20698
rect 22828 20646 22842 20698
rect 22842 20646 22854 20698
rect 22854 20646 22884 20698
rect 22908 20646 22918 20698
rect 22918 20646 22964 20698
rect 22668 20644 22724 20646
rect 22748 20644 22804 20646
rect 22828 20644 22884 20646
rect 22908 20644 22964 20646
rect 3670 20154 3726 20156
rect 3750 20154 3806 20156
rect 3830 20154 3886 20156
rect 3910 20154 3966 20156
rect 3670 20102 3716 20154
rect 3716 20102 3726 20154
rect 3750 20102 3780 20154
rect 3780 20102 3792 20154
rect 3792 20102 3806 20154
rect 3830 20102 3844 20154
rect 3844 20102 3856 20154
rect 3856 20102 3886 20154
rect 3910 20102 3920 20154
rect 3920 20102 3966 20154
rect 3670 20100 3726 20102
rect 3750 20100 3806 20102
rect 3830 20100 3886 20102
rect 3910 20100 3966 20102
rect 9098 20154 9154 20156
rect 9178 20154 9234 20156
rect 9258 20154 9314 20156
rect 9338 20154 9394 20156
rect 9098 20102 9144 20154
rect 9144 20102 9154 20154
rect 9178 20102 9208 20154
rect 9208 20102 9220 20154
rect 9220 20102 9234 20154
rect 9258 20102 9272 20154
rect 9272 20102 9284 20154
rect 9284 20102 9314 20154
rect 9338 20102 9348 20154
rect 9348 20102 9394 20154
rect 9098 20100 9154 20102
rect 9178 20100 9234 20102
rect 9258 20100 9314 20102
rect 9338 20100 9394 20102
rect 14526 20154 14582 20156
rect 14606 20154 14662 20156
rect 14686 20154 14742 20156
rect 14766 20154 14822 20156
rect 14526 20102 14572 20154
rect 14572 20102 14582 20154
rect 14606 20102 14636 20154
rect 14636 20102 14648 20154
rect 14648 20102 14662 20154
rect 14686 20102 14700 20154
rect 14700 20102 14712 20154
rect 14712 20102 14742 20154
rect 14766 20102 14776 20154
rect 14776 20102 14822 20154
rect 14526 20100 14582 20102
rect 14606 20100 14662 20102
rect 14686 20100 14742 20102
rect 14766 20100 14822 20102
rect 19954 20154 20010 20156
rect 20034 20154 20090 20156
rect 20114 20154 20170 20156
rect 20194 20154 20250 20156
rect 19954 20102 20000 20154
rect 20000 20102 20010 20154
rect 20034 20102 20064 20154
rect 20064 20102 20076 20154
rect 20076 20102 20090 20154
rect 20114 20102 20128 20154
rect 20128 20102 20140 20154
rect 20140 20102 20170 20154
rect 20194 20102 20204 20154
rect 20204 20102 20250 20154
rect 19954 20100 20010 20102
rect 20034 20100 20090 20102
rect 20114 20100 20170 20102
rect 20194 20100 20250 20102
rect 2134 19760 2190 19816
rect 6384 19610 6440 19612
rect 6464 19610 6520 19612
rect 6544 19610 6600 19612
rect 6624 19610 6680 19612
rect 6384 19558 6430 19610
rect 6430 19558 6440 19610
rect 6464 19558 6494 19610
rect 6494 19558 6506 19610
rect 6506 19558 6520 19610
rect 6544 19558 6558 19610
rect 6558 19558 6570 19610
rect 6570 19558 6600 19610
rect 6624 19558 6634 19610
rect 6634 19558 6680 19610
rect 6384 19556 6440 19558
rect 6464 19556 6520 19558
rect 6544 19556 6600 19558
rect 6624 19556 6680 19558
rect 11812 19610 11868 19612
rect 11892 19610 11948 19612
rect 11972 19610 12028 19612
rect 12052 19610 12108 19612
rect 11812 19558 11858 19610
rect 11858 19558 11868 19610
rect 11892 19558 11922 19610
rect 11922 19558 11934 19610
rect 11934 19558 11948 19610
rect 11972 19558 11986 19610
rect 11986 19558 11998 19610
rect 11998 19558 12028 19610
rect 12052 19558 12062 19610
rect 12062 19558 12108 19610
rect 11812 19556 11868 19558
rect 11892 19556 11948 19558
rect 11972 19556 12028 19558
rect 12052 19556 12108 19558
rect 17240 19610 17296 19612
rect 17320 19610 17376 19612
rect 17400 19610 17456 19612
rect 17480 19610 17536 19612
rect 17240 19558 17286 19610
rect 17286 19558 17296 19610
rect 17320 19558 17350 19610
rect 17350 19558 17362 19610
rect 17362 19558 17376 19610
rect 17400 19558 17414 19610
rect 17414 19558 17426 19610
rect 17426 19558 17456 19610
rect 17480 19558 17490 19610
rect 17490 19558 17536 19610
rect 17240 19556 17296 19558
rect 17320 19556 17376 19558
rect 17400 19556 17456 19558
rect 17480 19556 17536 19558
rect 22668 19610 22724 19612
rect 22748 19610 22804 19612
rect 22828 19610 22884 19612
rect 22908 19610 22964 19612
rect 22668 19558 22714 19610
rect 22714 19558 22724 19610
rect 22748 19558 22778 19610
rect 22778 19558 22790 19610
rect 22790 19558 22804 19610
rect 22828 19558 22842 19610
rect 22842 19558 22854 19610
rect 22854 19558 22884 19610
rect 22908 19558 22918 19610
rect 22918 19558 22964 19610
rect 22668 19556 22724 19558
rect 22748 19556 22804 19558
rect 22828 19556 22884 19558
rect 22908 19556 22964 19558
rect 3670 19066 3726 19068
rect 3750 19066 3806 19068
rect 3830 19066 3886 19068
rect 3910 19066 3966 19068
rect 3670 19014 3716 19066
rect 3716 19014 3726 19066
rect 3750 19014 3780 19066
rect 3780 19014 3792 19066
rect 3792 19014 3806 19066
rect 3830 19014 3844 19066
rect 3844 19014 3856 19066
rect 3856 19014 3886 19066
rect 3910 19014 3920 19066
rect 3920 19014 3966 19066
rect 3670 19012 3726 19014
rect 3750 19012 3806 19014
rect 3830 19012 3886 19014
rect 3910 19012 3966 19014
rect 9098 19066 9154 19068
rect 9178 19066 9234 19068
rect 9258 19066 9314 19068
rect 9338 19066 9394 19068
rect 9098 19014 9144 19066
rect 9144 19014 9154 19066
rect 9178 19014 9208 19066
rect 9208 19014 9220 19066
rect 9220 19014 9234 19066
rect 9258 19014 9272 19066
rect 9272 19014 9284 19066
rect 9284 19014 9314 19066
rect 9338 19014 9348 19066
rect 9348 19014 9394 19066
rect 9098 19012 9154 19014
rect 9178 19012 9234 19014
rect 9258 19012 9314 19014
rect 9338 19012 9394 19014
rect 14526 19066 14582 19068
rect 14606 19066 14662 19068
rect 14686 19066 14742 19068
rect 14766 19066 14822 19068
rect 14526 19014 14572 19066
rect 14572 19014 14582 19066
rect 14606 19014 14636 19066
rect 14636 19014 14648 19066
rect 14648 19014 14662 19066
rect 14686 19014 14700 19066
rect 14700 19014 14712 19066
rect 14712 19014 14742 19066
rect 14766 19014 14776 19066
rect 14776 19014 14822 19066
rect 14526 19012 14582 19014
rect 14606 19012 14662 19014
rect 14686 19012 14742 19014
rect 14766 19012 14822 19014
rect 19954 19066 20010 19068
rect 20034 19066 20090 19068
rect 20114 19066 20170 19068
rect 20194 19066 20250 19068
rect 19954 19014 20000 19066
rect 20000 19014 20010 19066
rect 20034 19014 20064 19066
rect 20064 19014 20076 19066
rect 20076 19014 20090 19066
rect 20114 19014 20128 19066
rect 20128 19014 20140 19066
rect 20140 19014 20170 19066
rect 20194 19014 20204 19066
rect 20204 19014 20250 19066
rect 19954 19012 20010 19014
rect 20034 19012 20090 19014
rect 20114 19012 20170 19014
rect 20194 19012 20250 19014
rect 6384 18522 6440 18524
rect 6464 18522 6520 18524
rect 6544 18522 6600 18524
rect 6624 18522 6680 18524
rect 6384 18470 6430 18522
rect 6430 18470 6440 18522
rect 6464 18470 6494 18522
rect 6494 18470 6506 18522
rect 6506 18470 6520 18522
rect 6544 18470 6558 18522
rect 6558 18470 6570 18522
rect 6570 18470 6600 18522
rect 6624 18470 6634 18522
rect 6634 18470 6680 18522
rect 6384 18468 6440 18470
rect 6464 18468 6520 18470
rect 6544 18468 6600 18470
rect 6624 18468 6680 18470
rect 11812 18522 11868 18524
rect 11892 18522 11948 18524
rect 11972 18522 12028 18524
rect 12052 18522 12108 18524
rect 11812 18470 11858 18522
rect 11858 18470 11868 18522
rect 11892 18470 11922 18522
rect 11922 18470 11934 18522
rect 11934 18470 11948 18522
rect 11972 18470 11986 18522
rect 11986 18470 11998 18522
rect 11998 18470 12028 18522
rect 12052 18470 12062 18522
rect 12062 18470 12108 18522
rect 11812 18468 11868 18470
rect 11892 18468 11948 18470
rect 11972 18468 12028 18470
rect 12052 18468 12108 18470
rect 17240 18522 17296 18524
rect 17320 18522 17376 18524
rect 17400 18522 17456 18524
rect 17480 18522 17536 18524
rect 17240 18470 17286 18522
rect 17286 18470 17296 18522
rect 17320 18470 17350 18522
rect 17350 18470 17362 18522
rect 17362 18470 17376 18522
rect 17400 18470 17414 18522
rect 17414 18470 17426 18522
rect 17426 18470 17456 18522
rect 17480 18470 17490 18522
rect 17490 18470 17536 18522
rect 17240 18468 17296 18470
rect 17320 18468 17376 18470
rect 17400 18468 17456 18470
rect 17480 18468 17536 18470
rect 22668 18522 22724 18524
rect 22748 18522 22804 18524
rect 22828 18522 22884 18524
rect 22908 18522 22964 18524
rect 22668 18470 22714 18522
rect 22714 18470 22724 18522
rect 22748 18470 22778 18522
rect 22778 18470 22790 18522
rect 22790 18470 22804 18522
rect 22828 18470 22842 18522
rect 22842 18470 22854 18522
rect 22854 18470 22884 18522
rect 22908 18470 22918 18522
rect 22918 18470 22964 18522
rect 22668 18468 22724 18470
rect 22748 18468 22804 18470
rect 22828 18468 22884 18470
rect 22908 18468 22964 18470
rect 3670 17978 3726 17980
rect 3750 17978 3806 17980
rect 3830 17978 3886 17980
rect 3910 17978 3966 17980
rect 3670 17926 3716 17978
rect 3716 17926 3726 17978
rect 3750 17926 3780 17978
rect 3780 17926 3792 17978
rect 3792 17926 3806 17978
rect 3830 17926 3844 17978
rect 3844 17926 3856 17978
rect 3856 17926 3886 17978
rect 3910 17926 3920 17978
rect 3920 17926 3966 17978
rect 3670 17924 3726 17926
rect 3750 17924 3806 17926
rect 3830 17924 3886 17926
rect 3910 17924 3966 17926
rect 9098 17978 9154 17980
rect 9178 17978 9234 17980
rect 9258 17978 9314 17980
rect 9338 17978 9394 17980
rect 9098 17926 9144 17978
rect 9144 17926 9154 17978
rect 9178 17926 9208 17978
rect 9208 17926 9220 17978
rect 9220 17926 9234 17978
rect 9258 17926 9272 17978
rect 9272 17926 9284 17978
rect 9284 17926 9314 17978
rect 9338 17926 9348 17978
rect 9348 17926 9394 17978
rect 9098 17924 9154 17926
rect 9178 17924 9234 17926
rect 9258 17924 9314 17926
rect 9338 17924 9394 17926
rect 14526 17978 14582 17980
rect 14606 17978 14662 17980
rect 14686 17978 14742 17980
rect 14766 17978 14822 17980
rect 14526 17926 14572 17978
rect 14572 17926 14582 17978
rect 14606 17926 14636 17978
rect 14636 17926 14648 17978
rect 14648 17926 14662 17978
rect 14686 17926 14700 17978
rect 14700 17926 14712 17978
rect 14712 17926 14742 17978
rect 14766 17926 14776 17978
rect 14776 17926 14822 17978
rect 14526 17924 14582 17926
rect 14606 17924 14662 17926
rect 14686 17924 14742 17926
rect 14766 17924 14822 17926
rect 19954 17978 20010 17980
rect 20034 17978 20090 17980
rect 20114 17978 20170 17980
rect 20194 17978 20250 17980
rect 19954 17926 20000 17978
rect 20000 17926 20010 17978
rect 20034 17926 20064 17978
rect 20064 17926 20076 17978
rect 20076 17926 20090 17978
rect 20114 17926 20128 17978
rect 20128 17926 20140 17978
rect 20140 17926 20170 17978
rect 20194 17926 20204 17978
rect 20204 17926 20250 17978
rect 19954 17924 20010 17926
rect 20034 17924 20090 17926
rect 20114 17924 20170 17926
rect 20194 17924 20250 17926
rect 6384 17434 6440 17436
rect 6464 17434 6520 17436
rect 6544 17434 6600 17436
rect 6624 17434 6680 17436
rect 6384 17382 6430 17434
rect 6430 17382 6440 17434
rect 6464 17382 6494 17434
rect 6494 17382 6506 17434
rect 6506 17382 6520 17434
rect 6544 17382 6558 17434
rect 6558 17382 6570 17434
rect 6570 17382 6600 17434
rect 6624 17382 6634 17434
rect 6634 17382 6680 17434
rect 6384 17380 6440 17382
rect 6464 17380 6520 17382
rect 6544 17380 6600 17382
rect 6624 17380 6680 17382
rect 11812 17434 11868 17436
rect 11892 17434 11948 17436
rect 11972 17434 12028 17436
rect 12052 17434 12108 17436
rect 11812 17382 11858 17434
rect 11858 17382 11868 17434
rect 11892 17382 11922 17434
rect 11922 17382 11934 17434
rect 11934 17382 11948 17434
rect 11972 17382 11986 17434
rect 11986 17382 11998 17434
rect 11998 17382 12028 17434
rect 12052 17382 12062 17434
rect 12062 17382 12108 17434
rect 11812 17380 11868 17382
rect 11892 17380 11948 17382
rect 11972 17380 12028 17382
rect 12052 17380 12108 17382
rect 17240 17434 17296 17436
rect 17320 17434 17376 17436
rect 17400 17434 17456 17436
rect 17480 17434 17536 17436
rect 17240 17382 17286 17434
rect 17286 17382 17296 17434
rect 17320 17382 17350 17434
rect 17350 17382 17362 17434
rect 17362 17382 17376 17434
rect 17400 17382 17414 17434
rect 17414 17382 17426 17434
rect 17426 17382 17456 17434
rect 17480 17382 17490 17434
rect 17490 17382 17536 17434
rect 17240 17380 17296 17382
rect 17320 17380 17376 17382
rect 17400 17380 17456 17382
rect 17480 17380 17536 17382
rect 22668 17434 22724 17436
rect 22748 17434 22804 17436
rect 22828 17434 22884 17436
rect 22908 17434 22964 17436
rect 22668 17382 22714 17434
rect 22714 17382 22724 17434
rect 22748 17382 22778 17434
rect 22778 17382 22790 17434
rect 22790 17382 22804 17434
rect 22828 17382 22842 17434
rect 22842 17382 22854 17434
rect 22854 17382 22884 17434
rect 22908 17382 22918 17434
rect 22918 17382 22964 17434
rect 22668 17380 22724 17382
rect 22748 17380 22804 17382
rect 22828 17380 22884 17382
rect 22908 17380 22964 17382
rect 3670 16890 3726 16892
rect 3750 16890 3806 16892
rect 3830 16890 3886 16892
rect 3910 16890 3966 16892
rect 3670 16838 3716 16890
rect 3716 16838 3726 16890
rect 3750 16838 3780 16890
rect 3780 16838 3792 16890
rect 3792 16838 3806 16890
rect 3830 16838 3844 16890
rect 3844 16838 3856 16890
rect 3856 16838 3886 16890
rect 3910 16838 3920 16890
rect 3920 16838 3966 16890
rect 3670 16836 3726 16838
rect 3750 16836 3806 16838
rect 3830 16836 3886 16838
rect 3910 16836 3966 16838
rect 9098 16890 9154 16892
rect 9178 16890 9234 16892
rect 9258 16890 9314 16892
rect 9338 16890 9394 16892
rect 9098 16838 9144 16890
rect 9144 16838 9154 16890
rect 9178 16838 9208 16890
rect 9208 16838 9220 16890
rect 9220 16838 9234 16890
rect 9258 16838 9272 16890
rect 9272 16838 9284 16890
rect 9284 16838 9314 16890
rect 9338 16838 9348 16890
rect 9348 16838 9394 16890
rect 9098 16836 9154 16838
rect 9178 16836 9234 16838
rect 9258 16836 9314 16838
rect 9338 16836 9394 16838
rect 14526 16890 14582 16892
rect 14606 16890 14662 16892
rect 14686 16890 14742 16892
rect 14766 16890 14822 16892
rect 14526 16838 14572 16890
rect 14572 16838 14582 16890
rect 14606 16838 14636 16890
rect 14636 16838 14648 16890
rect 14648 16838 14662 16890
rect 14686 16838 14700 16890
rect 14700 16838 14712 16890
rect 14712 16838 14742 16890
rect 14766 16838 14776 16890
rect 14776 16838 14822 16890
rect 14526 16836 14582 16838
rect 14606 16836 14662 16838
rect 14686 16836 14742 16838
rect 14766 16836 14822 16838
rect 19954 16890 20010 16892
rect 20034 16890 20090 16892
rect 20114 16890 20170 16892
rect 20194 16890 20250 16892
rect 19954 16838 20000 16890
rect 20000 16838 20010 16890
rect 20034 16838 20064 16890
rect 20064 16838 20076 16890
rect 20076 16838 20090 16890
rect 20114 16838 20128 16890
rect 20128 16838 20140 16890
rect 20140 16838 20170 16890
rect 20194 16838 20204 16890
rect 20204 16838 20250 16890
rect 19954 16836 20010 16838
rect 20034 16836 20090 16838
rect 20114 16836 20170 16838
rect 20194 16836 20250 16838
rect 6384 16346 6440 16348
rect 6464 16346 6520 16348
rect 6544 16346 6600 16348
rect 6624 16346 6680 16348
rect 6384 16294 6430 16346
rect 6430 16294 6440 16346
rect 6464 16294 6494 16346
rect 6494 16294 6506 16346
rect 6506 16294 6520 16346
rect 6544 16294 6558 16346
rect 6558 16294 6570 16346
rect 6570 16294 6600 16346
rect 6624 16294 6634 16346
rect 6634 16294 6680 16346
rect 6384 16292 6440 16294
rect 6464 16292 6520 16294
rect 6544 16292 6600 16294
rect 6624 16292 6680 16294
rect 11812 16346 11868 16348
rect 11892 16346 11948 16348
rect 11972 16346 12028 16348
rect 12052 16346 12108 16348
rect 11812 16294 11858 16346
rect 11858 16294 11868 16346
rect 11892 16294 11922 16346
rect 11922 16294 11934 16346
rect 11934 16294 11948 16346
rect 11972 16294 11986 16346
rect 11986 16294 11998 16346
rect 11998 16294 12028 16346
rect 12052 16294 12062 16346
rect 12062 16294 12108 16346
rect 11812 16292 11868 16294
rect 11892 16292 11948 16294
rect 11972 16292 12028 16294
rect 12052 16292 12108 16294
rect 17240 16346 17296 16348
rect 17320 16346 17376 16348
rect 17400 16346 17456 16348
rect 17480 16346 17536 16348
rect 17240 16294 17286 16346
rect 17286 16294 17296 16346
rect 17320 16294 17350 16346
rect 17350 16294 17362 16346
rect 17362 16294 17376 16346
rect 17400 16294 17414 16346
rect 17414 16294 17426 16346
rect 17426 16294 17456 16346
rect 17480 16294 17490 16346
rect 17490 16294 17536 16346
rect 17240 16292 17296 16294
rect 17320 16292 17376 16294
rect 17400 16292 17456 16294
rect 17480 16292 17536 16294
rect 22668 16346 22724 16348
rect 22748 16346 22804 16348
rect 22828 16346 22884 16348
rect 22908 16346 22964 16348
rect 22668 16294 22714 16346
rect 22714 16294 22724 16346
rect 22748 16294 22778 16346
rect 22778 16294 22790 16346
rect 22790 16294 22804 16346
rect 22828 16294 22842 16346
rect 22842 16294 22854 16346
rect 22854 16294 22884 16346
rect 22908 16294 22918 16346
rect 22918 16294 22964 16346
rect 22668 16292 22724 16294
rect 22748 16292 22804 16294
rect 22828 16292 22884 16294
rect 22908 16292 22964 16294
rect 3670 15802 3726 15804
rect 3750 15802 3806 15804
rect 3830 15802 3886 15804
rect 3910 15802 3966 15804
rect 3670 15750 3716 15802
rect 3716 15750 3726 15802
rect 3750 15750 3780 15802
rect 3780 15750 3792 15802
rect 3792 15750 3806 15802
rect 3830 15750 3844 15802
rect 3844 15750 3856 15802
rect 3856 15750 3886 15802
rect 3910 15750 3920 15802
rect 3920 15750 3966 15802
rect 3670 15748 3726 15750
rect 3750 15748 3806 15750
rect 3830 15748 3886 15750
rect 3910 15748 3966 15750
rect 3514 14900 3516 14920
rect 3516 14900 3568 14920
rect 3568 14900 3570 14920
rect 3514 14864 3570 14900
rect 3670 14714 3726 14716
rect 3750 14714 3806 14716
rect 3830 14714 3886 14716
rect 3910 14714 3966 14716
rect 3670 14662 3716 14714
rect 3716 14662 3726 14714
rect 3750 14662 3780 14714
rect 3780 14662 3792 14714
rect 3792 14662 3806 14714
rect 3830 14662 3844 14714
rect 3844 14662 3856 14714
rect 3856 14662 3886 14714
rect 3910 14662 3920 14714
rect 3920 14662 3966 14714
rect 3670 14660 3726 14662
rect 3750 14660 3806 14662
rect 3830 14660 3886 14662
rect 3910 14660 3966 14662
rect 2778 11872 2834 11928
rect 3670 13626 3726 13628
rect 3750 13626 3806 13628
rect 3830 13626 3886 13628
rect 3910 13626 3966 13628
rect 3670 13574 3716 13626
rect 3716 13574 3726 13626
rect 3750 13574 3780 13626
rect 3780 13574 3792 13626
rect 3792 13574 3806 13626
rect 3830 13574 3844 13626
rect 3844 13574 3856 13626
rect 3856 13574 3886 13626
rect 3910 13574 3920 13626
rect 3920 13574 3966 13626
rect 3670 13572 3726 13574
rect 3750 13572 3806 13574
rect 3830 13572 3886 13574
rect 3910 13572 3966 13574
rect 3670 12538 3726 12540
rect 3750 12538 3806 12540
rect 3830 12538 3886 12540
rect 3910 12538 3966 12540
rect 3670 12486 3716 12538
rect 3716 12486 3726 12538
rect 3750 12486 3780 12538
rect 3780 12486 3792 12538
rect 3792 12486 3806 12538
rect 3830 12486 3844 12538
rect 3844 12486 3856 12538
rect 3856 12486 3886 12538
rect 3910 12486 3920 12538
rect 3920 12486 3966 12538
rect 3670 12484 3726 12486
rect 3750 12484 3806 12486
rect 3830 12484 3886 12486
rect 3910 12484 3966 12486
rect 3670 11450 3726 11452
rect 3750 11450 3806 11452
rect 3830 11450 3886 11452
rect 3910 11450 3966 11452
rect 3670 11398 3716 11450
rect 3716 11398 3726 11450
rect 3750 11398 3780 11450
rect 3780 11398 3792 11450
rect 3792 11398 3806 11450
rect 3830 11398 3844 11450
rect 3844 11398 3856 11450
rect 3856 11398 3886 11450
rect 3910 11398 3920 11450
rect 3920 11398 3966 11450
rect 3670 11396 3726 11398
rect 3750 11396 3806 11398
rect 3830 11396 3886 11398
rect 3910 11396 3966 11398
rect 6384 15258 6440 15260
rect 6464 15258 6520 15260
rect 6544 15258 6600 15260
rect 6624 15258 6680 15260
rect 6384 15206 6430 15258
rect 6430 15206 6440 15258
rect 6464 15206 6494 15258
rect 6494 15206 6506 15258
rect 6506 15206 6520 15258
rect 6544 15206 6558 15258
rect 6558 15206 6570 15258
rect 6570 15206 6600 15258
rect 6624 15206 6634 15258
rect 6634 15206 6680 15258
rect 6384 15204 6440 15206
rect 6464 15204 6520 15206
rect 6544 15204 6600 15206
rect 6624 15204 6680 15206
rect 3670 10362 3726 10364
rect 3750 10362 3806 10364
rect 3830 10362 3886 10364
rect 3910 10362 3966 10364
rect 3670 10310 3716 10362
rect 3716 10310 3726 10362
rect 3750 10310 3780 10362
rect 3780 10310 3792 10362
rect 3792 10310 3806 10362
rect 3830 10310 3844 10362
rect 3844 10310 3856 10362
rect 3856 10310 3886 10362
rect 3910 10310 3920 10362
rect 3920 10310 3966 10362
rect 3670 10308 3726 10310
rect 3750 10308 3806 10310
rect 3830 10308 3886 10310
rect 3910 10308 3966 10310
rect 3670 9274 3726 9276
rect 3750 9274 3806 9276
rect 3830 9274 3886 9276
rect 3910 9274 3966 9276
rect 3670 9222 3716 9274
rect 3716 9222 3726 9274
rect 3750 9222 3780 9274
rect 3780 9222 3792 9274
rect 3792 9222 3806 9274
rect 3830 9222 3844 9274
rect 3844 9222 3856 9274
rect 3856 9222 3886 9274
rect 3910 9222 3920 9274
rect 3920 9222 3966 9274
rect 3670 9220 3726 9222
rect 3750 9220 3806 9222
rect 3830 9220 3886 9222
rect 3910 9220 3966 9222
rect 9098 15802 9154 15804
rect 9178 15802 9234 15804
rect 9258 15802 9314 15804
rect 9338 15802 9394 15804
rect 9098 15750 9144 15802
rect 9144 15750 9154 15802
rect 9178 15750 9208 15802
rect 9208 15750 9220 15802
rect 9220 15750 9234 15802
rect 9258 15750 9272 15802
rect 9272 15750 9284 15802
rect 9284 15750 9314 15802
rect 9338 15750 9348 15802
rect 9348 15750 9394 15802
rect 9098 15748 9154 15750
rect 9178 15748 9234 15750
rect 9258 15748 9314 15750
rect 9338 15748 9394 15750
rect 14526 15802 14582 15804
rect 14606 15802 14662 15804
rect 14686 15802 14742 15804
rect 14766 15802 14822 15804
rect 14526 15750 14572 15802
rect 14572 15750 14582 15802
rect 14606 15750 14636 15802
rect 14636 15750 14648 15802
rect 14648 15750 14662 15802
rect 14686 15750 14700 15802
rect 14700 15750 14712 15802
rect 14712 15750 14742 15802
rect 14766 15750 14776 15802
rect 14776 15750 14822 15802
rect 14526 15748 14582 15750
rect 14606 15748 14662 15750
rect 14686 15748 14742 15750
rect 14766 15748 14822 15750
rect 19954 15802 20010 15804
rect 20034 15802 20090 15804
rect 20114 15802 20170 15804
rect 20194 15802 20250 15804
rect 19954 15750 20000 15802
rect 20000 15750 20010 15802
rect 20034 15750 20064 15802
rect 20064 15750 20076 15802
rect 20076 15750 20090 15802
rect 20114 15750 20128 15802
rect 20128 15750 20140 15802
rect 20140 15750 20170 15802
rect 20194 15750 20204 15802
rect 20204 15750 20250 15802
rect 19954 15748 20010 15750
rect 20034 15748 20090 15750
rect 20114 15748 20170 15750
rect 20194 15748 20250 15750
rect 6384 14170 6440 14172
rect 6464 14170 6520 14172
rect 6544 14170 6600 14172
rect 6624 14170 6680 14172
rect 6384 14118 6430 14170
rect 6430 14118 6440 14170
rect 6464 14118 6494 14170
rect 6494 14118 6506 14170
rect 6506 14118 6520 14170
rect 6544 14118 6558 14170
rect 6558 14118 6570 14170
rect 6570 14118 6600 14170
rect 6624 14118 6634 14170
rect 6634 14118 6680 14170
rect 6384 14116 6440 14118
rect 6464 14116 6520 14118
rect 6544 14116 6600 14118
rect 6624 14116 6680 14118
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6430 13082
rect 6430 13030 6440 13082
rect 6464 13030 6494 13082
rect 6494 13030 6506 13082
rect 6506 13030 6520 13082
rect 6544 13030 6558 13082
rect 6558 13030 6570 13082
rect 6570 13030 6600 13082
rect 6624 13030 6634 13082
rect 6634 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 3670 8186 3726 8188
rect 3750 8186 3806 8188
rect 3830 8186 3886 8188
rect 3910 8186 3966 8188
rect 3670 8134 3716 8186
rect 3716 8134 3726 8186
rect 3750 8134 3780 8186
rect 3780 8134 3792 8186
rect 3792 8134 3806 8186
rect 3830 8134 3844 8186
rect 3844 8134 3856 8186
rect 3856 8134 3886 8186
rect 3910 8134 3920 8186
rect 3920 8134 3966 8186
rect 3670 8132 3726 8134
rect 3750 8132 3806 8134
rect 3830 8132 3886 8134
rect 3910 8132 3966 8134
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6430 11994
rect 6430 11942 6440 11994
rect 6464 11942 6494 11994
rect 6494 11942 6506 11994
rect 6506 11942 6520 11994
rect 6544 11942 6558 11994
rect 6558 11942 6570 11994
rect 6570 11942 6600 11994
rect 6624 11942 6634 11994
rect 6634 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6430 10906
rect 6430 10854 6440 10906
rect 6464 10854 6494 10906
rect 6494 10854 6506 10906
rect 6506 10854 6520 10906
rect 6544 10854 6558 10906
rect 6558 10854 6570 10906
rect 6570 10854 6600 10906
rect 6624 10854 6634 10906
rect 6634 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6430 9818
rect 6430 9766 6440 9818
rect 6464 9766 6494 9818
rect 6494 9766 6506 9818
rect 6506 9766 6520 9818
rect 6544 9766 6558 9818
rect 6558 9766 6570 9818
rect 6570 9766 6600 9818
rect 6624 9766 6634 9818
rect 6634 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6430 8730
rect 6430 8678 6440 8730
rect 6464 8678 6494 8730
rect 6494 8678 6506 8730
rect 6506 8678 6520 8730
rect 6544 8678 6558 8730
rect 6558 8678 6570 8730
rect 6570 8678 6600 8730
rect 6624 8678 6634 8730
rect 6634 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6430 7642
rect 6430 7590 6440 7642
rect 6464 7590 6494 7642
rect 6494 7590 6506 7642
rect 6506 7590 6520 7642
rect 6544 7590 6558 7642
rect 6558 7590 6570 7642
rect 6570 7590 6600 7642
rect 6624 7590 6634 7642
rect 6634 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 4066 3984 4122 4040
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6430 6554
rect 6430 6502 6440 6554
rect 6464 6502 6494 6554
rect 6494 6502 6506 6554
rect 6506 6502 6520 6554
rect 6544 6502 6558 6554
rect 6558 6502 6570 6554
rect 6570 6502 6600 6554
rect 6624 6502 6634 6554
rect 6634 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6430 5466
rect 6430 5414 6440 5466
rect 6464 5414 6494 5466
rect 6494 5414 6506 5466
rect 6506 5414 6520 5466
rect 6544 5414 6558 5466
rect 6558 5414 6570 5466
rect 6570 5414 6600 5466
rect 6624 5414 6634 5466
rect 6634 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6430 4378
rect 6430 4326 6440 4378
rect 6464 4326 6494 4378
rect 6494 4326 6506 4378
rect 6506 4326 6520 4378
rect 6544 4326 6558 4378
rect 6558 4326 6570 4378
rect 6570 4326 6600 4378
rect 6624 4326 6634 4378
rect 6634 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6430 3290
rect 6430 3238 6440 3290
rect 6464 3238 6494 3290
rect 6494 3238 6506 3290
rect 6506 3238 6520 3290
rect 6544 3238 6558 3290
rect 6558 3238 6570 3290
rect 6570 3238 6600 3290
rect 6624 3238 6634 3290
rect 6634 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 8942 14884 8998 14920
rect 8942 14864 8944 14884
rect 8944 14864 8996 14884
rect 8996 14864 8998 14884
rect 11812 15258 11868 15260
rect 11892 15258 11948 15260
rect 11972 15258 12028 15260
rect 12052 15258 12108 15260
rect 11812 15206 11858 15258
rect 11858 15206 11868 15258
rect 11892 15206 11922 15258
rect 11922 15206 11934 15258
rect 11934 15206 11948 15258
rect 11972 15206 11986 15258
rect 11986 15206 11998 15258
rect 11998 15206 12028 15258
rect 12052 15206 12062 15258
rect 12062 15206 12108 15258
rect 11812 15204 11868 15206
rect 11892 15204 11948 15206
rect 11972 15204 12028 15206
rect 12052 15204 12108 15206
rect 17240 15258 17296 15260
rect 17320 15258 17376 15260
rect 17400 15258 17456 15260
rect 17480 15258 17536 15260
rect 17240 15206 17286 15258
rect 17286 15206 17296 15258
rect 17320 15206 17350 15258
rect 17350 15206 17362 15258
rect 17362 15206 17376 15258
rect 17400 15206 17414 15258
rect 17414 15206 17426 15258
rect 17426 15206 17456 15258
rect 17480 15206 17490 15258
rect 17490 15206 17536 15258
rect 17240 15204 17296 15206
rect 17320 15204 17376 15206
rect 17400 15204 17456 15206
rect 17480 15204 17536 15206
rect 22668 15258 22724 15260
rect 22748 15258 22804 15260
rect 22828 15258 22884 15260
rect 22908 15258 22964 15260
rect 22668 15206 22714 15258
rect 22714 15206 22724 15258
rect 22748 15206 22778 15258
rect 22778 15206 22790 15258
rect 22790 15206 22804 15258
rect 22828 15206 22842 15258
rect 22842 15206 22854 15258
rect 22854 15206 22884 15258
rect 22908 15206 22918 15258
rect 22918 15206 22964 15258
rect 22668 15204 22724 15206
rect 22748 15204 22804 15206
rect 22828 15204 22884 15206
rect 22908 15204 22964 15206
rect 9098 14714 9154 14716
rect 9178 14714 9234 14716
rect 9258 14714 9314 14716
rect 9338 14714 9394 14716
rect 9098 14662 9144 14714
rect 9144 14662 9154 14714
rect 9178 14662 9208 14714
rect 9208 14662 9220 14714
rect 9220 14662 9234 14714
rect 9258 14662 9272 14714
rect 9272 14662 9284 14714
rect 9284 14662 9314 14714
rect 9338 14662 9348 14714
rect 9348 14662 9394 14714
rect 9098 14660 9154 14662
rect 9178 14660 9234 14662
rect 9258 14660 9314 14662
rect 9338 14660 9394 14662
rect 14526 14714 14582 14716
rect 14606 14714 14662 14716
rect 14686 14714 14742 14716
rect 14766 14714 14822 14716
rect 14526 14662 14572 14714
rect 14572 14662 14582 14714
rect 14606 14662 14636 14714
rect 14636 14662 14648 14714
rect 14648 14662 14662 14714
rect 14686 14662 14700 14714
rect 14700 14662 14712 14714
rect 14712 14662 14742 14714
rect 14766 14662 14776 14714
rect 14776 14662 14822 14714
rect 14526 14660 14582 14662
rect 14606 14660 14662 14662
rect 14686 14660 14742 14662
rect 14766 14660 14822 14662
rect 19954 14714 20010 14716
rect 20034 14714 20090 14716
rect 20114 14714 20170 14716
rect 20194 14714 20250 14716
rect 19954 14662 20000 14714
rect 20000 14662 20010 14714
rect 20034 14662 20064 14714
rect 20064 14662 20076 14714
rect 20076 14662 20090 14714
rect 20114 14662 20128 14714
rect 20128 14662 20140 14714
rect 20140 14662 20170 14714
rect 20194 14662 20204 14714
rect 20204 14662 20250 14714
rect 19954 14660 20010 14662
rect 20034 14660 20090 14662
rect 20114 14660 20170 14662
rect 20194 14660 20250 14662
rect 11812 14170 11868 14172
rect 11892 14170 11948 14172
rect 11972 14170 12028 14172
rect 12052 14170 12108 14172
rect 11812 14118 11858 14170
rect 11858 14118 11868 14170
rect 11892 14118 11922 14170
rect 11922 14118 11934 14170
rect 11934 14118 11948 14170
rect 11972 14118 11986 14170
rect 11986 14118 11998 14170
rect 11998 14118 12028 14170
rect 12052 14118 12062 14170
rect 12062 14118 12108 14170
rect 11812 14116 11868 14118
rect 11892 14116 11948 14118
rect 11972 14116 12028 14118
rect 12052 14116 12108 14118
rect 17240 14170 17296 14172
rect 17320 14170 17376 14172
rect 17400 14170 17456 14172
rect 17480 14170 17536 14172
rect 17240 14118 17286 14170
rect 17286 14118 17296 14170
rect 17320 14118 17350 14170
rect 17350 14118 17362 14170
rect 17362 14118 17376 14170
rect 17400 14118 17414 14170
rect 17414 14118 17426 14170
rect 17426 14118 17456 14170
rect 17480 14118 17490 14170
rect 17490 14118 17536 14170
rect 17240 14116 17296 14118
rect 17320 14116 17376 14118
rect 17400 14116 17456 14118
rect 17480 14116 17536 14118
rect 22668 14170 22724 14172
rect 22748 14170 22804 14172
rect 22828 14170 22884 14172
rect 22908 14170 22964 14172
rect 22668 14118 22714 14170
rect 22714 14118 22724 14170
rect 22748 14118 22778 14170
rect 22778 14118 22790 14170
rect 22790 14118 22804 14170
rect 22828 14118 22842 14170
rect 22842 14118 22854 14170
rect 22854 14118 22884 14170
rect 22908 14118 22918 14170
rect 22918 14118 22964 14170
rect 22668 14116 22724 14118
rect 22748 14116 22804 14118
rect 22828 14116 22884 14118
rect 22908 14116 22964 14118
rect 9098 13626 9154 13628
rect 9178 13626 9234 13628
rect 9258 13626 9314 13628
rect 9338 13626 9394 13628
rect 9098 13574 9144 13626
rect 9144 13574 9154 13626
rect 9178 13574 9208 13626
rect 9208 13574 9220 13626
rect 9220 13574 9234 13626
rect 9258 13574 9272 13626
rect 9272 13574 9284 13626
rect 9284 13574 9314 13626
rect 9338 13574 9348 13626
rect 9348 13574 9394 13626
rect 9098 13572 9154 13574
rect 9178 13572 9234 13574
rect 9258 13572 9314 13574
rect 9338 13572 9394 13574
rect 9098 12538 9154 12540
rect 9178 12538 9234 12540
rect 9258 12538 9314 12540
rect 9338 12538 9394 12540
rect 9098 12486 9144 12538
rect 9144 12486 9154 12538
rect 9178 12486 9208 12538
rect 9208 12486 9220 12538
rect 9220 12486 9234 12538
rect 9258 12486 9272 12538
rect 9272 12486 9284 12538
rect 9284 12486 9314 12538
rect 9338 12486 9348 12538
rect 9348 12486 9394 12538
rect 9098 12484 9154 12486
rect 9178 12484 9234 12486
rect 9258 12484 9314 12486
rect 9338 12484 9394 12486
rect 9098 11450 9154 11452
rect 9178 11450 9234 11452
rect 9258 11450 9314 11452
rect 9338 11450 9394 11452
rect 9098 11398 9144 11450
rect 9144 11398 9154 11450
rect 9178 11398 9208 11450
rect 9208 11398 9220 11450
rect 9220 11398 9234 11450
rect 9258 11398 9272 11450
rect 9272 11398 9284 11450
rect 9284 11398 9314 11450
rect 9338 11398 9348 11450
rect 9348 11398 9394 11450
rect 9098 11396 9154 11398
rect 9178 11396 9234 11398
rect 9258 11396 9314 11398
rect 9338 11396 9394 11398
rect 9098 10362 9154 10364
rect 9178 10362 9234 10364
rect 9258 10362 9314 10364
rect 9338 10362 9394 10364
rect 9098 10310 9144 10362
rect 9144 10310 9154 10362
rect 9178 10310 9208 10362
rect 9208 10310 9220 10362
rect 9220 10310 9234 10362
rect 9258 10310 9272 10362
rect 9272 10310 9284 10362
rect 9284 10310 9314 10362
rect 9338 10310 9348 10362
rect 9348 10310 9394 10362
rect 9098 10308 9154 10310
rect 9178 10308 9234 10310
rect 9258 10308 9314 10310
rect 9338 10308 9394 10310
rect 9098 9274 9154 9276
rect 9178 9274 9234 9276
rect 9258 9274 9314 9276
rect 9338 9274 9394 9276
rect 9098 9222 9144 9274
rect 9144 9222 9154 9274
rect 9178 9222 9208 9274
rect 9208 9222 9220 9274
rect 9220 9222 9234 9274
rect 9258 9222 9272 9274
rect 9272 9222 9284 9274
rect 9284 9222 9314 9274
rect 9338 9222 9348 9274
rect 9348 9222 9394 9274
rect 9098 9220 9154 9222
rect 9178 9220 9234 9222
rect 9258 9220 9314 9222
rect 9338 9220 9394 9222
rect 9098 8186 9154 8188
rect 9178 8186 9234 8188
rect 9258 8186 9314 8188
rect 9338 8186 9394 8188
rect 9098 8134 9144 8186
rect 9144 8134 9154 8186
rect 9178 8134 9208 8186
rect 9208 8134 9220 8186
rect 9220 8134 9234 8186
rect 9258 8134 9272 8186
rect 9272 8134 9284 8186
rect 9284 8134 9314 8186
rect 9338 8134 9348 8186
rect 9348 8134 9394 8186
rect 9098 8132 9154 8134
rect 9178 8132 9234 8134
rect 9258 8132 9314 8134
rect 9338 8132 9394 8134
rect 9098 7098 9154 7100
rect 9178 7098 9234 7100
rect 9258 7098 9314 7100
rect 9338 7098 9394 7100
rect 9098 7046 9144 7098
rect 9144 7046 9154 7098
rect 9178 7046 9208 7098
rect 9208 7046 9220 7098
rect 9220 7046 9234 7098
rect 9258 7046 9272 7098
rect 9272 7046 9284 7098
rect 9284 7046 9314 7098
rect 9338 7046 9348 7098
rect 9348 7046 9394 7098
rect 9098 7044 9154 7046
rect 9178 7044 9234 7046
rect 9258 7044 9314 7046
rect 9338 7044 9394 7046
rect 9098 6010 9154 6012
rect 9178 6010 9234 6012
rect 9258 6010 9314 6012
rect 9338 6010 9394 6012
rect 9098 5958 9144 6010
rect 9144 5958 9154 6010
rect 9178 5958 9208 6010
rect 9208 5958 9220 6010
rect 9220 5958 9234 6010
rect 9258 5958 9272 6010
rect 9272 5958 9284 6010
rect 9284 5958 9314 6010
rect 9338 5958 9348 6010
rect 9348 5958 9394 6010
rect 9098 5956 9154 5958
rect 9178 5956 9234 5958
rect 9258 5956 9314 5958
rect 9338 5956 9394 5958
rect 10230 7384 10286 7440
rect 11812 13082 11868 13084
rect 11892 13082 11948 13084
rect 11972 13082 12028 13084
rect 12052 13082 12108 13084
rect 11812 13030 11858 13082
rect 11858 13030 11868 13082
rect 11892 13030 11922 13082
rect 11922 13030 11934 13082
rect 11934 13030 11948 13082
rect 11972 13030 11986 13082
rect 11986 13030 11998 13082
rect 11998 13030 12028 13082
rect 12052 13030 12062 13082
rect 12062 13030 12108 13082
rect 11812 13028 11868 13030
rect 11892 13028 11948 13030
rect 11972 13028 12028 13030
rect 12052 13028 12108 13030
rect 11812 11994 11868 11996
rect 11892 11994 11948 11996
rect 11972 11994 12028 11996
rect 12052 11994 12108 11996
rect 11812 11942 11858 11994
rect 11858 11942 11868 11994
rect 11892 11942 11922 11994
rect 11922 11942 11934 11994
rect 11934 11942 11948 11994
rect 11972 11942 11986 11994
rect 11986 11942 11998 11994
rect 11998 11942 12028 11994
rect 12052 11942 12062 11994
rect 12062 11942 12108 11994
rect 11812 11940 11868 11942
rect 11892 11940 11948 11942
rect 11972 11940 12028 11942
rect 12052 11940 12108 11942
rect 14526 13626 14582 13628
rect 14606 13626 14662 13628
rect 14686 13626 14742 13628
rect 14766 13626 14822 13628
rect 14526 13574 14572 13626
rect 14572 13574 14582 13626
rect 14606 13574 14636 13626
rect 14636 13574 14648 13626
rect 14648 13574 14662 13626
rect 14686 13574 14700 13626
rect 14700 13574 14712 13626
rect 14712 13574 14742 13626
rect 14766 13574 14776 13626
rect 14776 13574 14822 13626
rect 14526 13572 14582 13574
rect 14606 13572 14662 13574
rect 14686 13572 14742 13574
rect 14766 13572 14822 13574
rect 19954 13626 20010 13628
rect 20034 13626 20090 13628
rect 20114 13626 20170 13628
rect 20194 13626 20250 13628
rect 19954 13574 20000 13626
rect 20000 13574 20010 13626
rect 20034 13574 20064 13626
rect 20064 13574 20076 13626
rect 20076 13574 20090 13626
rect 20114 13574 20128 13626
rect 20128 13574 20140 13626
rect 20140 13574 20170 13626
rect 20194 13574 20204 13626
rect 20204 13574 20250 13626
rect 19954 13572 20010 13574
rect 20034 13572 20090 13574
rect 20114 13572 20170 13574
rect 20194 13572 20250 13574
rect 17240 13082 17296 13084
rect 17320 13082 17376 13084
rect 17400 13082 17456 13084
rect 17480 13082 17536 13084
rect 17240 13030 17286 13082
rect 17286 13030 17296 13082
rect 17320 13030 17350 13082
rect 17350 13030 17362 13082
rect 17362 13030 17376 13082
rect 17400 13030 17414 13082
rect 17414 13030 17426 13082
rect 17426 13030 17456 13082
rect 17480 13030 17490 13082
rect 17490 13030 17536 13082
rect 17240 13028 17296 13030
rect 17320 13028 17376 13030
rect 17400 13028 17456 13030
rect 17480 13028 17536 13030
rect 22668 13082 22724 13084
rect 22748 13082 22804 13084
rect 22828 13082 22884 13084
rect 22908 13082 22964 13084
rect 22668 13030 22714 13082
rect 22714 13030 22724 13082
rect 22748 13030 22778 13082
rect 22778 13030 22790 13082
rect 22790 13030 22804 13082
rect 22828 13030 22842 13082
rect 22842 13030 22854 13082
rect 22854 13030 22884 13082
rect 22908 13030 22918 13082
rect 22918 13030 22964 13082
rect 22668 13028 22724 13030
rect 22748 13028 22804 13030
rect 22828 13028 22884 13030
rect 22908 13028 22964 13030
rect 11812 10906 11868 10908
rect 11892 10906 11948 10908
rect 11972 10906 12028 10908
rect 12052 10906 12108 10908
rect 11812 10854 11858 10906
rect 11858 10854 11868 10906
rect 11892 10854 11922 10906
rect 11922 10854 11934 10906
rect 11934 10854 11948 10906
rect 11972 10854 11986 10906
rect 11986 10854 11998 10906
rect 11998 10854 12028 10906
rect 12052 10854 12062 10906
rect 12062 10854 12108 10906
rect 11812 10852 11868 10854
rect 11892 10852 11948 10854
rect 11972 10852 12028 10854
rect 12052 10852 12108 10854
rect 11812 9818 11868 9820
rect 11892 9818 11948 9820
rect 11972 9818 12028 9820
rect 12052 9818 12108 9820
rect 11812 9766 11858 9818
rect 11858 9766 11868 9818
rect 11892 9766 11922 9818
rect 11922 9766 11934 9818
rect 11934 9766 11948 9818
rect 11972 9766 11986 9818
rect 11986 9766 11998 9818
rect 11998 9766 12028 9818
rect 12052 9766 12062 9818
rect 12062 9766 12108 9818
rect 11812 9764 11868 9766
rect 11892 9764 11948 9766
rect 11972 9764 12028 9766
rect 12052 9764 12108 9766
rect 11812 8730 11868 8732
rect 11892 8730 11948 8732
rect 11972 8730 12028 8732
rect 12052 8730 12108 8732
rect 11812 8678 11858 8730
rect 11858 8678 11868 8730
rect 11892 8678 11922 8730
rect 11922 8678 11934 8730
rect 11934 8678 11948 8730
rect 11972 8678 11986 8730
rect 11986 8678 11998 8730
rect 11998 8678 12028 8730
rect 12052 8678 12062 8730
rect 12062 8678 12108 8730
rect 11812 8676 11868 8678
rect 11892 8676 11948 8678
rect 11972 8676 12028 8678
rect 12052 8676 12108 8678
rect 14526 12538 14582 12540
rect 14606 12538 14662 12540
rect 14686 12538 14742 12540
rect 14766 12538 14822 12540
rect 14526 12486 14572 12538
rect 14572 12486 14582 12538
rect 14606 12486 14636 12538
rect 14636 12486 14648 12538
rect 14648 12486 14662 12538
rect 14686 12486 14700 12538
rect 14700 12486 14712 12538
rect 14712 12486 14742 12538
rect 14766 12486 14776 12538
rect 14776 12486 14822 12538
rect 14526 12484 14582 12486
rect 14606 12484 14662 12486
rect 14686 12484 14742 12486
rect 14766 12484 14822 12486
rect 14526 11450 14582 11452
rect 14606 11450 14662 11452
rect 14686 11450 14742 11452
rect 14766 11450 14822 11452
rect 14526 11398 14572 11450
rect 14572 11398 14582 11450
rect 14606 11398 14636 11450
rect 14636 11398 14648 11450
rect 14648 11398 14662 11450
rect 14686 11398 14700 11450
rect 14700 11398 14712 11450
rect 14712 11398 14742 11450
rect 14766 11398 14776 11450
rect 14776 11398 14822 11450
rect 14526 11396 14582 11398
rect 14606 11396 14662 11398
rect 14686 11396 14742 11398
rect 14766 11396 14822 11398
rect 14526 10362 14582 10364
rect 14606 10362 14662 10364
rect 14686 10362 14742 10364
rect 14766 10362 14822 10364
rect 14526 10310 14572 10362
rect 14572 10310 14582 10362
rect 14606 10310 14636 10362
rect 14636 10310 14648 10362
rect 14648 10310 14662 10362
rect 14686 10310 14700 10362
rect 14700 10310 14712 10362
rect 14712 10310 14742 10362
rect 14766 10310 14776 10362
rect 14776 10310 14822 10362
rect 14526 10308 14582 10310
rect 14606 10308 14662 10310
rect 14686 10308 14742 10310
rect 14766 10308 14822 10310
rect 15198 10512 15254 10568
rect 19954 12538 20010 12540
rect 20034 12538 20090 12540
rect 20114 12538 20170 12540
rect 20194 12538 20250 12540
rect 19954 12486 20000 12538
rect 20000 12486 20010 12538
rect 20034 12486 20064 12538
rect 20064 12486 20076 12538
rect 20076 12486 20090 12538
rect 20114 12486 20128 12538
rect 20128 12486 20140 12538
rect 20140 12486 20170 12538
rect 20194 12486 20204 12538
rect 20204 12486 20250 12538
rect 19954 12484 20010 12486
rect 20034 12484 20090 12486
rect 20114 12484 20170 12486
rect 20194 12484 20250 12486
rect 17240 11994 17296 11996
rect 17320 11994 17376 11996
rect 17400 11994 17456 11996
rect 17480 11994 17536 11996
rect 17240 11942 17286 11994
rect 17286 11942 17296 11994
rect 17320 11942 17350 11994
rect 17350 11942 17362 11994
rect 17362 11942 17376 11994
rect 17400 11942 17414 11994
rect 17414 11942 17426 11994
rect 17426 11942 17456 11994
rect 17480 11942 17490 11994
rect 17490 11942 17536 11994
rect 17240 11940 17296 11942
rect 17320 11940 17376 11942
rect 17400 11940 17456 11942
rect 17480 11940 17536 11942
rect 22668 11994 22724 11996
rect 22748 11994 22804 11996
rect 22828 11994 22884 11996
rect 22908 11994 22964 11996
rect 22668 11942 22714 11994
rect 22714 11942 22724 11994
rect 22748 11942 22778 11994
rect 22778 11942 22790 11994
rect 22790 11942 22804 11994
rect 22828 11942 22842 11994
rect 22842 11942 22854 11994
rect 22854 11942 22884 11994
rect 22908 11942 22918 11994
rect 22918 11942 22964 11994
rect 22668 11940 22724 11942
rect 22748 11940 22804 11942
rect 22828 11940 22884 11942
rect 22908 11940 22964 11942
rect 19954 11450 20010 11452
rect 20034 11450 20090 11452
rect 20114 11450 20170 11452
rect 20194 11450 20250 11452
rect 19954 11398 20000 11450
rect 20000 11398 20010 11450
rect 20034 11398 20064 11450
rect 20064 11398 20076 11450
rect 20076 11398 20090 11450
rect 20114 11398 20128 11450
rect 20128 11398 20140 11450
rect 20140 11398 20170 11450
rect 20194 11398 20204 11450
rect 20204 11398 20250 11450
rect 19954 11396 20010 11398
rect 20034 11396 20090 11398
rect 20114 11396 20170 11398
rect 20194 11396 20250 11398
rect 17240 10906 17296 10908
rect 17320 10906 17376 10908
rect 17400 10906 17456 10908
rect 17480 10906 17536 10908
rect 17240 10854 17286 10906
rect 17286 10854 17296 10906
rect 17320 10854 17350 10906
rect 17350 10854 17362 10906
rect 17362 10854 17376 10906
rect 17400 10854 17414 10906
rect 17414 10854 17426 10906
rect 17426 10854 17456 10906
rect 17480 10854 17490 10906
rect 17490 10854 17536 10906
rect 17240 10852 17296 10854
rect 17320 10852 17376 10854
rect 17400 10852 17456 10854
rect 17480 10852 17536 10854
rect 22668 10906 22724 10908
rect 22748 10906 22804 10908
rect 22828 10906 22884 10908
rect 22908 10906 22964 10908
rect 22668 10854 22714 10906
rect 22714 10854 22724 10906
rect 22748 10854 22778 10906
rect 22778 10854 22790 10906
rect 22790 10854 22804 10906
rect 22828 10854 22842 10906
rect 22842 10854 22854 10906
rect 22854 10854 22884 10906
rect 22908 10854 22918 10906
rect 22918 10854 22964 10906
rect 22668 10852 22724 10854
rect 22748 10852 22804 10854
rect 22828 10852 22884 10854
rect 22908 10852 22964 10854
rect 19954 10362 20010 10364
rect 20034 10362 20090 10364
rect 20114 10362 20170 10364
rect 20194 10362 20250 10364
rect 19954 10310 20000 10362
rect 20000 10310 20010 10362
rect 20034 10310 20064 10362
rect 20064 10310 20076 10362
rect 20076 10310 20090 10362
rect 20114 10310 20128 10362
rect 20128 10310 20140 10362
rect 20140 10310 20170 10362
rect 20194 10310 20204 10362
rect 20204 10310 20250 10362
rect 19954 10308 20010 10310
rect 20034 10308 20090 10310
rect 20114 10308 20170 10310
rect 20194 10308 20250 10310
rect 14526 9274 14582 9276
rect 14606 9274 14662 9276
rect 14686 9274 14742 9276
rect 14766 9274 14822 9276
rect 14526 9222 14572 9274
rect 14572 9222 14582 9274
rect 14606 9222 14636 9274
rect 14636 9222 14648 9274
rect 14648 9222 14662 9274
rect 14686 9222 14700 9274
rect 14700 9222 14712 9274
rect 14712 9222 14742 9274
rect 14766 9222 14776 9274
rect 14776 9222 14822 9274
rect 14526 9220 14582 9222
rect 14606 9220 14662 9222
rect 14686 9220 14742 9222
rect 14766 9220 14822 9222
rect 11812 7642 11868 7644
rect 11892 7642 11948 7644
rect 11972 7642 12028 7644
rect 12052 7642 12108 7644
rect 11812 7590 11858 7642
rect 11858 7590 11868 7642
rect 11892 7590 11922 7642
rect 11922 7590 11934 7642
rect 11934 7590 11948 7642
rect 11972 7590 11986 7642
rect 11986 7590 11998 7642
rect 11998 7590 12028 7642
rect 12052 7590 12062 7642
rect 12062 7590 12108 7642
rect 11812 7588 11868 7590
rect 11892 7588 11948 7590
rect 11972 7588 12028 7590
rect 12052 7588 12108 7590
rect 11150 6704 11206 6760
rect 11812 6554 11868 6556
rect 11892 6554 11948 6556
rect 11972 6554 12028 6556
rect 12052 6554 12108 6556
rect 11812 6502 11858 6554
rect 11858 6502 11868 6554
rect 11892 6502 11922 6554
rect 11922 6502 11934 6554
rect 11934 6502 11948 6554
rect 11972 6502 11986 6554
rect 11986 6502 11998 6554
rect 11998 6502 12028 6554
rect 12052 6502 12062 6554
rect 12062 6502 12108 6554
rect 11812 6500 11868 6502
rect 11892 6500 11948 6502
rect 11972 6500 12028 6502
rect 12052 6500 12108 6502
rect 11812 5466 11868 5468
rect 11892 5466 11948 5468
rect 11972 5466 12028 5468
rect 12052 5466 12108 5468
rect 11812 5414 11858 5466
rect 11858 5414 11868 5466
rect 11892 5414 11922 5466
rect 11922 5414 11934 5466
rect 11934 5414 11948 5466
rect 11972 5414 11986 5466
rect 11986 5414 11998 5466
rect 11998 5414 12028 5466
rect 12052 5414 12062 5466
rect 12062 5414 12108 5466
rect 11812 5412 11868 5414
rect 11892 5412 11948 5414
rect 11972 5412 12028 5414
rect 12052 5412 12108 5414
rect 9098 4922 9154 4924
rect 9178 4922 9234 4924
rect 9258 4922 9314 4924
rect 9338 4922 9394 4924
rect 9098 4870 9144 4922
rect 9144 4870 9154 4922
rect 9178 4870 9208 4922
rect 9208 4870 9220 4922
rect 9220 4870 9234 4922
rect 9258 4870 9272 4922
rect 9272 4870 9284 4922
rect 9284 4870 9314 4922
rect 9338 4870 9348 4922
rect 9348 4870 9394 4922
rect 9098 4868 9154 4870
rect 9178 4868 9234 4870
rect 9258 4868 9314 4870
rect 9338 4868 9394 4870
rect 9098 3834 9154 3836
rect 9178 3834 9234 3836
rect 9258 3834 9314 3836
rect 9338 3834 9394 3836
rect 9098 3782 9144 3834
rect 9144 3782 9154 3834
rect 9178 3782 9208 3834
rect 9208 3782 9220 3834
rect 9220 3782 9234 3834
rect 9258 3782 9272 3834
rect 9272 3782 9284 3834
rect 9284 3782 9314 3834
rect 9338 3782 9348 3834
rect 9348 3782 9394 3834
rect 9098 3780 9154 3782
rect 9178 3780 9234 3782
rect 9258 3780 9314 3782
rect 9338 3780 9394 3782
rect 11812 4378 11868 4380
rect 11892 4378 11948 4380
rect 11972 4378 12028 4380
rect 12052 4378 12108 4380
rect 11812 4326 11858 4378
rect 11858 4326 11868 4378
rect 11892 4326 11922 4378
rect 11922 4326 11934 4378
rect 11934 4326 11948 4378
rect 11972 4326 11986 4378
rect 11986 4326 11998 4378
rect 11998 4326 12028 4378
rect 12052 4326 12062 4378
rect 12062 4326 12108 4378
rect 11812 4324 11868 4326
rect 11892 4324 11948 4326
rect 11972 4324 12028 4326
rect 12052 4324 12108 4326
rect 9098 2746 9154 2748
rect 9178 2746 9234 2748
rect 9258 2746 9314 2748
rect 9338 2746 9394 2748
rect 9098 2694 9144 2746
rect 9144 2694 9154 2746
rect 9178 2694 9208 2746
rect 9208 2694 9220 2746
rect 9220 2694 9234 2746
rect 9258 2694 9272 2746
rect 9272 2694 9284 2746
rect 9284 2694 9314 2746
rect 9338 2694 9348 2746
rect 9348 2694 9394 2746
rect 9098 2692 9154 2694
rect 9178 2692 9234 2694
rect 9258 2692 9314 2694
rect 9338 2692 9394 2694
rect 11812 3290 11868 3292
rect 11892 3290 11948 3292
rect 11972 3290 12028 3292
rect 12052 3290 12108 3292
rect 11812 3238 11858 3290
rect 11858 3238 11868 3290
rect 11892 3238 11922 3290
rect 11922 3238 11934 3290
rect 11934 3238 11948 3290
rect 11972 3238 11986 3290
rect 11986 3238 11998 3290
rect 11998 3238 12028 3290
rect 12052 3238 12062 3290
rect 12062 3238 12108 3290
rect 11812 3236 11868 3238
rect 11892 3236 11948 3238
rect 11972 3236 12028 3238
rect 12052 3236 12108 3238
rect 14526 8186 14582 8188
rect 14606 8186 14662 8188
rect 14686 8186 14742 8188
rect 14766 8186 14822 8188
rect 14526 8134 14572 8186
rect 14572 8134 14582 8186
rect 14606 8134 14636 8186
rect 14636 8134 14648 8186
rect 14648 8134 14662 8186
rect 14686 8134 14700 8186
rect 14700 8134 14712 8186
rect 14712 8134 14742 8186
rect 14766 8134 14776 8186
rect 14776 8134 14822 8186
rect 14526 8132 14582 8134
rect 14606 8132 14662 8134
rect 14686 8132 14742 8134
rect 14766 8132 14822 8134
rect 14526 7098 14582 7100
rect 14606 7098 14662 7100
rect 14686 7098 14742 7100
rect 14766 7098 14822 7100
rect 14526 7046 14572 7098
rect 14572 7046 14582 7098
rect 14606 7046 14636 7098
rect 14636 7046 14648 7098
rect 14648 7046 14662 7098
rect 14686 7046 14700 7098
rect 14700 7046 14712 7098
rect 14712 7046 14742 7098
rect 14766 7046 14776 7098
rect 14776 7046 14822 7098
rect 14526 7044 14582 7046
rect 14606 7044 14662 7046
rect 14686 7044 14742 7046
rect 14766 7044 14822 7046
rect 14526 6010 14582 6012
rect 14606 6010 14662 6012
rect 14686 6010 14742 6012
rect 14766 6010 14822 6012
rect 14526 5958 14572 6010
rect 14572 5958 14582 6010
rect 14606 5958 14636 6010
rect 14636 5958 14648 6010
rect 14648 5958 14662 6010
rect 14686 5958 14700 6010
rect 14700 5958 14712 6010
rect 14712 5958 14742 6010
rect 14766 5958 14776 6010
rect 14776 5958 14822 6010
rect 14526 5956 14582 5958
rect 14606 5956 14662 5958
rect 14686 5956 14742 5958
rect 14766 5956 14822 5958
rect 13910 3984 13966 4040
rect 14526 4922 14582 4924
rect 14606 4922 14662 4924
rect 14686 4922 14742 4924
rect 14766 4922 14822 4924
rect 14526 4870 14572 4922
rect 14572 4870 14582 4922
rect 14606 4870 14636 4922
rect 14636 4870 14648 4922
rect 14648 4870 14662 4922
rect 14686 4870 14700 4922
rect 14700 4870 14712 4922
rect 14712 4870 14742 4922
rect 14766 4870 14776 4922
rect 14776 4870 14822 4922
rect 14526 4868 14582 4870
rect 14606 4868 14662 4870
rect 14686 4868 14742 4870
rect 14766 4868 14822 4870
rect 14526 3834 14582 3836
rect 14606 3834 14662 3836
rect 14686 3834 14742 3836
rect 14766 3834 14822 3836
rect 14526 3782 14572 3834
rect 14572 3782 14582 3834
rect 14606 3782 14636 3834
rect 14636 3782 14648 3834
rect 14648 3782 14662 3834
rect 14686 3782 14700 3834
rect 14700 3782 14712 3834
rect 14712 3782 14742 3834
rect 14766 3782 14776 3834
rect 14776 3782 14822 3834
rect 14526 3780 14582 3782
rect 14606 3780 14662 3782
rect 14686 3780 14742 3782
rect 14766 3780 14822 3782
rect 14526 2746 14582 2748
rect 14606 2746 14662 2748
rect 14686 2746 14742 2748
rect 14766 2746 14822 2748
rect 14526 2694 14572 2746
rect 14572 2694 14582 2746
rect 14606 2694 14636 2746
rect 14636 2694 14648 2746
rect 14648 2694 14662 2746
rect 14686 2694 14700 2746
rect 14700 2694 14712 2746
rect 14712 2694 14742 2746
rect 14766 2694 14776 2746
rect 14776 2694 14822 2746
rect 14526 2692 14582 2694
rect 14606 2692 14662 2694
rect 14686 2692 14742 2694
rect 14766 2692 14822 2694
rect 17240 9818 17296 9820
rect 17320 9818 17376 9820
rect 17400 9818 17456 9820
rect 17480 9818 17536 9820
rect 17240 9766 17286 9818
rect 17286 9766 17296 9818
rect 17320 9766 17350 9818
rect 17350 9766 17362 9818
rect 17362 9766 17376 9818
rect 17400 9766 17414 9818
rect 17414 9766 17426 9818
rect 17426 9766 17456 9818
rect 17480 9766 17490 9818
rect 17490 9766 17536 9818
rect 17240 9764 17296 9766
rect 17320 9764 17376 9766
rect 17400 9764 17456 9766
rect 17480 9764 17536 9766
rect 22668 9818 22724 9820
rect 22748 9818 22804 9820
rect 22828 9818 22884 9820
rect 22908 9818 22964 9820
rect 22668 9766 22714 9818
rect 22714 9766 22724 9818
rect 22748 9766 22778 9818
rect 22778 9766 22790 9818
rect 22790 9766 22804 9818
rect 22828 9766 22842 9818
rect 22842 9766 22854 9818
rect 22854 9766 22884 9818
rect 22908 9766 22918 9818
rect 22918 9766 22964 9818
rect 22668 9764 22724 9766
rect 22748 9764 22804 9766
rect 22828 9764 22884 9766
rect 22908 9764 22964 9766
rect 19954 9274 20010 9276
rect 20034 9274 20090 9276
rect 20114 9274 20170 9276
rect 20194 9274 20250 9276
rect 19954 9222 20000 9274
rect 20000 9222 20010 9274
rect 20034 9222 20064 9274
rect 20064 9222 20076 9274
rect 20076 9222 20090 9274
rect 20114 9222 20128 9274
rect 20128 9222 20140 9274
rect 20140 9222 20170 9274
rect 20194 9222 20204 9274
rect 20204 9222 20250 9274
rect 19954 9220 20010 9222
rect 20034 9220 20090 9222
rect 20114 9220 20170 9222
rect 20194 9220 20250 9222
rect 17240 8730 17296 8732
rect 17320 8730 17376 8732
rect 17400 8730 17456 8732
rect 17480 8730 17536 8732
rect 17240 8678 17286 8730
rect 17286 8678 17296 8730
rect 17320 8678 17350 8730
rect 17350 8678 17362 8730
rect 17362 8678 17376 8730
rect 17400 8678 17414 8730
rect 17414 8678 17426 8730
rect 17426 8678 17456 8730
rect 17480 8678 17490 8730
rect 17490 8678 17536 8730
rect 17240 8676 17296 8678
rect 17320 8676 17376 8678
rect 17400 8676 17456 8678
rect 17480 8676 17536 8678
rect 17240 7642 17296 7644
rect 17320 7642 17376 7644
rect 17400 7642 17456 7644
rect 17480 7642 17536 7644
rect 17240 7590 17286 7642
rect 17286 7590 17296 7642
rect 17320 7590 17350 7642
rect 17350 7590 17362 7642
rect 17362 7590 17376 7642
rect 17400 7590 17414 7642
rect 17414 7590 17426 7642
rect 17426 7590 17456 7642
rect 17480 7590 17490 7642
rect 17490 7590 17536 7642
rect 17240 7588 17296 7590
rect 17320 7588 17376 7590
rect 17400 7588 17456 7590
rect 17480 7588 17536 7590
rect 17406 7384 17462 7440
rect 17240 6554 17296 6556
rect 17320 6554 17376 6556
rect 17400 6554 17456 6556
rect 17480 6554 17536 6556
rect 17240 6502 17286 6554
rect 17286 6502 17296 6554
rect 17320 6502 17350 6554
rect 17350 6502 17362 6554
rect 17362 6502 17376 6554
rect 17400 6502 17414 6554
rect 17414 6502 17426 6554
rect 17426 6502 17456 6554
rect 17480 6502 17490 6554
rect 17490 6502 17536 6554
rect 17240 6500 17296 6502
rect 17320 6500 17376 6502
rect 17400 6500 17456 6502
rect 17480 6500 17536 6502
rect 17240 5466 17296 5468
rect 17320 5466 17376 5468
rect 17400 5466 17456 5468
rect 17480 5466 17536 5468
rect 17240 5414 17286 5466
rect 17286 5414 17296 5466
rect 17320 5414 17350 5466
rect 17350 5414 17362 5466
rect 17362 5414 17376 5466
rect 17400 5414 17414 5466
rect 17414 5414 17426 5466
rect 17426 5414 17456 5466
rect 17480 5414 17490 5466
rect 17490 5414 17536 5466
rect 17240 5412 17296 5414
rect 17320 5412 17376 5414
rect 17400 5412 17456 5414
rect 17480 5412 17536 5414
rect 17240 4378 17296 4380
rect 17320 4378 17376 4380
rect 17400 4378 17456 4380
rect 17480 4378 17536 4380
rect 17240 4326 17286 4378
rect 17286 4326 17296 4378
rect 17320 4326 17350 4378
rect 17350 4326 17362 4378
rect 17362 4326 17376 4378
rect 17400 4326 17414 4378
rect 17414 4326 17426 4378
rect 17426 4326 17456 4378
rect 17480 4326 17490 4378
rect 17490 4326 17536 4378
rect 17240 4324 17296 4326
rect 17320 4324 17376 4326
rect 17400 4324 17456 4326
rect 17480 4324 17536 4326
rect 17240 3290 17296 3292
rect 17320 3290 17376 3292
rect 17400 3290 17456 3292
rect 17480 3290 17536 3292
rect 17240 3238 17286 3290
rect 17286 3238 17296 3290
rect 17320 3238 17350 3290
rect 17350 3238 17362 3290
rect 17362 3238 17376 3290
rect 17400 3238 17414 3290
rect 17414 3238 17426 3290
rect 17426 3238 17456 3290
rect 17480 3238 17490 3290
rect 17490 3238 17536 3290
rect 17240 3236 17296 3238
rect 17320 3236 17376 3238
rect 17400 3236 17456 3238
rect 17480 3236 17536 3238
rect 19430 5752 19486 5808
rect 22668 8730 22724 8732
rect 22748 8730 22804 8732
rect 22828 8730 22884 8732
rect 22908 8730 22964 8732
rect 22668 8678 22714 8730
rect 22714 8678 22724 8730
rect 22748 8678 22778 8730
rect 22778 8678 22790 8730
rect 22790 8678 22804 8730
rect 22828 8678 22842 8730
rect 22842 8678 22854 8730
rect 22854 8678 22884 8730
rect 22908 8678 22918 8730
rect 22918 8678 22964 8730
rect 22668 8676 22724 8678
rect 22748 8676 22804 8678
rect 22828 8676 22884 8678
rect 22908 8676 22964 8678
rect 19954 8186 20010 8188
rect 20034 8186 20090 8188
rect 20114 8186 20170 8188
rect 20194 8186 20250 8188
rect 19954 8134 20000 8186
rect 20000 8134 20010 8186
rect 20034 8134 20064 8186
rect 20064 8134 20076 8186
rect 20076 8134 20090 8186
rect 20114 8134 20128 8186
rect 20128 8134 20140 8186
rect 20140 8134 20170 8186
rect 20194 8134 20204 8186
rect 20204 8134 20250 8186
rect 19954 8132 20010 8134
rect 20034 8132 20090 8134
rect 20114 8132 20170 8134
rect 20194 8132 20250 8134
rect 19954 7098 20010 7100
rect 20034 7098 20090 7100
rect 20114 7098 20170 7100
rect 20194 7098 20250 7100
rect 19954 7046 20000 7098
rect 20000 7046 20010 7098
rect 20034 7046 20064 7098
rect 20064 7046 20076 7098
rect 20076 7046 20090 7098
rect 20114 7046 20128 7098
rect 20128 7046 20140 7098
rect 20140 7046 20170 7098
rect 20194 7046 20204 7098
rect 20204 7046 20250 7098
rect 19954 7044 20010 7046
rect 20034 7044 20090 7046
rect 20114 7044 20170 7046
rect 20194 7044 20250 7046
rect 19614 6296 19670 6352
rect 19614 5652 19616 5672
rect 19616 5652 19668 5672
rect 19668 5652 19670 5672
rect 19614 5616 19670 5652
rect 19062 3984 19118 4040
rect 19954 6010 20010 6012
rect 20034 6010 20090 6012
rect 20114 6010 20170 6012
rect 20194 6010 20250 6012
rect 19954 5958 20000 6010
rect 20000 5958 20010 6010
rect 20034 5958 20064 6010
rect 20064 5958 20076 6010
rect 20076 5958 20090 6010
rect 20114 5958 20128 6010
rect 20128 5958 20140 6010
rect 20140 5958 20170 6010
rect 20194 5958 20204 6010
rect 20204 5958 20250 6010
rect 19954 5956 20010 5958
rect 20034 5956 20090 5958
rect 20114 5956 20170 5958
rect 20194 5956 20250 5958
rect 22668 7642 22724 7644
rect 22748 7642 22804 7644
rect 22828 7642 22884 7644
rect 22908 7642 22964 7644
rect 22668 7590 22714 7642
rect 22714 7590 22724 7642
rect 22748 7590 22778 7642
rect 22778 7590 22790 7642
rect 22790 7590 22804 7642
rect 22828 7590 22842 7642
rect 22842 7590 22854 7642
rect 22854 7590 22884 7642
rect 22908 7590 22918 7642
rect 22918 7590 22964 7642
rect 22668 7588 22724 7590
rect 22748 7588 22804 7590
rect 22828 7588 22884 7590
rect 22908 7588 22964 7590
rect 19954 4922 20010 4924
rect 20034 4922 20090 4924
rect 20114 4922 20170 4924
rect 20194 4922 20250 4924
rect 19954 4870 20000 4922
rect 20000 4870 20010 4922
rect 20034 4870 20064 4922
rect 20064 4870 20076 4922
rect 20076 4870 20090 4922
rect 20114 4870 20128 4922
rect 20128 4870 20140 4922
rect 20140 4870 20170 4922
rect 20194 4870 20204 4922
rect 20204 4870 20250 4922
rect 19954 4868 20010 4870
rect 20034 4868 20090 4870
rect 20114 4868 20170 4870
rect 20194 4868 20250 4870
rect 19954 3834 20010 3836
rect 20034 3834 20090 3836
rect 20114 3834 20170 3836
rect 20194 3834 20250 3836
rect 19954 3782 20000 3834
rect 20000 3782 20010 3834
rect 20034 3782 20064 3834
rect 20064 3782 20076 3834
rect 20076 3782 20090 3834
rect 20114 3782 20128 3834
rect 20128 3782 20140 3834
rect 20140 3782 20170 3834
rect 20194 3782 20204 3834
rect 20204 3782 20250 3834
rect 19954 3780 20010 3782
rect 20034 3780 20090 3782
rect 20114 3780 20170 3782
rect 20194 3780 20250 3782
rect 22668 6554 22724 6556
rect 22748 6554 22804 6556
rect 22828 6554 22884 6556
rect 22908 6554 22964 6556
rect 22668 6502 22714 6554
rect 22714 6502 22724 6554
rect 22748 6502 22778 6554
rect 22778 6502 22790 6554
rect 22790 6502 22804 6554
rect 22828 6502 22842 6554
rect 22842 6502 22854 6554
rect 22854 6502 22884 6554
rect 22908 6502 22918 6554
rect 22918 6502 22964 6554
rect 22668 6500 22724 6502
rect 22748 6500 22804 6502
rect 22828 6500 22884 6502
rect 22908 6500 22964 6502
rect 22668 5466 22724 5468
rect 22748 5466 22804 5468
rect 22828 5466 22884 5468
rect 22908 5466 22964 5468
rect 22668 5414 22714 5466
rect 22714 5414 22724 5466
rect 22748 5414 22778 5466
rect 22778 5414 22790 5466
rect 22790 5414 22804 5466
rect 22828 5414 22842 5466
rect 22842 5414 22854 5466
rect 22854 5414 22884 5466
rect 22908 5414 22918 5466
rect 22918 5414 22964 5466
rect 22668 5412 22724 5414
rect 22748 5412 22804 5414
rect 22828 5412 22884 5414
rect 22908 5412 22964 5414
rect 22668 4378 22724 4380
rect 22748 4378 22804 4380
rect 22828 4378 22884 4380
rect 22908 4378 22964 4380
rect 22668 4326 22714 4378
rect 22714 4326 22724 4378
rect 22748 4326 22778 4378
rect 22778 4326 22790 4378
rect 22790 4326 22804 4378
rect 22828 4326 22842 4378
rect 22842 4326 22854 4378
rect 22854 4326 22884 4378
rect 22908 4326 22918 4378
rect 22918 4326 22964 4378
rect 22668 4324 22724 4326
rect 22748 4324 22804 4326
rect 22828 4324 22884 4326
rect 22908 4324 22964 4326
rect 22668 3290 22724 3292
rect 22748 3290 22804 3292
rect 22828 3290 22884 3292
rect 22908 3290 22964 3292
rect 22668 3238 22714 3290
rect 22714 3238 22724 3290
rect 22748 3238 22778 3290
rect 22778 3238 22790 3290
rect 22790 3238 22804 3290
rect 22828 3238 22842 3290
rect 22842 3238 22854 3290
rect 22854 3238 22884 3290
rect 22908 3238 22918 3290
rect 22918 3238 22964 3290
rect 22668 3236 22724 3238
rect 22748 3236 22804 3238
rect 22828 3236 22884 3238
rect 22908 3236 22964 3238
rect 19954 2746 20010 2748
rect 20034 2746 20090 2748
rect 20114 2746 20170 2748
rect 20194 2746 20250 2748
rect 19954 2694 20000 2746
rect 20000 2694 20010 2746
rect 20034 2694 20064 2746
rect 20064 2694 20076 2746
rect 20076 2694 20090 2746
rect 20114 2694 20128 2746
rect 20128 2694 20140 2746
rect 20140 2694 20170 2746
rect 20194 2694 20204 2746
rect 20204 2694 20250 2746
rect 19954 2692 20010 2694
rect 20034 2692 20090 2694
rect 20114 2692 20170 2694
rect 20194 2692 20250 2694
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6430 2202
rect 6430 2150 6440 2202
rect 6464 2150 6494 2202
rect 6494 2150 6506 2202
rect 6506 2150 6520 2202
rect 6544 2150 6558 2202
rect 6558 2150 6570 2202
rect 6570 2150 6600 2202
rect 6624 2150 6634 2202
rect 6634 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 11812 2202 11868 2204
rect 11892 2202 11948 2204
rect 11972 2202 12028 2204
rect 12052 2202 12108 2204
rect 11812 2150 11858 2202
rect 11858 2150 11868 2202
rect 11892 2150 11922 2202
rect 11922 2150 11934 2202
rect 11934 2150 11948 2202
rect 11972 2150 11986 2202
rect 11986 2150 11998 2202
rect 11998 2150 12028 2202
rect 12052 2150 12062 2202
rect 12062 2150 12108 2202
rect 11812 2148 11868 2150
rect 11892 2148 11948 2150
rect 11972 2148 12028 2150
rect 12052 2148 12108 2150
rect 17240 2202 17296 2204
rect 17320 2202 17376 2204
rect 17400 2202 17456 2204
rect 17480 2202 17536 2204
rect 17240 2150 17286 2202
rect 17286 2150 17296 2202
rect 17320 2150 17350 2202
rect 17350 2150 17362 2202
rect 17362 2150 17376 2202
rect 17400 2150 17414 2202
rect 17414 2150 17426 2202
rect 17426 2150 17456 2202
rect 17480 2150 17490 2202
rect 17490 2150 17536 2202
rect 17240 2148 17296 2150
rect 17320 2148 17376 2150
rect 17400 2148 17456 2150
rect 17480 2148 17536 2150
rect 22668 2202 22724 2204
rect 22748 2202 22804 2204
rect 22828 2202 22884 2204
rect 22908 2202 22964 2204
rect 22668 2150 22714 2202
rect 22714 2150 22724 2202
rect 22748 2150 22778 2202
rect 22778 2150 22790 2202
rect 22790 2150 22804 2202
rect 22828 2150 22842 2202
rect 22842 2150 22854 2202
rect 22854 2150 22884 2202
rect 22908 2150 22918 2202
rect 22918 2150 22964 2202
rect 22668 2148 22724 2150
rect 22748 2148 22804 2150
rect 22828 2148 22884 2150
rect 22908 2148 22964 2150
<< metal3 >>
rect 6374 21792 6690 21793
rect 6374 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6690 21792
rect 6374 21727 6690 21728
rect 11802 21792 12118 21793
rect 11802 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12118 21792
rect 11802 21727 12118 21728
rect 17230 21792 17546 21793
rect 17230 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17546 21792
rect 17230 21727 17546 21728
rect 22658 21792 22974 21793
rect 22658 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22974 21792
rect 22658 21727 22974 21728
rect 3660 21248 3976 21249
rect 3660 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3976 21248
rect 3660 21183 3976 21184
rect 9088 21248 9404 21249
rect 9088 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9404 21248
rect 9088 21183 9404 21184
rect 14516 21248 14832 21249
rect 14516 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14832 21248
rect 14516 21183 14832 21184
rect 19944 21248 20260 21249
rect 19944 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20260 21248
rect 19944 21183 20260 21184
rect 6374 20704 6690 20705
rect 6374 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6690 20704
rect 6374 20639 6690 20640
rect 11802 20704 12118 20705
rect 11802 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12118 20704
rect 11802 20639 12118 20640
rect 17230 20704 17546 20705
rect 17230 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17546 20704
rect 17230 20639 17546 20640
rect 22658 20704 22974 20705
rect 22658 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22974 20704
rect 22658 20639 22974 20640
rect 3660 20160 3976 20161
rect 3660 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3976 20160
rect 3660 20095 3976 20096
rect 9088 20160 9404 20161
rect 9088 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9404 20160
rect 9088 20095 9404 20096
rect 14516 20160 14832 20161
rect 14516 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14832 20160
rect 14516 20095 14832 20096
rect 19944 20160 20260 20161
rect 19944 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20260 20160
rect 19944 20095 20260 20096
rect 0 19818 800 19908
rect 2129 19818 2195 19821
rect 0 19816 2195 19818
rect 0 19760 2134 19816
rect 2190 19760 2195 19816
rect 0 19758 2195 19760
rect 0 19668 800 19758
rect 2129 19755 2195 19758
rect 6374 19616 6690 19617
rect 6374 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6690 19616
rect 6374 19551 6690 19552
rect 11802 19616 12118 19617
rect 11802 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12118 19616
rect 11802 19551 12118 19552
rect 17230 19616 17546 19617
rect 17230 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17546 19616
rect 17230 19551 17546 19552
rect 22658 19616 22974 19617
rect 22658 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22974 19616
rect 22658 19551 22974 19552
rect 3660 19072 3976 19073
rect 3660 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3976 19072
rect 3660 19007 3976 19008
rect 9088 19072 9404 19073
rect 9088 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9404 19072
rect 9088 19007 9404 19008
rect 14516 19072 14832 19073
rect 14516 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14832 19072
rect 14516 19007 14832 19008
rect 19944 19072 20260 19073
rect 19944 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20260 19072
rect 19944 19007 20260 19008
rect 6374 18528 6690 18529
rect 6374 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6690 18528
rect 6374 18463 6690 18464
rect 11802 18528 12118 18529
rect 11802 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12118 18528
rect 11802 18463 12118 18464
rect 17230 18528 17546 18529
rect 17230 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17546 18528
rect 17230 18463 17546 18464
rect 22658 18528 22974 18529
rect 22658 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22974 18528
rect 22658 18463 22974 18464
rect 3660 17984 3976 17985
rect 3660 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3976 17984
rect 3660 17919 3976 17920
rect 9088 17984 9404 17985
rect 9088 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9404 17984
rect 9088 17919 9404 17920
rect 14516 17984 14832 17985
rect 14516 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14832 17984
rect 14516 17919 14832 17920
rect 19944 17984 20260 17985
rect 19944 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20260 17984
rect 19944 17919 20260 17920
rect 6374 17440 6690 17441
rect 6374 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6690 17440
rect 6374 17375 6690 17376
rect 11802 17440 12118 17441
rect 11802 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12118 17440
rect 11802 17375 12118 17376
rect 17230 17440 17546 17441
rect 17230 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17546 17440
rect 17230 17375 17546 17376
rect 22658 17440 22974 17441
rect 22658 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22974 17440
rect 22658 17375 22974 17376
rect 3660 16896 3976 16897
rect 3660 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3976 16896
rect 3660 16831 3976 16832
rect 9088 16896 9404 16897
rect 9088 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9404 16896
rect 9088 16831 9404 16832
rect 14516 16896 14832 16897
rect 14516 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14832 16896
rect 14516 16831 14832 16832
rect 19944 16896 20260 16897
rect 19944 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20260 16896
rect 19944 16831 20260 16832
rect 6374 16352 6690 16353
rect 6374 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6690 16352
rect 6374 16287 6690 16288
rect 11802 16352 12118 16353
rect 11802 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12118 16352
rect 11802 16287 12118 16288
rect 17230 16352 17546 16353
rect 17230 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17546 16352
rect 17230 16287 17546 16288
rect 22658 16352 22974 16353
rect 22658 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22974 16352
rect 22658 16287 22974 16288
rect 3660 15808 3976 15809
rect 3660 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3976 15808
rect 3660 15743 3976 15744
rect 9088 15808 9404 15809
rect 9088 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9404 15808
rect 9088 15743 9404 15744
rect 14516 15808 14832 15809
rect 14516 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14832 15808
rect 14516 15743 14832 15744
rect 19944 15808 20260 15809
rect 19944 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20260 15808
rect 19944 15743 20260 15744
rect 6374 15264 6690 15265
rect 6374 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6690 15264
rect 6374 15199 6690 15200
rect 11802 15264 12118 15265
rect 11802 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12118 15264
rect 11802 15199 12118 15200
rect 17230 15264 17546 15265
rect 17230 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17546 15264
rect 17230 15199 17546 15200
rect 22658 15264 22974 15265
rect 22658 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22974 15264
rect 22658 15199 22974 15200
rect 3509 14922 3575 14925
rect 8937 14922 9003 14925
rect 3509 14920 9003 14922
rect 3509 14864 3514 14920
rect 3570 14864 8942 14920
rect 8998 14864 9003 14920
rect 3509 14862 9003 14864
rect 3509 14859 3575 14862
rect 8937 14859 9003 14862
rect 3660 14720 3976 14721
rect 3660 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3976 14720
rect 3660 14655 3976 14656
rect 9088 14720 9404 14721
rect 9088 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9404 14720
rect 9088 14655 9404 14656
rect 14516 14720 14832 14721
rect 14516 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14832 14720
rect 14516 14655 14832 14656
rect 19944 14720 20260 14721
rect 19944 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20260 14720
rect 19944 14655 20260 14656
rect 6374 14176 6690 14177
rect 6374 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6690 14176
rect 6374 14111 6690 14112
rect 11802 14176 12118 14177
rect 11802 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12118 14176
rect 11802 14111 12118 14112
rect 17230 14176 17546 14177
rect 17230 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17546 14176
rect 17230 14111 17546 14112
rect 22658 14176 22974 14177
rect 22658 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22974 14176
rect 22658 14111 22974 14112
rect 3660 13632 3976 13633
rect 3660 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3976 13632
rect 3660 13567 3976 13568
rect 9088 13632 9404 13633
rect 9088 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9404 13632
rect 9088 13567 9404 13568
rect 14516 13632 14832 13633
rect 14516 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14832 13632
rect 14516 13567 14832 13568
rect 19944 13632 20260 13633
rect 19944 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20260 13632
rect 19944 13567 20260 13568
rect 6374 13088 6690 13089
rect 6374 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6690 13088
rect 6374 13023 6690 13024
rect 11802 13088 12118 13089
rect 11802 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12118 13088
rect 11802 13023 12118 13024
rect 17230 13088 17546 13089
rect 17230 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17546 13088
rect 17230 13023 17546 13024
rect 22658 13088 22974 13089
rect 22658 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22974 13088
rect 22658 13023 22974 13024
rect 3660 12544 3976 12545
rect 3660 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3976 12544
rect 3660 12479 3976 12480
rect 9088 12544 9404 12545
rect 9088 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9404 12544
rect 9088 12479 9404 12480
rect 14516 12544 14832 12545
rect 14516 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14832 12544
rect 14516 12479 14832 12480
rect 19944 12544 20260 12545
rect 19944 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20260 12544
rect 19944 12479 20260 12480
rect 0 11930 800 12020
rect 6374 12000 6690 12001
rect 6374 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6690 12000
rect 6374 11935 6690 11936
rect 11802 12000 12118 12001
rect 11802 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12118 12000
rect 11802 11935 12118 11936
rect 17230 12000 17546 12001
rect 17230 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17546 12000
rect 17230 11935 17546 11936
rect 22658 12000 22974 12001
rect 22658 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22974 12000
rect 22658 11935 22974 11936
rect 2773 11930 2839 11933
rect 0 11928 2839 11930
rect 0 11872 2778 11928
rect 2834 11872 2839 11928
rect 0 11870 2839 11872
rect 0 11780 800 11870
rect 2773 11867 2839 11870
rect 3660 11456 3976 11457
rect 3660 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3976 11456
rect 3660 11391 3976 11392
rect 9088 11456 9404 11457
rect 9088 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9404 11456
rect 9088 11391 9404 11392
rect 14516 11456 14832 11457
rect 14516 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14832 11456
rect 14516 11391 14832 11392
rect 19944 11456 20260 11457
rect 19944 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20260 11456
rect 19944 11391 20260 11392
rect 6374 10912 6690 10913
rect 6374 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6690 10912
rect 6374 10847 6690 10848
rect 11802 10912 12118 10913
rect 11802 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12118 10912
rect 11802 10847 12118 10848
rect 17230 10912 17546 10913
rect 17230 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17546 10912
rect 17230 10847 17546 10848
rect 22658 10912 22974 10913
rect 22658 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22974 10912
rect 22658 10847 22974 10848
rect 15193 10572 15259 10573
rect 15142 10508 15148 10572
rect 15212 10570 15259 10572
rect 15212 10568 15304 10570
rect 15254 10512 15304 10568
rect 15212 10510 15304 10512
rect 15212 10508 15259 10510
rect 15193 10507 15259 10508
rect 3660 10368 3976 10369
rect 3660 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3976 10368
rect 3660 10303 3976 10304
rect 9088 10368 9404 10369
rect 9088 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9404 10368
rect 9088 10303 9404 10304
rect 14516 10368 14832 10369
rect 14516 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14832 10368
rect 14516 10303 14832 10304
rect 19944 10368 20260 10369
rect 19944 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20260 10368
rect 19944 10303 20260 10304
rect 6374 9824 6690 9825
rect 6374 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6690 9824
rect 6374 9759 6690 9760
rect 11802 9824 12118 9825
rect 11802 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12118 9824
rect 11802 9759 12118 9760
rect 17230 9824 17546 9825
rect 17230 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17546 9824
rect 17230 9759 17546 9760
rect 22658 9824 22974 9825
rect 22658 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22974 9824
rect 22658 9759 22974 9760
rect 3660 9280 3976 9281
rect 3660 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3976 9280
rect 3660 9215 3976 9216
rect 9088 9280 9404 9281
rect 9088 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9404 9280
rect 9088 9215 9404 9216
rect 14516 9280 14832 9281
rect 14516 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14832 9280
rect 14516 9215 14832 9216
rect 19944 9280 20260 9281
rect 19944 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20260 9280
rect 19944 9215 20260 9216
rect 6374 8736 6690 8737
rect 6374 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6690 8736
rect 6374 8671 6690 8672
rect 11802 8736 12118 8737
rect 11802 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12118 8736
rect 11802 8671 12118 8672
rect 17230 8736 17546 8737
rect 17230 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17546 8736
rect 17230 8671 17546 8672
rect 22658 8736 22974 8737
rect 22658 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22974 8736
rect 22658 8671 22974 8672
rect 3660 8192 3976 8193
rect 3660 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3976 8192
rect 3660 8127 3976 8128
rect 9088 8192 9404 8193
rect 9088 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9404 8192
rect 9088 8127 9404 8128
rect 14516 8192 14832 8193
rect 14516 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14832 8192
rect 14516 8127 14832 8128
rect 19944 8192 20260 8193
rect 19944 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20260 8192
rect 19944 8127 20260 8128
rect 6374 7648 6690 7649
rect 6374 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6690 7648
rect 6374 7583 6690 7584
rect 11802 7648 12118 7649
rect 11802 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12118 7648
rect 11802 7583 12118 7584
rect 17230 7648 17546 7649
rect 17230 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17546 7648
rect 17230 7583 17546 7584
rect 22658 7648 22974 7649
rect 22658 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22974 7648
rect 22658 7583 22974 7584
rect 10225 7442 10291 7445
rect 17401 7442 17467 7445
rect 10225 7440 17467 7442
rect 10225 7384 10230 7440
rect 10286 7384 17406 7440
rect 17462 7384 17467 7440
rect 10225 7382 17467 7384
rect 10225 7379 10291 7382
rect 17401 7379 17467 7382
rect 3660 7104 3976 7105
rect 3660 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3976 7104
rect 3660 7039 3976 7040
rect 9088 7104 9404 7105
rect 9088 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9404 7104
rect 9088 7039 9404 7040
rect 14516 7104 14832 7105
rect 14516 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14832 7104
rect 14516 7039 14832 7040
rect 19944 7104 20260 7105
rect 19944 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20260 7104
rect 19944 7039 20260 7040
rect 11145 6762 11211 6765
rect 15142 6762 15148 6764
rect 11145 6760 15148 6762
rect 11145 6704 11150 6760
rect 11206 6704 15148 6760
rect 11145 6702 15148 6704
rect 11145 6699 11211 6702
rect 15142 6700 15148 6702
rect 15212 6700 15218 6764
rect 6374 6560 6690 6561
rect 6374 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6690 6560
rect 6374 6495 6690 6496
rect 11802 6560 12118 6561
rect 11802 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12118 6560
rect 11802 6495 12118 6496
rect 17230 6560 17546 6561
rect 17230 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17546 6560
rect 17230 6495 17546 6496
rect 22658 6560 22974 6561
rect 22658 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22974 6560
rect 22658 6495 22974 6496
rect 19609 6354 19675 6357
rect 19566 6352 19675 6354
rect 19566 6296 19614 6352
rect 19670 6296 19675 6352
rect 19566 6291 19675 6296
rect 3660 6016 3976 6017
rect 3660 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3976 6016
rect 3660 5951 3976 5952
rect 9088 6016 9404 6017
rect 9088 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9404 6016
rect 9088 5951 9404 5952
rect 14516 6016 14832 6017
rect 14516 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14832 6016
rect 14516 5951 14832 5952
rect 19425 5810 19491 5813
rect 19566 5810 19626 6291
rect 19944 6016 20260 6017
rect 19944 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20260 6016
rect 19944 5951 20260 5952
rect 19425 5808 19626 5810
rect 19425 5752 19430 5808
rect 19486 5752 19626 5808
rect 19425 5750 19626 5752
rect 19425 5747 19491 5750
rect 19609 5676 19675 5677
rect 19558 5612 19564 5676
rect 19628 5674 19675 5676
rect 19628 5672 19720 5674
rect 19670 5616 19720 5672
rect 19628 5614 19720 5616
rect 19628 5612 19675 5614
rect 19609 5611 19675 5612
rect 6374 5472 6690 5473
rect 6374 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6690 5472
rect 6374 5407 6690 5408
rect 11802 5472 12118 5473
rect 11802 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12118 5472
rect 11802 5407 12118 5408
rect 17230 5472 17546 5473
rect 17230 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17546 5472
rect 17230 5407 17546 5408
rect 22658 5472 22974 5473
rect 22658 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22974 5472
rect 22658 5407 22974 5408
rect 3660 4928 3976 4929
rect 3660 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3976 4928
rect 3660 4863 3976 4864
rect 9088 4928 9404 4929
rect 9088 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9404 4928
rect 9088 4863 9404 4864
rect 14516 4928 14832 4929
rect 14516 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14832 4928
rect 14516 4863 14832 4864
rect 19944 4928 20260 4929
rect 19944 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20260 4928
rect 19944 4863 20260 4864
rect 6374 4384 6690 4385
rect 6374 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6690 4384
rect 6374 4319 6690 4320
rect 11802 4384 12118 4385
rect 11802 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12118 4384
rect 11802 4319 12118 4320
rect 17230 4384 17546 4385
rect 17230 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17546 4384
rect 17230 4319 17546 4320
rect 22658 4384 22974 4385
rect 22658 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22974 4384
rect 22658 4319 22974 4320
rect 0 4042 800 4132
rect 4061 4042 4127 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3892 800 3982
rect 4061 3979 4127 3982
rect 13905 4042 13971 4045
rect 19057 4042 19123 4045
rect 19558 4042 19564 4044
rect 13905 4040 19564 4042
rect 13905 3984 13910 4040
rect 13966 3984 19062 4040
rect 19118 3984 19564 4040
rect 13905 3982 19564 3984
rect 13905 3979 13971 3982
rect 19057 3979 19123 3982
rect 19558 3980 19564 3982
rect 19628 3980 19634 4044
rect 3660 3840 3976 3841
rect 3660 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3976 3840
rect 3660 3775 3976 3776
rect 9088 3840 9404 3841
rect 9088 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9404 3840
rect 9088 3775 9404 3776
rect 14516 3840 14832 3841
rect 14516 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14832 3840
rect 14516 3775 14832 3776
rect 19944 3840 20260 3841
rect 19944 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20260 3840
rect 19944 3775 20260 3776
rect 6374 3296 6690 3297
rect 6374 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6690 3296
rect 6374 3231 6690 3232
rect 11802 3296 12118 3297
rect 11802 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12118 3296
rect 11802 3231 12118 3232
rect 17230 3296 17546 3297
rect 17230 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17546 3296
rect 17230 3231 17546 3232
rect 22658 3296 22974 3297
rect 22658 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22974 3296
rect 22658 3231 22974 3232
rect 3660 2752 3976 2753
rect 3660 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3976 2752
rect 3660 2687 3976 2688
rect 9088 2752 9404 2753
rect 9088 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9404 2752
rect 9088 2687 9404 2688
rect 14516 2752 14832 2753
rect 14516 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14832 2752
rect 14516 2687 14832 2688
rect 19944 2752 20260 2753
rect 19944 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20260 2752
rect 19944 2687 20260 2688
rect 6374 2208 6690 2209
rect 6374 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6690 2208
rect 6374 2143 6690 2144
rect 11802 2208 12118 2209
rect 11802 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12118 2208
rect 11802 2143 12118 2144
rect 17230 2208 17546 2209
rect 17230 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17546 2208
rect 17230 2143 17546 2144
rect 22658 2208 22974 2209
rect 22658 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22974 2208
rect 22658 2143 22974 2144
<< via3 >>
rect 6380 21788 6444 21792
rect 6380 21732 6384 21788
rect 6384 21732 6440 21788
rect 6440 21732 6444 21788
rect 6380 21728 6444 21732
rect 6460 21788 6524 21792
rect 6460 21732 6464 21788
rect 6464 21732 6520 21788
rect 6520 21732 6524 21788
rect 6460 21728 6524 21732
rect 6540 21788 6604 21792
rect 6540 21732 6544 21788
rect 6544 21732 6600 21788
rect 6600 21732 6604 21788
rect 6540 21728 6604 21732
rect 6620 21788 6684 21792
rect 6620 21732 6624 21788
rect 6624 21732 6680 21788
rect 6680 21732 6684 21788
rect 6620 21728 6684 21732
rect 11808 21788 11872 21792
rect 11808 21732 11812 21788
rect 11812 21732 11868 21788
rect 11868 21732 11872 21788
rect 11808 21728 11872 21732
rect 11888 21788 11952 21792
rect 11888 21732 11892 21788
rect 11892 21732 11948 21788
rect 11948 21732 11952 21788
rect 11888 21728 11952 21732
rect 11968 21788 12032 21792
rect 11968 21732 11972 21788
rect 11972 21732 12028 21788
rect 12028 21732 12032 21788
rect 11968 21728 12032 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 17316 21788 17380 21792
rect 17316 21732 17320 21788
rect 17320 21732 17376 21788
rect 17376 21732 17380 21788
rect 17316 21728 17380 21732
rect 17396 21788 17460 21792
rect 17396 21732 17400 21788
rect 17400 21732 17456 21788
rect 17456 21732 17460 21788
rect 17396 21728 17460 21732
rect 17476 21788 17540 21792
rect 17476 21732 17480 21788
rect 17480 21732 17536 21788
rect 17536 21732 17540 21788
rect 17476 21728 17540 21732
rect 22664 21788 22728 21792
rect 22664 21732 22668 21788
rect 22668 21732 22724 21788
rect 22724 21732 22728 21788
rect 22664 21728 22728 21732
rect 22744 21788 22808 21792
rect 22744 21732 22748 21788
rect 22748 21732 22804 21788
rect 22804 21732 22808 21788
rect 22744 21728 22808 21732
rect 22824 21788 22888 21792
rect 22824 21732 22828 21788
rect 22828 21732 22884 21788
rect 22884 21732 22888 21788
rect 22824 21728 22888 21732
rect 22904 21788 22968 21792
rect 22904 21732 22908 21788
rect 22908 21732 22964 21788
rect 22964 21732 22968 21788
rect 22904 21728 22968 21732
rect 3666 21244 3730 21248
rect 3666 21188 3670 21244
rect 3670 21188 3726 21244
rect 3726 21188 3730 21244
rect 3666 21184 3730 21188
rect 3746 21244 3810 21248
rect 3746 21188 3750 21244
rect 3750 21188 3806 21244
rect 3806 21188 3810 21244
rect 3746 21184 3810 21188
rect 3826 21244 3890 21248
rect 3826 21188 3830 21244
rect 3830 21188 3886 21244
rect 3886 21188 3890 21244
rect 3826 21184 3890 21188
rect 3906 21244 3970 21248
rect 3906 21188 3910 21244
rect 3910 21188 3966 21244
rect 3966 21188 3970 21244
rect 3906 21184 3970 21188
rect 9094 21244 9158 21248
rect 9094 21188 9098 21244
rect 9098 21188 9154 21244
rect 9154 21188 9158 21244
rect 9094 21184 9158 21188
rect 9174 21244 9238 21248
rect 9174 21188 9178 21244
rect 9178 21188 9234 21244
rect 9234 21188 9238 21244
rect 9174 21184 9238 21188
rect 9254 21244 9318 21248
rect 9254 21188 9258 21244
rect 9258 21188 9314 21244
rect 9314 21188 9318 21244
rect 9254 21184 9318 21188
rect 9334 21244 9398 21248
rect 9334 21188 9338 21244
rect 9338 21188 9394 21244
rect 9394 21188 9398 21244
rect 9334 21184 9398 21188
rect 14522 21244 14586 21248
rect 14522 21188 14526 21244
rect 14526 21188 14582 21244
rect 14582 21188 14586 21244
rect 14522 21184 14586 21188
rect 14602 21244 14666 21248
rect 14602 21188 14606 21244
rect 14606 21188 14662 21244
rect 14662 21188 14666 21244
rect 14602 21184 14666 21188
rect 14682 21244 14746 21248
rect 14682 21188 14686 21244
rect 14686 21188 14742 21244
rect 14742 21188 14746 21244
rect 14682 21184 14746 21188
rect 14762 21244 14826 21248
rect 14762 21188 14766 21244
rect 14766 21188 14822 21244
rect 14822 21188 14826 21244
rect 14762 21184 14826 21188
rect 19950 21244 20014 21248
rect 19950 21188 19954 21244
rect 19954 21188 20010 21244
rect 20010 21188 20014 21244
rect 19950 21184 20014 21188
rect 20030 21244 20094 21248
rect 20030 21188 20034 21244
rect 20034 21188 20090 21244
rect 20090 21188 20094 21244
rect 20030 21184 20094 21188
rect 20110 21244 20174 21248
rect 20110 21188 20114 21244
rect 20114 21188 20170 21244
rect 20170 21188 20174 21244
rect 20110 21184 20174 21188
rect 20190 21244 20254 21248
rect 20190 21188 20194 21244
rect 20194 21188 20250 21244
rect 20250 21188 20254 21244
rect 20190 21184 20254 21188
rect 6380 20700 6444 20704
rect 6380 20644 6384 20700
rect 6384 20644 6440 20700
rect 6440 20644 6444 20700
rect 6380 20640 6444 20644
rect 6460 20700 6524 20704
rect 6460 20644 6464 20700
rect 6464 20644 6520 20700
rect 6520 20644 6524 20700
rect 6460 20640 6524 20644
rect 6540 20700 6604 20704
rect 6540 20644 6544 20700
rect 6544 20644 6600 20700
rect 6600 20644 6604 20700
rect 6540 20640 6604 20644
rect 6620 20700 6684 20704
rect 6620 20644 6624 20700
rect 6624 20644 6680 20700
rect 6680 20644 6684 20700
rect 6620 20640 6684 20644
rect 11808 20700 11872 20704
rect 11808 20644 11812 20700
rect 11812 20644 11868 20700
rect 11868 20644 11872 20700
rect 11808 20640 11872 20644
rect 11888 20700 11952 20704
rect 11888 20644 11892 20700
rect 11892 20644 11948 20700
rect 11948 20644 11952 20700
rect 11888 20640 11952 20644
rect 11968 20700 12032 20704
rect 11968 20644 11972 20700
rect 11972 20644 12028 20700
rect 12028 20644 12032 20700
rect 11968 20640 12032 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 17316 20700 17380 20704
rect 17316 20644 17320 20700
rect 17320 20644 17376 20700
rect 17376 20644 17380 20700
rect 17316 20640 17380 20644
rect 17396 20700 17460 20704
rect 17396 20644 17400 20700
rect 17400 20644 17456 20700
rect 17456 20644 17460 20700
rect 17396 20640 17460 20644
rect 17476 20700 17540 20704
rect 17476 20644 17480 20700
rect 17480 20644 17536 20700
rect 17536 20644 17540 20700
rect 17476 20640 17540 20644
rect 22664 20700 22728 20704
rect 22664 20644 22668 20700
rect 22668 20644 22724 20700
rect 22724 20644 22728 20700
rect 22664 20640 22728 20644
rect 22744 20700 22808 20704
rect 22744 20644 22748 20700
rect 22748 20644 22804 20700
rect 22804 20644 22808 20700
rect 22744 20640 22808 20644
rect 22824 20700 22888 20704
rect 22824 20644 22828 20700
rect 22828 20644 22884 20700
rect 22884 20644 22888 20700
rect 22824 20640 22888 20644
rect 22904 20700 22968 20704
rect 22904 20644 22908 20700
rect 22908 20644 22964 20700
rect 22964 20644 22968 20700
rect 22904 20640 22968 20644
rect 3666 20156 3730 20160
rect 3666 20100 3670 20156
rect 3670 20100 3726 20156
rect 3726 20100 3730 20156
rect 3666 20096 3730 20100
rect 3746 20156 3810 20160
rect 3746 20100 3750 20156
rect 3750 20100 3806 20156
rect 3806 20100 3810 20156
rect 3746 20096 3810 20100
rect 3826 20156 3890 20160
rect 3826 20100 3830 20156
rect 3830 20100 3886 20156
rect 3886 20100 3890 20156
rect 3826 20096 3890 20100
rect 3906 20156 3970 20160
rect 3906 20100 3910 20156
rect 3910 20100 3966 20156
rect 3966 20100 3970 20156
rect 3906 20096 3970 20100
rect 9094 20156 9158 20160
rect 9094 20100 9098 20156
rect 9098 20100 9154 20156
rect 9154 20100 9158 20156
rect 9094 20096 9158 20100
rect 9174 20156 9238 20160
rect 9174 20100 9178 20156
rect 9178 20100 9234 20156
rect 9234 20100 9238 20156
rect 9174 20096 9238 20100
rect 9254 20156 9318 20160
rect 9254 20100 9258 20156
rect 9258 20100 9314 20156
rect 9314 20100 9318 20156
rect 9254 20096 9318 20100
rect 9334 20156 9398 20160
rect 9334 20100 9338 20156
rect 9338 20100 9394 20156
rect 9394 20100 9398 20156
rect 9334 20096 9398 20100
rect 14522 20156 14586 20160
rect 14522 20100 14526 20156
rect 14526 20100 14582 20156
rect 14582 20100 14586 20156
rect 14522 20096 14586 20100
rect 14602 20156 14666 20160
rect 14602 20100 14606 20156
rect 14606 20100 14662 20156
rect 14662 20100 14666 20156
rect 14602 20096 14666 20100
rect 14682 20156 14746 20160
rect 14682 20100 14686 20156
rect 14686 20100 14742 20156
rect 14742 20100 14746 20156
rect 14682 20096 14746 20100
rect 14762 20156 14826 20160
rect 14762 20100 14766 20156
rect 14766 20100 14822 20156
rect 14822 20100 14826 20156
rect 14762 20096 14826 20100
rect 19950 20156 20014 20160
rect 19950 20100 19954 20156
rect 19954 20100 20010 20156
rect 20010 20100 20014 20156
rect 19950 20096 20014 20100
rect 20030 20156 20094 20160
rect 20030 20100 20034 20156
rect 20034 20100 20090 20156
rect 20090 20100 20094 20156
rect 20030 20096 20094 20100
rect 20110 20156 20174 20160
rect 20110 20100 20114 20156
rect 20114 20100 20170 20156
rect 20170 20100 20174 20156
rect 20110 20096 20174 20100
rect 20190 20156 20254 20160
rect 20190 20100 20194 20156
rect 20194 20100 20250 20156
rect 20250 20100 20254 20156
rect 20190 20096 20254 20100
rect 6380 19612 6444 19616
rect 6380 19556 6384 19612
rect 6384 19556 6440 19612
rect 6440 19556 6444 19612
rect 6380 19552 6444 19556
rect 6460 19612 6524 19616
rect 6460 19556 6464 19612
rect 6464 19556 6520 19612
rect 6520 19556 6524 19612
rect 6460 19552 6524 19556
rect 6540 19612 6604 19616
rect 6540 19556 6544 19612
rect 6544 19556 6600 19612
rect 6600 19556 6604 19612
rect 6540 19552 6604 19556
rect 6620 19612 6684 19616
rect 6620 19556 6624 19612
rect 6624 19556 6680 19612
rect 6680 19556 6684 19612
rect 6620 19552 6684 19556
rect 11808 19612 11872 19616
rect 11808 19556 11812 19612
rect 11812 19556 11868 19612
rect 11868 19556 11872 19612
rect 11808 19552 11872 19556
rect 11888 19612 11952 19616
rect 11888 19556 11892 19612
rect 11892 19556 11948 19612
rect 11948 19556 11952 19612
rect 11888 19552 11952 19556
rect 11968 19612 12032 19616
rect 11968 19556 11972 19612
rect 11972 19556 12028 19612
rect 12028 19556 12032 19612
rect 11968 19552 12032 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 17316 19612 17380 19616
rect 17316 19556 17320 19612
rect 17320 19556 17376 19612
rect 17376 19556 17380 19612
rect 17316 19552 17380 19556
rect 17396 19612 17460 19616
rect 17396 19556 17400 19612
rect 17400 19556 17456 19612
rect 17456 19556 17460 19612
rect 17396 19552 17460 19556
rect 17476 19612 17540 19616
rect 17476 19556 17480 19612
rect 17480 19556 17536 19612
rect 17536 19556 17540 19612
rect 17476 19552 17540 19556
rect 22664 19612 22728 19616
rect 22664 19556 22668 19612
rect 22668 19556 22724 19612
rect 22724 19556 22728 19612
rect 22664 19552 22728 19556
rect 22744 19612 22808 19616
rect 22744 19556 22748 19612
rect 22748 19556 22804 19612
rect 22804 19556 22808 19612
rect 22744 19552 22808 19556
rect 22824 19612 22888 19616
rect 22824 19556 22828 19612
rect 22828 19556 22884 19612
rect 22884 19556 22888 19612
rect 22824 19552 22888 19556
rect 22904 19612 22968 19616
rect 22904 19556 22908 19612
rect 22908 19556 22964 19612
rect 22964 19556 22968 19612
rect 22904 19552 22968 19556
rect 3666 19068 3730 19072
rect 3666 19012 3670 19068
rect 3670 19012 3726 19068
rect 3726 19012 3730 19068
rect 3666 19008 3730 19012
rect 3746 19068 3810 19072
rect 3746 19012 3750 19068
rect 3750 19012 3806 19068
rect 3806 19012 3810 19068
rect 3746 19008 3810 19012
rect 3826 19068 3890 19072
rect 3826 19012 3830 19068
rect 3830 19012 3886 19068
rect 3886 19012 3890 19068
rect 3826 19008 3890 19012
rect 3906 19068 3970 19072
rect 3906 19012 3910 19068
rect 3910 19012 3966 19068
rect 3966 19012 3970 19068
rect 3906 19008 3970 19012
rect 9094 19068 9158 19072
rect 9094 19012 9098 19068
rect 9098 19012 9154 19068
rect 9154 19012 9158 19068
rect 9094 19008 9158 19012
rect 9174 19068 9238 19072
rect 9174 19012 9178 19068
rect 9178 19012 9234 19068
rect 9234 19012 9238 19068
rect 9174 19008 9238 19012
rect 9254 19068 9318 19072
rect 9254 19012 9258 19068
rect 9258 19012 9314 19068
rect 9314 19012 9318 19068
rect 9254 19008 9318 19012
rect 9334 19068 9398 19072
rect 9334 19012 9338 19068
rect 9338 19012 9394 19068
rect 9394 19012 9398 19068
rect 9334 19008 9398 19012
rect 14522 19068 14586 19072
rect 14522 19012 14526 19068
rect 14526 19012 14582 19068
rect 14582 19012 14586 19068
rect 14522 19008 14586 19012
rect 14602 19068 14666 19072
rect 14602 19012 14606 19068
rect 14606 19012 14662 19068
rect 14662 19012 14666 19068
rect 14602 19008 14666 19012
rect 14682 19068 14746 19072
rect 14682 19012 14686 19068
rect 14686 19012 14742 19068
rect 14742 19012 14746 19068
rect 14682 19008 14746 19012
rect 14762 19068 14826 19072
rect 14762 19012 14766 19068
rect 14766 19012 14822 19068
rect 14822 19012 14826 19068
rect 14762 19008 14826 19012
rect 19950 19068 20014 19072
rect 19950 19012 19954 19068
rect 19954 19012 20010 19068
rect 20010 19012 20014 19068
rect 19950 19008 20014 19012
rect 20030 19068 20094 19072
rect 20030 19012 20034 19068
rect 20034 19012 20090 19068
rect 20090 19012 20094 19068
rect 20030 19008 20094 19012
rect 20110 19068 20174 19072
rect 20110 19012 20114 19068
rect 20114 19012 20170 19068
rect 20170 19012 20174 19068
rect 20110 19008 20174 19012
rect 20190 19068 20254 19072
rect 20190 19012 20194 19068
rect 20194 19012 20250 19068
rect 20250 19012 20254 19068
rect 20190 19008 20254 19012
rect 6380 18524 6444 18528
rect 6380 18468 6384 18524
rect 6384 18468 6440 18524
rect 6440 18468 6444 18524
rect 6380 18464 6444 18468
rect 6460 18524 6524 18528
rect 6460 18468 6464 18524
rect 6464 18468 6520 18524
rect 6520 18468 6524 18524
rect 6460 18464 6524 18468
rect 6540 18524 6604 18528
rect 6540 18468 6544 18524
rect 6544 18468 6600 18524
rect 6600 18468 6604 18524
rect 6540 18464 6604 18468
rect 6620 18524 6684 18528
rect 6620 18468 6624 18524
rect 6624 18468 6680 18524
rect 6680 18468 6684 18524
rect 6620 18464 6684 18468
rect 11808 18524 11872 18528
rect 11808 18468 11812 18524
rect 11812 18468 11868 18524
rect 11868 18468 11872 18524
rect 11808 18464 11872 18468
rect 11888 18524 11952 18528
rect 11888 18468 11892 18524
rect 11892 18468 11948 18524
rect 11948 18468 11952 18524
rect 11888 18464 11952 18468
rect 11968 18524 12032 18528
rect 11968 18468 11972 18524
rect 11972 18468 12028 18524
rect 12028 18468 12032 18524
rect 11968 18464 12032 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 17316 18524 17380 18528
rect 17316 18468 17320 18524
rect 17320 18468 17376 18524
rect 17376 18468 17380 18524
rect 17316 18464 17380 18468
rect 17396 18524 17460 18528
rect 17396 18468 17400 18524
rect 17400 18468 17456 18524
rect 17456 18468 17460 18524
rect 17396 18464 17460 18468
rect 17476 18524 17540 18528
rect 17476 18468 17480 18524
rect 17480 18468 17536 18524
rect 17536 18468 17540 18524
rect 17476 18464 17540 18468
rect 22664 18524 22728 18528
rect 22664 18468 22668 18524
rect 22668 18468 22724 18524
rect 22724 18468 22728 18524
rect 22664 18464 22728 18468
rect 22744 18524 22808 18528
rect 22744 18468 22748 18524
rect 22748 18468 22804 18524
rect 22804 18468 22808 18524
rect 22744 18464 22808 18468
rect 22824 18524 22888 18528
rect 22824 18468 22828 18524
rect 22828 18468 22884 18524
rect 22884 18468 22888 18524
rect 22824 18464 22888 18468
rect 22904 18524 22968 18528
rect 22904 18468 22908 18524
rect 22908 18468 22964 18524
rect 22964 18468 22968 18524
rect 22904 18464 22968 18468
rect 3666 17980 3730 17984
rect 3666 17924 3670 17980
rect 3670 17924 3726 17980
rect 3726 17924 3730 17980
rect 3666 17920 3730 17924
rect 3746 17980 3810 17984
rect 3746 17924 3750 17980
rect 3750 17924 3806 17980
rect 3806 17924 3810 17980
rect 3746 17920 3810 17924
rect 3826 17980 3890 17984
rect 3826 17924 3830 17980
rect 3830 17924 3886 17980
rect 3886 17924 3890 17980
rect 3826 17920 3890 17924
rect 3906 17980 3970 17984
rect 3906 17924 3910 17980
rect 3910 17924 3966 17980
rect 3966 17924 3970 17980
rect 3906 17920 3970 17924
rect 9094 17980 9158 17984
rect 9094 17924 9098 17980
rect 9098 17924 9154 17980
rect 9154 17924 9158 17980
rect 9094 17920 9158 17924
rect 9174 17980 9238 17984
rect 9174 17924 9178 17980
rect 9178 17924 9234 17980
rect 9234 17924 9238 17980
rect 9174 17920 9238 17924
rect 9254 17980 9318 17984
rect 9254 17924 9258 17980
rect 9258 17924 9314 17980
rect 9314 17924 9318 17980
rect 9254 17920 9318 17924
rect 9334 17980 9398 17984
rect 9334 17924 9338 17980
rect 9338 17924 9394 17980
rect 9394 17924 9398 17980
rect 9334 17920 9398 17924
rect 14522 17980 14586 17984
rect 14522 17924 14526 17980
rect 14526 17924 14582 17980
rect 14582 17924 14586 17980
rect 14522 17920 14586 17924
rect 14602 17980 14666 17984
rect 14602 17924 14606 17980
rect 14606 17924 14662 17980
rect 14662 17924 14666 17980
rect 14602 17920 14666 17924
rect 14682 17980 14746 17984
rect 14682 17924 14686 17980
rect 14686 17924 14742 17980
rect 14742 17924 14746 17980
rect 14682 17920 14746 17924
rect 14762 17980 14826 17984
rect 14762 17924 14766 17980
rect 14766 17924 14822 17980
rect 14822 17924 14826 17980
rect 14762 17920 14826 17924
rect 19950 17980 20014 17984
rect 19950 17924 19954 17980
rect 19954 17924 20010 17980
rect 20010 17924 20014 17980
rect 19950 17920 20014 17924
rect 20030 17980 20094 17984
rect 20030 17924 20034 17980
rect 20034 17924 20090 17980
rect 20090 17924 20094 17980
rect 20030 17920 20094 17924
rect 20110 17980 20174 17984
rect 20110 17924 20114 17980
rect 20114 17924 20170 17980
rect 20170 17924 20174 17980
rect 20110 17920 20174 17924
rect 20190 17980 20254 17984
rect 20190 17924 20194 17980
rect 20194 17924 20250 17980
rect 20250 17924 20254 17980
rect 20190 17920 20254 17924
rect 6380 17436 6444 17440
rect 6380 17380 6384 17436
rect 6384 17380 6440 17436
rect 6440 17380 6444 17436
rect 6380 17376 6444 17380
rect 6460 17436 6524 17440
rect 6460 17380 6464 17436
rect 6464 17380 6520 17436
rect 6520 17380 6524 17436
rect 6460 17376 6524 17380
rect 6540 17436 6604 17440
rect 6540 17380 6544 17436
rect 6544 17380 6600 17436
rect 6600 17380 6604 17436
rect 6540 17376 6604 17380
rect 6620 17436 6684 17440
rect 6620 17380 6624 17436
rect 6624 17380 6680 17436
rect 6680 17380 6684 17436
rect 6620 17376 6684 17380
rect 11808 17436 11872 17440
rect 11808 17380 11812 17436
rect 11812 17380 11868 17436
rect 11868 17380 11872 17436
rect 11808 17376 11872 17380
rect 11888 17436 11952 17440
rect 11888 17380 11892 17436
rect 11892 17380 11948 17436
rect 11948 17380 11952 17436
rect 11888 17376 11952 17380
rect 11968 17436 12032 17440
rect 11968 17380 11972 17436
rect 11972 17380 12028 17436
rect 12028 17380 12032 17436
rect 11968 17376 12032 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 17316 17436 17380 17440
rect 17316 17380 17320 17436
rect 17320 17380 17376 17436
rect 17376 17380 17380 17436
rect 17316 17376 17380 17380
rect 17396 17436 17460 17440
rect 17396 17380 17400 17436
rect 17400 17380 17456 17436
rect 17456 17380 17460 17436
rect 17396 17376 17460 17380
rect 17476 17436 17540 17440
rect 17476 17380 17480 17436
rect 17480 17380 17536 17436
rect 17536 17380 17540 17436
rect 17476 17376 17540 17380
rect 22664 17436 22728 17440
rect 22664 17380 22668 17436
rect 22668 17380 22724 17436
rect 22724 17380 22728 17436
rect 22664 17376 22728 17380
rect 22744 17436 22808 17440
rect 22744 17380 22748 17436
rect 22748 17380 22804 17436
rect 22804 17380 22808 17436
rect 22744 17376 22808 17380
rect 22824 17436 22888 17440
rect 22824 17380 22828 17436
rect 22828 17380 22884 17436
rect 22884 17380 22888 17436
rect 22824 17376 22888 17380
rect 22904 17436 22968 17440
rect 22904 17380 22908 17436
rect 22908 17380 22964 17436
rect 22964 17380 22968 17436
rect 22904 17376 22968 17380
rect 3666 16892 3730 16896
rect 3666 16836 3670 16892
rect 3670 16836 3726 16892
rect 3726 16836 3730 16892
rect 3666 16832 3730 16836
rect 3746 16892 3810 16896
rect 3746 16836 3750 16892
rect 3750 16836 3806 16892
rect 3806 16836 3810 16892
rect 3746 16832 3810 16836
rect 3826 16892 3890 16896
rect 3826 16836 3830 16892
rect 3830 16836 3886 16892
rect 3886 16836 3890 16892
rect 3826 16832 3890 16836
rect 3906 16892 3970 16896
rect 3906 16836 3910 16892
rect 3910 16836 3966 16892
rect 3966 16836 3970 16892
rect 3906 16832 3970 16836
rect 9094 16892 9158 16896
rect 9094 16836 9098 16892
rect 9098 16836 9154 16892
rect 9154 16836 9158 16892
rect 9094 16832 9158 16836
rect 9174 16892 9238 16896
rect 9174 16836 9178 16892
rect 9178 16836 9234 16892
rect 9234 16836 9238 16892
rect 9174 16832 9238 16836
rect 9254 16892 9318 16896
rect 9254 16836 9258 16892
rect 9258 16836 9314 16892
rect 9314 16836 9318 16892
rect 9254 16832 9318 16836
rect 9334 16892 9398 16896
rect 9334 16836 9338 16892
rect 9338 16836 9394 16892
rect 9394 16836 9398 16892
rect 9334 16832 9398 16836
rect 14522 16892 14586 16896
rect 14522 16836 14526 16892
rect 14526 16836 14582 16892
rect 14582 16836 14586 16892
rect 14522 16832 14586 16836
rect 14602 16892 14666 16896
rect 14602 16836 14606 16892
rect 14606 16836 14662 16892
rect 14662 16836 14666 16892
rect 14602 16832 14666 16836
rect 14682 16892 14746 16896
rect 14682 16836 14686 16892
rect 14686 16836 14742 16892
rect 14742 16836 14746 16892
rect 14682 16832 14746 16836
rect 14762 16892 14826 16896
rect 14762 16836 14766 16892
rect 14766 16836 14822 16892
rect 14822 16836 14826 16892
rect 14762 16832 14826 16836
rect 19950 16892 20014 16896
rect 19950 16836 19954 16892
rect 19954 16836 20010 16892
rect 20010 16836 20014 16892
rect 19950 16832 20014 16836
rect 20030 16892 20094 16896
rect 20030 16836 20034 16892
rect 20034 16836 20090 16892
rect 20090 16836 20094 16892
rect 20030 16832 20094 16836
rect 20110 16892 20174 16896
rect 20110 16836 20114 16892
rect 20114 16836 20170 16892
rect 20170 16836 20174 16892
rect 20110 16832 20174 16836
rect 20190 16892 20254 16896
rect 20190 16836 20194 16892
rect 20194 16836 20250 16892
rect 20250 16836 20254 16892
rect 20190 16832 20254 16836
rect 6380 16348 6444 16352
rect 6380 16292 6384 16348
rect 6384 16292 6440 16348
rect 6440 16292 6444 16348
rect 6380 16288 6444 16292
rect 6460 16348 6524 16352
rect 6460 16292 6464 16348
rect 6464 16292 6520 16348
rect 6520 16292 6524 16348
rect 6460 16288 6524 16292
rect 6540 16348 6604 16352
rect 6540 16292 6544 16348
rect 6544 16292 6600 16348
rect 6600 16292 6604 16348
rect 6540 16288 6604 16292
rect 6620 16348 6684 16352
rect 6620 16292 6624 16348
rect 6624 16292 6680 16348
rect 6680 16292 6684 16348
rect 6620 16288 6684 16292
rect 11808 16348 11872 16352
rect 11808 16292 11812 16348
rect 11812 16292 11868 16348
rect 11868 16292 11872 16348
rect 11808 16288 11872 16292
rect 11888 16348 11952 16352
rect 11888 16292 11892 16348
rect 11892 16292 11948 16348
rect 11948 16292 11952 16348
rect 11888 16288 11952 16292
rect 11968 16348 12032 16352
rect 11968 16292 11972 16348
rect 11972 16292 12028 16348
rect 12028 16292 12032 16348
rect 11968 16288 12032 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 17316 16348 17380 16352
rect 17316 16292 17320 16348
rect 17320 16292 17376 16348
rect 17376 16292 17380 16348
rect 17316 16288 17380 16292
rect 17396 16348 17460 16352
rect 17396 16292 17400 16348
rect 17400 16292 17456 16348
rect 17456 16292 17460 16348
rect 17396 16288 17460 16292
rect 17476 16348 17540 16352
rect 17476 16292 17480 16348
rect 17480 16292 17536 16348
rect 17536 16292 17540 16348
rect 17476 16288 17540 16292
rect 22664 16348 22728 16352
rect 22664 16292 22668 16348
rect 22668 16292 22724 16348
rect 22724 16292 22728 16348
rect 22664 16288 22728 16292
rect 22744 16348 22808 16352
rect 22744 16292 22748 16348
rect 22748 16292 22804 16348
rect 22804 16292 22808 16348
rect 22744 16288 22808 16292
rect 22824 16348 22888 16352
rect 22824 16292 22828 16348
rect 22828 16292 22884 16348
rect 22884 16292 22888 16348
rect 22824 16288 22888 16292
rect 22904 16348 22968 16352
rect 22904 16292 22908 16348
rect 22908 16292 22964 16348
rect 22964 16292 22968 16348
rect 22904 16288 22968 16292
rect 3666 15804 3730 15808
rect 3666 15748 3670 15804
rect 3670 15748 3726 15804
rect 3726 15748 3730 15804
rect 3666 15744 3730 15748
rect 3746 15804 3810 15808
rect 3746 15748 3750 15804
rect 3750 15748 3806 15804
rect 3806 15748 3810 15804
rect 3746 15744 3810 15748
rect 3826 15804 3890 15808
rect 3826 15748 3830 15804
rect 3830 15748 3886 15804
rect 3886 15748 3890 15804
rect 3826 15744 3890 15748
rect 3906 15804 3970 15808
rect 3906 15748 3910 15804
rect 3910 15748 3966 15804
rect 3966 15748 3970 15804
rect 3906 15744 3970 15748
rect 9094 15804 9158 15808
rect 9094 15748 9098 15804
rect 9098 15748 9154 15804
rect 9154 15748 9158 15804
rect 9094 15744 9158 15748
rect 9174 15804 9238 15808
rect 9174 15748 9178 15804
rect 9178 15748 9234 15804
rect 9234 15748 9238 15804
rect 9174 15744 9238 15748
rect 9254 15804 9318 15808
rect 9254 15748 9258 15804
rect 9258 15748 9314 15804
rect 9314 15748 9318 15804
rect 9254 15744 9318 15748
rect 9334 15804 9398 15808
rect 9334 15748 9338 15804
rect 9338 15748 9394 15804
rect 9394 15748 9398 15804
rect 9334 15744 9398 15748
rect 14522 15804 14586 15808
rect 14522 15748 14526 15804
rect 14526 15748 14582 15804
rect 14582 15748 14586 15804
rect 14522 15744 14586 15748
rect 14602 15804 14666 15808
rect 14602 15748 14606 15804
rect 14606 15748 14662 15804
rect 14662 15748 14666 15804
rect 14602 15744 14666 15748
rect 14682 15804 14746 15808
rect 14682 15748 14686 15804
rect 14686 15748 14742 15804
rect 14742 15748 14746 15804
rect 14682 15744 14746 15748
rect 14762 15804 14826 15808
rect 14762 15748 14766 15804
rect 14766 15748 14822 15804
rect 14822 15748 14826 15804
rect 14762 15744 14826 15748
rect 19950 15804 20014 15808
rect 19950 15748 19954 15804
rect 19954 15748 20010 15804
rect 20010 15748 20014 15804
rect 19950 15744 20014 15748
rect 20030 15804 20094 15808
rect 20030 15748 20034 15804
rect 20034 15748 20090 15804
rect 20090 15748 20094 15804
rect 20030 15744 20094 15748
rect 20110 15804 20174 15808
rect 20110 15748 20114 15804
rect 20114 15748 20170 15804
rect 20170 15748 20174 15804
rect 20110 15744 20174 15748
rect 20190 15804 20254 15808
rect 20190 15748 20194 15804
rect 20194 15748 20250 15804
rect 20250 15748 20254 15804
rect 20190 15744 20254 15748
rect 6380 15260 6444 15264
rect 6380 15204 6384 15260
rect 6384 15204 6440 15260
rect 6440 15204 6444 15260
rect 6380 15200 6444 15204
rect 6460 15260 6524 15264
rect 6460 15204 6464 15260
rect 6464 15204 6520 15260
rect 6520 15204 6524 15260
rect 6460 15200 6524 15204
rect 6540 15260 6604 15264
rect 6540 15204 6544 15260
rect 6544 15204 6600 15260
rect 6600 15204 6604 15260
rect 6540 15200 6604 15204
rect 6620 15260 6684 15264
rect 6620 15204 6624 15260
rect 6624 15204 6680 15260
rect 6680 15204 6684 15260
rect 6620 15200 6684 15204
rect 11808 15260 11872 15264
rect 11808 15204 11812 15260
rect 11812 15204 11868 15260
rect 11868 15204 11872 15260
rect 11808 15200 11872 15204
rect 11888 15260 11952 15264
rect 11888 15204 11892 15260
rect 11892 15204 11948 15260
rect 11948 15204 11952 15260
rect 11888 15200 11952 15204
rect 11968 15260 12032 15264
rect 11968 15204 11972 15260
rect 11972 15204 12028 15260
rect 12028 15204 12032 15260
rect 11968 15200 12032 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 17316 15260 17380 15264
rect 17316 15204 17320 15260
rect 17320 15204 17376 15260
rect 17376 15204 17380 15260
rect 17316 15200 17380 15204
rect 17396 15260 17460 15264
rect 17396 15204 17400 15260
rect 17400 15204 17456 15260
rect 17456 15204 17460 15260
rect 17396 15200 17460 15204
rect 17476 15260 17540 15264
rect 17476 15204 17480 15260
rect 17480 15204 17536 15260
rect 17536 15204 17540 15260
rect 17476 15200 17540 15204
rect 22664 15260 22728 15264
rect 22664 15204 22668 15260
rect 22668 15204 22724 15260
rect 22724 15204 22728 15260
rect 22664 15200 22728 15204
rect 22744 15260 22808 15264
rect 22744 15204 22748 15260
rect 22748 15204 22804 15260
rect 22804 15204 22808 15260
rect 22744 15200 22808 15204
rect 22824 15260 22888 15264
rect 22824 15204 22828 15260
rect 22828 15204 22884 15260
rect 22884 15204 22888 15260
rect 22824 15200 22888 15204
rect 22904 15260 22968 15264
rect 22904 15204 22908 15260
rect 22908 15204 22964 15260
rect 22964 15204 22968 15260
rect 22904 15200 22968 15204
rect 3666 14716 3730 14720
rect 3666 14660 3670 14716
rect 3670 14660 3726 14716
rect 3726 14660 3730 14716
rect 3666 14656 3730 14660
rect 3746 14716 3810 14720
rect 3746 14660 3750 14716
rect 3750 14660 3806 14716
rect 3806 14660 3810 14716
rect 3746 14656 3810 14660
rect 3826 14716 3890 14720
rect 3826 14660 3830 14716
rect 3830 14660 3886 14716
rect 3886 14660 3890 14716
rect 3826 14656 3890 14660
rect 3906 14716 3970 14720
rect 3906 14660 3910 14716
rect 3910 14660 3966 14716
rect 3966 14660 3970 14716
rect 3906 14656 3970 14660
rect 9094 14716 9158 14720
rect 9094 14660 9098 14716
rect 9098 14660 9154 14716
rect 9154 14660 9158 14716
rect 9094 14656 9158 14660
rect 9174 14716 9238 14720
rect 9174 14660 9178 14716
rect 9178 14660 9234 14716
rect 9234 14660 9238 14716
rect 9174 14656 9238 14660
rect 9254 14716 9318 14720
rect 9254 14660 9258 14716
rect 9258 14660 9314 14716
rect 9314 14660 9318 14716
rect 9254 14656 9318 14660
rect 9334 14716 9398 14720
rect 9334 14660 9338 14716
rect 9338 14660 9394 14716
rect 9394 14660 9398 14716
rect 9334 14656 9398 14660
rect 14522 14716 14586 14720
rect 14522 14660 14526 14716
rect 14526 14660 14582 14716
rect 14582 14660 14586 14716
rect 14522 14656 14586 14660
rect 14602 14716 14666 14720
rect 14602 14660 14606 14716
rect 14606 14660 14662 14716
rect 14662 14660 14666 14716
rect 14602 14656 14666 14660
rect 14682 14716 14746 14720
rect 14682 14660 14686 14716
rect 14686 14660 14742 14716
rect 14742 14660 14746 14716
rect 14682 14656 14746 14660
rect 14762 14716 14826 14720
rect 14762 14660 14766 14716
rect 14766 14660 14822 14716
rect 14822 14660 14826 14716
rect 14762 14656 14826 14660
rect 19950 14716 20014 14720
rect 19950 14660 19954 14716
rect 19954 14660 20010 14716
rect 20010 14660 20014 14716
rect 19950 14656 20014 14660
rect 20030 14716 20094 14720
rect 20030 14660 20034 14716
rect 20034 14660 20090 14716
rect 20090 14660 20094 14716
rect 20030 14656 20094 14660
rect 20110 14716 20174 14720
rect 20110 14660 20114 14716
rect 20114 14660 20170 14716
rect 20170 14660 20174 14716
rect 20110 14656 20174 14660
rect 20190 14716 20254 14720
rect 20190 14660 20194 14716
rect 20194 14660 20250 14716
rect 20250 14660 20254 14716
rect 20190 14656 20254 14660
rect 6380 14172 6444 14176
rect 6380 14116 6384 14172
rect 6384 14116 6440 14172
rect 6440 14116 6444 14172
rect 6380 14112 6444 14116
rect 6460 14172 6524 14176
rect 6460 14116 6464 14172
rect 6464 14116 6520 14172
rect 6520 14116 6524 14172
rect 6460 14112 6524 14116
rect 6540 14172 6604 14176
rect 6540 14116 6544 14172
rect 6544 14116 6600 14172
rect 6600 14116 6604 14172
rect 6540 14112 6604 14116
rect 6620 14172 6684 14176
rect 6620 14116 6624 14172
rect 6624 14116 6680 14172
rect 6680 14116 6684 14172
rect 6620 14112 6684 14116
rect 11808 14172 11872 14176
rect 11808 14116 11812 14172
rect 11812 14116 11868 14172
rect 11868 14116 11872 14172
rect 11808 14112 11872 14116
rect 11888 14172 11952 14176
rect 11888 14116 11892 14172
rect 11892 14116 11948 14172
rect 11948 14116 11952 14172
rect 11888 14112 11952 14116
rect 11968 14172 12032 14176
rect 11968 14116 11972 14172
rect 11972 14116 12028 14172
rect 12028 14116 12032 14172
rect 11968 14112 12032 14116
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 17316 14172 17380 14176
rect 17316 14116 17320 14172
rect 17320 14116 17376 14172
rect 17376 14116 17380 14172
rect 17316 14112 17380 14116
rect 17396 14172 17460 14176
rect 17396 14116 17400 14172
rect 17400 14116 17456 14172
rect 17456 14116 17460 14172
rect 17396 14112 17460 14116
rect 17476 14172 17540 14176
rect 17476 14116 17480 14172
rect 17480 14116 17536 14172
rect 17536 14116 17540 14172
rect 17476 14112 17540 14116
rect 22664 14172 22728 14176
rect 22664 14116 22668 14172
rect 22668 14116 22724 14172
rect 22724 14116 22728 14172
rect 22664 14112 22728 14116
rect 22744 14172 22808 14176
rect 22744 14116 22748 14172
rect 22748 14116 22804 14172
rect 22804 14116 22808 14172
rect 22744 14112 22808 14116
rect 22824 14172 22888 14176
rect 22824 14116 22828 14172
rect 22828 14116 22884 14172
rect 22884 14116 22888 14172
rect 22824 14112 22888 14116
rect 22904 14172 22968 14176
rect 22904 14116 22908 14172
rect 22908 14116 22964 14172
rect 22964 14116 22968 14172
rect 22904 14112 22968 14116
rect 3666 13628 3730 13632
rect 3666 13572 3670 13628
rect 3670 13572 3726 13628
rect 3726 13572 3730 13628
rect 3666 13568 3730 13572
rect 3746 13628 3810 13632
rect 3746 13572 3750 13628
rect 3750 13572 3806 13628
rect 3806 13572 3810 13628
rect 3746 13568 3810 13572
rect 3826 13628 3890 13632
rect 3826 13572 3830 13628
rect 3830 13572 3886 13628
rect 3886 13572 3890 13628
rect 3826 13568 3890 13572
rect 3906 13628 3970 13632
rect 3906 13572 3910 13628
rect 3910 13572 3966 13628
rect 3966 13572 3970 13628
rect 3906 13568 3970 13572
rect 9094 13628 9158 13632
rect 9094 13572 9098 13628
rect 9098 13572 9154 13628
rect 9154 13572 9158 13628
rect 9094 13568 9158 13572
rect 9174 13628 9238 13632
rect 9174 13572 9178 13628
rect 9178 13572 9234 13628
rect 9234 13572 9238 13628
rect 9174 13568 9238 13572
rect 9254 13628 9318 13632
rect 9254 13572 9258 13628
rect 9258 13572 9314 13628
rect 9314 13572 9318 13628
rect 9254 13568 9318 13572
rect 9334 13628 9398 13632
rect 9334 13572 9338 13628
rect 9338 13572 9394 13628
rect 9394 13572 9398 13628
rect 9334 13568 9398 13572
rect 14522 13628 14586 13632
rect 14522 13572 14526 13628
rect 14526 13572 14582 13628
rect 14582 13572 14586 13628
rect 14522 13568 14586 13572
rect 14602 13628 14666 13632
rect 14602 13572 14606 13628
rect 14606 13572 14662 13628
rect 14662 13572 14666 13628
rect 14602 13568 14666 13572
rect 14682 13628 14746 13632
rect 14682 13572 14686 13628
rect 14686 13572 14742 13628
rect 14742 13572 14746 13628
rect 14682 13568 14746 13572
rect 14762 13628 14826 13632
rect 14762 13572 14766 13628
rect 14766 13572 14822 13628
rect 14822 13572 14826 13628
rect 14762 13568 14826 13572
rect 19950 13628 20014 13632
rect 19950 13572 19954 13628
rect 19954 13572 20010 13628
rect 20010 13572 20014 13628
rect 19950 13568 20014 13572
rect 20030 13628 20094 13632
rect 20030 13572 20034 13628
rect 20034 13572 20090 13628
rect 20090 13572 20094 13628
rect 20030 13568 20094 13572
rect 20110 13628 20174 13632
rect 20110 13572 20114 13628
rect 20114 13572 20170 13628
rect 20170 13572 20174 13628
rect 20110 13568 20174 13572
rect 20190 13628 20254 13632
rect 20190 13572 20194 13628
rect 20194 13572 20250 13628
rect 20250 13572 20254 13628
rect 20190 13568 20254 13572
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 11808 13084 11872 13088
rect 11808 13028 11812 13084
rect 11812 13028 11868 13084
rect 11868 13028 11872 13084
rect 11808 13024 11872 13028
rect 11888 13084 11952 13088
rect 11888 13028 11892 13084
rect 11892 13028 11948 13084
rect 11948 13028 11952 13084
rect 11888 13024 11952 13028
rect 11968 13084 12032 13088
rect 11968 13028 11972 13084
rect 11972 13028 12028 13084
rect 12028 13028 12032 13084
rect 11968 13024 12032 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 17316 13084 17380 13088
rect 17316 13028 17320 13084
rect 17320 13028 17376 13084
rect 17376 13028 17380 13084
rect 17316 13024 17380 13028
rect 17396 13084 17460 13088
rect 17396 13028 17400 13084
rect 17400 13028 17456 13084
rect 17456 13028 17460 13084
rect 17396 13024 17460 13028
rect 17476 13084 17540 13088
rect 17476 13028 17480 13084
rect 17480 13028 17536 13084
rect 17536 13028 17540 13084
rect 17476 13024 17540 13028
rect 22664 13084 22728 13088
rect 22664 13028 22668 13084
rect 22668 13028 22724 13084
rect 22724 13028 22728 13084
rect 22664 13024 22728 13028
rect 22744 13084 22808 13088
rect 22744 13028 22748 13084
rect 22748 13028 22804 13084
rect 22804 13028 22808 13084
rect 22744 13024 22808 13028
rect 22824 13084 22888 13088
rect 22824 13028 22828 13084
rect 22828 13028 22884 13084
rect 22884 13028 22888 13084
rect 22824 13024 22888 13028
rect 22904 13084 22968 13088
rect 22904 13028 22908 13084
rect 22908 13028 22964 13084
rect 22964 13028 22968 13084
rect 22904 13024 22968 13028
rect 3666 12540 3730 12544
rect 3666 12484 3670 12540
rect 3670 12484 3726 12540
rect 3726 12484 3730 12540
rect 3666 12480 3730 12484
rect 3746 12540 3810 12544
rect 3746 12484 3750 12540
rect 3750 12484 3806 12540
rect 3806 12484 3810 12540
rect 3746 12480 3810 12484
rect 3826 12540 3890 12544
rect 3826 12484 3830 12540
rect 3830 12484 3886 12540
rect 3886 12484 3890 12540
rect 3826 12480 3890 12484
rect 3906 12540 3970 12544
rect 3906 12484 3910 12540
rect 3910 12484 3966 12540
rect 3966 12484 3970 12540
rect 3906 12480 3970 12484
rect 9094 12540 9158 12544
rect 9094 12484 9098 12540
rect 9098 12484 9154 12540
rect 9154 12484 9158 12540
rect 9094 12480 9158 12484
rect 9174 12540 9238 12544
rect 9174 12484 9178 12540
rect 9178 12484 9234 12540
rect 9234 12484 9238 12540
rect 9174 12480 9238 12484
rect 9254 12540 9318 12544
rect 9254 12484 9258 12540
rect 9258 12484 9314 12540
rect 9314 12484 9318 12540
rect 9254 12480 9318 12484
rect 9334 12540 9398 12544
rect 9334 12484 9338 12540
rect 9338 12484 9394 12540
rect 9394 12484 9398 12540
rect 9334 12480 9398 12484
rect 14522 12540 14586 12544
rect 14522 12484 14526 12540
rect 14526 12484 14582 12540
rect 14582 12484 14586 12540
rect 14522 12480 14586 12484
rect 14602 12540 14666 12544
rect 14602 12484 14606 12540
rect 14606 12484 14662 12540
rect 14662 12484 14666 12540
rect 14602 12480 14666 12484
rect 14682 12540 14746 12544
rect 14682 12484 14686 12540
rect 14686 12484 14742 12540
rect 14742 12484 14746 12540
rect 14682 12480 14746 12484
rect 14762 12540 14826 12544
rect 14762 12484 14766 12540
rect 14766 12484 14822 12540
rect 14822 12484 14826 12540
rect 14762 12480 14826 12484
rect 19950 12540 20014 12544
rect 19950 12484 19954 12540
rect 19954 12484 20010 12540
rect 20010 12484 20014 12540
rect 19950 12480 20014 12484
rect 20030 12540 20094 12544
rect 20030 12484 20034 12540
rect 20034 12484 20090 12540
rect 20090 12484 20094 12540
rect 20030 12480 20094 12484
rect 20110 12540 20174 12544
rect 20110 12484 20114 12540
rect 20114 12484 20170 12540
rect 20170 12484 20174 12540
rect 20110 12480 20174 12484
rect 20190 12540 20254 12544
rect 20190 12484 20194 12540
rect 20194 12484 20250 12540
rect 20250 12484 20254 12540
rect 20190 12480 20254 12484
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 11808 11996 11872 12000
rect 11808 11940 11812 11996
rect 11812 11940 11868 11996
rect 11868 11940 11872 11996
rect 11808 11936 11872 11940
rect 11888 11996 11952 12000
rect 11888 11940 11892 11996
rect 11892 11940 11948 11996
rect 11948 11940 11952 11996
rect 11888 11936 11952 11940
rect 11968 11996 12032 12000
rect 11968 11940 11972 11996
rect 11972 11940 12028 11996
rect 12028 11940 12032 11996
rect 11968 11936 12032 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 17316 11996 17380 12000
rect 17316 11940 17320 11996
rect 17320 11940 17376 11996
rect 17376 11940 17380 11996
rect 17316 11936 17380 11940
rect 17396 11996 17460 12000
rect 17396 11940 17400 11996
rect 17400 11940 17456 11996
rect 17456 11940 17460 11996
rect 17396 11936 17460 11940
rect 17476 11996 17540 12000
rect 17476 11940 17480 11996
rect 17480 11940 17536 11996
rect 17536 11940 17540 11996
rect 17476 11936 17540 11940
rect 22664 11996 22728 12000
rect 22664 11940 22668 11996
rect 22668 11940 22724 11996
rect 22724 11940 22728 11996
rect 22664 11936 22728 11940
rect 22744 11996 22808 12000
rect 22744 11940 22748 11996
rect 22748 11940 22804 11996
rect 22804 11940 22808 11996
rect 22744 11936 22808 11940
rect 22824 11996 22888 12000
rect 22824 11940 22828 11996
rect 22828 11940 22884 11996
rect 22884 11940 22888 11996
rect 22824 11936 22888 11940
rect 22904 11996 22968 12000
rect 22904 11940 22908 11996
rect 22908 11940 22964 11996
rect 22964 11940 22968 11996
rect 22904 11936 22968 11940
rect 3666 11452 3730 11456
rect 3666 11396 3670 11452
rect 3670 11396 3726 11452
rect 3726 11396 3730 11452
rect 3666 11392 3730 11396
rect 3746 11452 3810 11456
rect 3746 11396 3750 11452
rect 3750 11396 3806 11452
rect 3806 11396 3810 11452
rect 3746 11392 3810 11396
rect 3826 11452 3890 11456
rect 3826 11396 3830 11452
rect 3830 11396 3886 11452
rect 3886 11396 3890 11452
rect 3826 11392 3890 11396
rect 3906 11452 3970 11456
rect 3906 11396 3910 11452
rect 3910 11396 3966 11452
rect 3966 11396 3970 11452
rect 3906 11392 3970 11396
rect 9094 11452 9158 11456
rect 9094 11396 9098 11452
rect 9098 11396 9154 11452
rect 9154 11396 9158 11452
rect 9094 11392 9158 11396
rect 9174 11452 9238 11456
rect 9174 11396 9178 11452
rect 9178 11396 9234 11452
rect 9234 11396 9238 11452
rect 9174 11392 9238 11396
rect 9254 11452 9318 11456
rect 9254 11396 9258 11452
rect 9258 11396 9314 11452
rect 9314 11396 9318 11452
rect 9254 11392 9318 11396
rect 9334 11452 9398 11456
rect 9334 11396 9338 11452
rect 9338 11396 9394 11452
rect 9394 11396 9398 11452
rect 9334 11392 9398 11396
rect 14522 11452 14586 11456
rect 14522 11396 14526 11452
rect 14526 11396 14582 11452
rect 14582 11396 14586 11452
rect 14522 11392 14586 11396
rect 14602 11452 14666 11456
rect 14602 11396 14606 11452
rect 14606 11396 14662 11452
rect 14662 11396 14666 11452
rect 14602 11392 14666 11396
rect 14682 11452 14746 11456
rect 14682 11396 14686 11452
rect 14686 11396 14742 11452
rect 14742 11396 14746 11452
rect 14682 11392 14746 11396
rect 14762 11452 14826 11456
rect 14762 11396 14766 11452
rect 14766 11396 14822 11452
rect 14822 11396 14826 11452
rect 14762 11392 14826 11396
rect 19950 11452 20014 11456
rect 19950 11396 19954 11452
rect 19954 11396 20010 11452
rect 20010 11396 20014 11452
rect 19950 11392 20014 11396
rect 20030 11452 20094 11456
rect 20030 11396 20034 11452
rect 20034 11396 20090 11452
rect 20090 11396 20094 11452
rect 20030 11392 20094 11396
rect 20110 11452 20174 11456
rect 20110 11396 20114 11452
rect 20114 11396 20170 11452
rect 20170 11396 20174 11452
rect 20110 11392 20174 11396
rect 20190 11452 20254 11456
rect 20190 11396 20194 11452
rect 20194 11396 20250 11452
rect 20250 11396 20254 11452
rect 20190 11392 20254 11396
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 11808 10908 11872 10912
rect 11808 10852 11812 10908
rect 11812 10852 11868 10908
rect 11868 10852 11872 10908
rect 11808 10848 11872 10852
rect 11888 10908 11952 10912
rect 11888 10852 11892 10908
rect 11892 10852 11948 10908
rect 11948 10852 11952 10908
rect 11888 10848 11952 10852
rect 11968 10908 12032 10912
rect 11968 10852 11972 10908
rect 11972 10852 12028 10908
rect 12028 10852 12032 10908
rect 11968 10848 12032 10852
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 17316 10908 17380 10912
rect 17316 10852 17320 10908
rect 17320 10852 17376 10908
rect 17376 10852 17380 10908
rect 17316 10848 17380 10852
rect 17396 10908 17460 10912
rect 17396 10852 17400 10908
rect 17400 10852 17456 10908
rect 17456 10852 17460 10908
rect 17396 10848 17460 10852
rect 17476 10908 17540 10912
rect 17476 10852 17480 10908
rect 17480 10852 17536 10908
rect 17536 10852 17540 10908
rect 17476 10848 17540 10852
rect 22664 10908 22728 10912
rect 22664 10852 22668 10908
rect 22668 10852 22724 10908
rect 22724 10852 22728 10908
rect 22664 10848 22728 10852
rect 22744 10908 22808 10912
rect 22744 10852 22748 10908
rect 22748 10852 22804 10908
rect 22804 10852 22808 10908
rect 22744 10848 22808 10852
rect 22824 10908 22888 10912
rect 22824 10852 22828 10908
rect 22828 10852 22884 10908
rect 22884 10852 22888 10908
rect 22824 10848 22888 10852
rect 22904 10908 22968 10912
rect 22904 10852 22908 10908
rect 22908 10852 22964 10908
rect 22964 10852 22968 10908
rect 22904 10848 22968 10852
rect 15148 10568 15212 10572
rect 15148 10512 15198 10568
rect 15198 10512 15212 10568
rect 15148 10508 15212 10512
rect 3666 10364 3730 10368
rect 3666 10308 3670 10364
rect 3670 10308 3726 10364
rect 3726 10308 3730 10364
rect 3666 10304 3730 10308
rect 3746 10364 3810 10368
rect 3746 10308 3750 10364
rect 3750 10308 3806 10364
rect 3806 10308 3810 10364
rect 3746 10304 3810 10308
rect 3826 10364 3890 10368
rect 3826 10308 3830 10364
rect 3830 10308 3886 10364
rect 3886 10308 3890 10364
rect 3826 10304 3890 10308
rect 3906 10364 3970 10368
rect 3906 10308 3910 10364
rect 3910 10308 3966 10364
rect 3966 10308 3970 10364
rect 3906 10304 3970 10308
rect 9094 10364 9158 10368
rect 9094 10308 9098 10364
rect 9098 10308 9154 10364
rect 9154 10308 9158 10364
rect 9094 10304 9158 10308
rect 9174 10364 9238 10368
rect 9174 10308 9178 10364
rect 9178 10308 9234 10364
rect 9234 10308 9238 10364
rect 9174 10304 9238 10308
rect 9254 10364 9318 10368
rect 9254 10308 9258 10364
rect 9258 10308 9314 10364
rect 9314 10308 9318 10364
rect 9254 10304 9318 10308
rect 9334 10364 9398 10368
rect 9334 10308 9338 10364
rect 9338 10308 9394 10364
rect 9394 10308 9398 10364
rect 9334 10304 9398 10308
rect 14522 10364 14586 10368
rect 14522 10308 14526 10364
rect 14526 10308 14582 10364
rect 14582 10308 14586 10364
rect 14522 10304 14586 10308
rect 14602 10364 14666 10368
rect 14602 10308 14606 10364
rect 14606 10308 14662 10364
rect 14662 10308 14666 10364
rect 14602 10304 14666 10308
rect 14682 10364 14746 10368
rect 14682 10308 14686 10364
rect 14686 10308 14742 10364
rect 14742 10308 14746 10364
rect 14682 10304 14746 10308
rect 14762 10364 14826 10368
rect 14762 10308 14766 10364
rect 14766 10308 14822 10364
rect 14822 10308 14826 10364
rect 14762 10304 14826 10308
rect 19950 10364 20014 10368
rect 19950 10308 19954 10364
rect 19954 10308 20010 10364
rect 20010 10308 20014 10364
rect 19950 10304 20014 10308
rect 20030 10364 20094 10368
rect 20030 10308 20034 10364
rect 20034 10308 20090 10364
rect 20090 10308 20094 10364
rect 20030 10304 20094 10308
rect 20110 10364 20174 10368
rect 20110 10308 20114 10364
rect 20114 10308 20170 10364
rect 20170 10308 20174 10364
rect 20110 10304 20174 10308
rect 20190 10364 20254 10368
rect 20190 10308 20194 10364
rect 20194 10308 20250 10364
rect 20250 10308 20254 10364
rect 20190 10304 20254 10308
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 11808 9820 11872 9824
rect 11808 9764 11812 9820
rect 11812 9764 11868 9820
rect 11868 9764 11872 9820
rect 11808 9760 11872 9764
rect 11888 9820 11952 9824
rect 11888 9764 11892 9820
rect 11892 9764 11948 9820
rect 11948 9764 11952 9820
rect 11888 9760 11952 9764
rect 11968 9820 12032 9824
rect 11968 9764 11972 9820
rect 11972 9764 12028 9820
rect 12028 9764 12032 9820
rect 11968 9760 12032 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 17316 9820 17380 9824
rect 17316 9764 17320 9820
rect 17320 9764 17376 9820
rect 17376 9764 17380 9820
rect 17316 9760 17380 9764
rect 17396 9820 17460 9824
rect 17396 9764 17400 9820
rect 17400 9764 17456 9820
rect 17456 9764 17460 9820
rect 17396 9760 17460 9764
rect 17476 9820 17540 9824
rect 17476 9764 17480 9820
rect 17480 9764 17536 9820
rect 17536 9764 17540 9820
rect 17476 9760 17540 9764
rect 22664 9820 22728 9824
rect 22664 9764 22668 9820
rect 22668 9764 22724 9820
rect 22724 9764 22728 9820
rect 22664 9760 22728 9764
rect 22744 9820 22808 9824
rect 22744 9764 22748 9820
rect 22748 9764 22804 9820
rect 22804 9764 22808 9820
rect 22744 9760 22808 9764
rect 22824 9820 22888 9824
rect 22824 9764 22828 9820
rect 22828 9764 22884 9820
rect 22884 9764 22888 9820
rect 22824 9760 22888 9764
rect 22904 9820 22968 9824
rect 22904 9764 22908 9820
rect 22908 9764 22964 9820
rect 22964 9764 22968 9820
rect 22904 9760 22968 9764
rect 3666 9276 3730 9280
rect 3666 9220 3670 9276
rect 3670 9220 3726 9276
rect 3726 9220 3730 9276
rect 3666 9216 3730 9220
rect 3746 9276 3810 9280
rect 3746 9220 3750 9276
rect 3750 9220 3806 9276
rect 3806 9220 3810 9276
rect 3746 9216 3810 9220
rect 3826 9276 3890 9280
rect 3826 9220 3830 9276
rect 3830 9220 3886 9276
rect 3886 9220 3890 9276
rect 3826 9216 3890 9220
rect 3906 9276 3970 9280
rect 3906 9220 3910 9276
rect 3910 9220 3966 9276
rect 3966 9220 3970 9276
rect 3906 9216 3970 9220
rect 9094 9276 9158 9280
rect 9094 9220 9098 9276
rect 9098 9220 9154 9276
rect 9154 9220 9158 9276
rect 9094 9216 9158 9220
rect 9174 9276 9238 9280
rect 9174 9220 9178 9276
rect 9178 9220 9234 9276
rect 9234 9220 9238 9276
rect 9174 9216 9238 9220
rect 9254 9276 9318 9280
rect 9254 9220 9258 9276
rect 9258 9220 9314 9276
rect 9314 9220 9318 9276
rect 9254 9216 9318 9220
rect 9334 9276 9398 9280
rect 9334 9220 9338 9276
rect 9338 9220 9394 9276
rect 9394 9220 9398 9276
rect 9334 9216 9398 9220
rect 14522 9276 14586 9280
rect 14522 9220 14526 9276
rect 14526 9220 14582 9276
rect 14582 9220 14586 9276
rect 14522 9216 14586 9220
rect 14602 9276 14666 9280
rect 14602 9220 14606 9276
rect 14606 9220 14662 9276
rect 14662 9220 14666 9276
rect 14602 9216 14666 9220
rect 14682 9276 14746 9280
rect 14682 9220 14686 9276
rect 14686 9220 14742 9276
rect 14742 9220 14746 9276
rect 14682 9216 14746 9220
rect 14762 9276 14826 9280
rect 14762 9220 14766 9276
rect 14766 9220 14822 9276
rect 14822 9220 14826 9276
rect 14762 9216 14826 9220
rect 19950 9276 20014 9280
rect 19950 9220 19954 9276
rect 19954 9220 20010 9276
rect 20010 9220 20014 9276
rect 19950 9216 20014 9220
rect 20030 9276 20094 9280
rect 20030 9220 20034 9276
rect 20034 9220 20090 9276
rect 20090 9220 20094 9276
rect 20030 9216 20094 9220
rect 20110 9276 20174 9280
rect 20110 9220 20114 9276
rect 20114 9220 20170 9276
rect 20170 9220 20174 9276
rect 20110 9216 20174 9220
rect 20190 9276 20254 9280
rect 20190 9220 20194 9276
rect 20194 9220 20250 9276
rect 20250 9220 20254 9276
rect 20190 9216 20254 9220
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 11808 8732 11872 8736
rect 11808 8676 11812 8732
rect 11812 8676 11868 8732
rect 11868 8676 11872 8732
rect 11808 8672 11872 8676
rect 11888 8732 11952 8736
rect 11888 8676 11892 8732
rect 11892 8676 11948 8732
rect 11948 8676 11952 8732
rect 11888 8672 11952 8676
rect 11968 8732 12032 8736
rect 11968 8676 11972 8732
rect 11972 8676 12028 8732
rect 12028 8676 12032 8732
rect 11968 8672 12032 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 17316 8732 17380 8736
rect 17316 8676 17320 8732
rect 17320 8676 17376 8732
rect 17376 8676 17380 8732
rect 17316 8672 17380 8676
rect 17396 8732 17460 8736
rect 17396 8676 17400 8732
rect 17400 8676 17456 8732
rect 17456 8676 17460 8732
rect 17396 8672 17460 8676
rect 17476 8732 17540 8736
rect 17476 8676 17480 8732
rect 17480 8676 17536 8732
rect 17536 8676 17540 8732
rect 17476 8672 17540 8676
rect 22664 8732 22728 8736
rect 22664 8676 22668 8732
rect 22668 8676 22724 8732
rect 22724 8676 22728 8732
rect 22664 8672 22728 8676
rect 22744 8732 22808 8736
rect 22744 8676 22748 8732
rect 22748 8676 22804 8732
rect 22804 8676 22808 8732
rect 22744 8672 22808 8676
rect 22824 8732 22888 8736
rect 22824 8676 22828 8732
rect 22828 8676 22884 8732
rect 22884 8676 22888 8732
rect 22824 8672 22888 8676
rect 22904 8732 22968 8736
rect 22904 8676 22908 8732
rect 22908 8676 22964 8732
rect 22964 8676 22968 8732
rect 22904 8672 22968 8676
rect 3666 8188 3730 8192
rect 3666 8132 3670 8188
rect 3670 8132 3726 8188
rect 3726 8132 3730 8188
rect 3666 8128 3730 8132
rect 3746 8188 3810 8192
rect 3746 8132 3750 8188
rect 3750 8132 3806 8188
rect 3806 8132 3810 8188
rect 3746 8128 3810 8132
rect 3826 8188 3890 8192
rect 3826 8132 3830 8188
rect 3830 8132 3886 8188
rect 3886 8132 3890 8188
rect 3826 8128 3890 8132
rect 3906 8188 3970 8192
rect 3906 8132 3910 8188
rect 3910 8132 3966 8188
rect 3966 8132 3970 8188
rect 3906 8128 3970 8132
rect 9094 8188 9158 8192
rect 9094 8132 9098 8188
rect 9098 8132 9154 8188
rect 9154 8132 9158 8188
rect 9094 8128 9158 8132
rect 9174 8188 9238 8192
rect 9174 8132 9178 8188
rect 9178 8132 9234 8188
rect 9234 8132 9238 8188
rect 9174 8128 9238 8132
rect 9254 8188 9318 8192
rect 9254 8132 9258 8188
rect 9258 8132 9314 8188
rect 9314 8132 9318 8188
rect 9254 8128 9318 8132
rect 9334 8188 9398 8192
rect 9334 8132 9338 8188
rect 9338 8132 9394 8188
rect 9394 8132 9398 8188
rect 9334 8128 9398 8132
rect 14522 8188 14586 8192
rect 14522 8132 14526 8188
rect 14526 8132 14582 8188
rect 14582 8132 14586 8188
rect 14522 8128 14586 8132
rect 14602 8188 14666 8192
rect 14602 8132 14606 8188
rect 14606 8132 14662 8188
rect 14662 8132 14666 8188
rect 14602 8128 14666 8132
rect 14682 8188 14746 8192
rect 14682 8132 14686 8188
rect 14686 8132 14742 8188
rect 14742 8132 14746 8188
rect 14682 8128 14746 8132
rect 14762 8188 14826 8192
rect 14762 8132 14766 8188
rect 14766 8132 14822 8188
rect 14822 8132 14826 8188
rect 14762 8128 14826 8132
rect 19950 8188 20014 8192
rect 19950 8132 19954 8188
rect 19954 8132 20010 8188
rect 20010 8132 20014 8188
rect 19950 8128 20014 8132
rect 20030 8188 20094 8192
rect 20030 8132 20034 8188
rect 20034 8132 20090 8188
rect 20090 8132 20094 8188
rect 20030 8128 20094 8132
rect 20110 8188 20174 8192
rect 20110 8132 20114 8188
rect 20114 8132 20170 8188
rect 20170 8132 20174 8188
rect 20110 8128 20174 8132
rect 20190 8188 20254 8192
rect 20190 8132 20194 8188
rect 20194 8132 20250 8188
rect 20250 8132 20254 8188
rect 20190 8128 20254 8132
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 11808 7644 11872 7648
rect 11808 7588 11812 7644
rect 11812 7588 11868 7644
rect 11868 7588 11872 7644
rect 11808 7584 11872 7588
rect 11888 7644 11952 7648
rect 11888 7588 11892 7644
rect 11892 7588 11948 7644
rect 11948 7588 11952 7644
rect 11888 7584 11952 7588
rect 11968 7644 12032 7648
rect 11968 7588 11972 7644
rect 11972 7588 12028 7644
rect 12028 7588 12032 7644
rect 11968 7584 12032 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 17316 7644 17380 7648
rect 17316 7588 17320 7644
rect 17320 7588 17376 7644
rect 17376 7588 17380 7644
rect 17316 7584 17380 7588
rect 17396 7644 17460 7648
rect 17396 7588 17400 7644
rect 17400 7588 17456 7644
rect 17456 7588 17460 7644
rect 17396 7584 17460 7588
rect 17476 7644 17540 7648
rect 17476 7588 17480 7644
rect 17480 7588 17536 7644
rect 17536 7588 17540 7644
rect 17476 7584 17540 7588
rect 22664 7644 22728 7648
rect 22664 7588 22668 7644
rect 22668 7588 22724 7644
rect 22724 7588 22728 7644
rect 22664 7584 22728 7588
rect 22744 7644 22808 7648
rect 22744 7588 22748 7644
rect 22748 7588 22804 7644
rect 22804 7588 22808 7644
rect 22744 7584 22808 7588
rect 22824 7644 22888 7648
rect 22824 7588 22828 7644
rect 22828 7588 22884 7644
rect 22884 7588 22888 7644
rect 22824 7584 22888 7588
rect 22904 7644 22968 7648
rect 22904 7588 22908 7644
rect 22908 7588 22964 7644
rect 22964 7588 22968 7644
rect 22904 7584 22968 7588
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 9094 7100 9158 7104
rect 9094 7044 9098 7100
rect 9098 7044 9154 7100
rect 9154 7044 9158 7100
rect 9094 7040 9158 7044
rect 9174 7100 9238 7104
rect 9174 7044 9178 7100
rect 9178 7044 9234 7100
rect 9234 7044 9238 7100
rect 9174 7040 9238 7044
rect 9254 7100 9318 7104
rect 9254 7044 9258 7100
rect 9258 7044 9314 7100
rect 9314 7044 9318 7100
rect 9254 7040 9318 7044
rect 9334 7100 9398 7104
rect 9334 7044 9338 7100
rect 9338 7044 9394 7100
rect 9394 7044 9398 7100
rect 9334 7040 9398 7044
rect 14522 7100 14586 7104
rect 14522 7044 14526 7100
rect 14526 7044 14582 7100
rect 14582 7044 14586 7100
rect 14522 7040 14586 7044
rect 14602 7100 14666 7104
rect 14602 7044 14606 7100
rect 14606 7044 14662 7100
rect 14662 7044 14666 7100
rect 14602 7040 14666 7044
rect 14682 7100 14746 7104
rect 14682 7044 14686 7100
rect 14686 7044 14742 7100
rect 14742 7044 14746 7100
rect 14682 7040 14746 7044
rect 14762 7100 14826 7104
rect 14762 7044 14766 7100
rect 14766 7044 14822 7100
rect 14822 7044 14826 7100
rect 14762 7040 14826 7044
rect 19950 7100 20014 7104
rect 19950 7044 19954 7100
rect 19954 7044 20010 7100
rect 20010 7044 20014 7100
rect 19950 7040 20014 7044
rect 20030 7100 20094 7104
rect 20030 7044 20034 7100
rect 20034 7044 20090 7100
rect 20090 7044 20094 7100
rect 20030 7040 20094 7044
rect 20110 7100 20174 7104
rect 20110 7044 20114 7100
rect 20114 7044 20170 7100
rect 20170 7044 20174 7100
rect 20110 7040 20174 7044
rect 20190 7100 20254 7104
rect 20190 7044 20194 7100
rect 20194 7044 20250 7100
rect 20250 7044 20254 7100
rect 20190 7040 20254 7044
rect 15148 6700 15212 6764
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 11808 6556 11872 6560
rect 11808 6500 11812 6556
rect 11812 6500 11868 6556
rect 11868 6500 11872 6556
rect 11808 6496 11872 6500
rect 11888 6556 11952 6560
rect 11888 6500 11892 6556
rect 11892 6500 11948 6556
rect 11948 6500 11952 6556
rect 11888 6496 11952 6500
rect 11968 6556 12032 6560
rect 11968 6500 11972 6556
rect 11972 6500 12028 6556
rect 12028 6500 12032 6556
rect 11968 6496 12032 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 17316 6556 17380 6560
rect 17316 6500 17320 6556
rect 17320 6500 17376 6556
rect 17376 6500 17380 6556
rect 17316 6496 17380 6500
rect 17396 6556 17460 6560
rect 17396 6500 17400 6556
rect 17400 6500 17456 6556
rect 17456 6500 17460 6556
rect 17396 6496 17460 6500
rect 17476 6556 17540 6560
rect 17476 6500 17480 6556
rect 17480 6500 17536 6556
rect 17536 6500 17540 6556
rect 17476 6496 17540 6500
rect 22664 6556 22728 6560
rect 22664 6500 22668 6556
rect 22668 6500 22724 6556
rect 22724 6500 22728 6556
rect 22664 6496 22728 6500
rect 22744 6556 22808 6560
rect 22744 6500 22748 6556
rect 22748 6500 22804 6556
rect 22804 6500 22808 6556
rect 22744 6496 22808 6500
rect 22824 6556 22888 6560
rect 22824 6500 22828 6556
rect 22828 6500 22884 6556
rect 22884 6500 22888 6556
rect 22824 6496 22888 6500
rect 22904 6556 22968 6560
rect 22904 6500 22908 6556
rect 22908 6500 22964 6556
rect 22964 6500 22968 6556
rect 22904 6496 22968 6500
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 9094 6012 9158 6016
rect 9094 5956 9098 6012
rect 9098 5956 9154 6012
rect 9154 5956 9158 6012
rect 9094 5952 9158 5956
rect 9174 6012 9238 6016
rect 9174 5956 9178 6012
rect 9178 5956 9234 6012
rect 9234 5956 9238 6012
rect 9174 5952 9238 5956
rect 9254 6012 9318 6016
rect 9254 5956 9258 6012
rect 9258 5956 9314 6012
rect 9314 5956 9318 6012
rect 9254 5952 9318 5956
rect 9334 6012 9398 6016
rect 9334 5956 9338 6012
rect 9338 5956 9394 6012
rect 9394 5956 9398 6012
rect 9334 5952 9398 5956
rect 14522 6012 14586 6016
rect 14522 5956 14526 6012
rect 14526 5956 14582 6012
rect 14582 5956 14586 6012
rect 14522 5952 14586 5956
rect 14602 6012 14666 6016
rect 14602 5956 14606 6012
rect 14606 5956 14662 6012
rect 14662 5956 14666 6012
rect 14602 5952 14666 5956
rect 14682 6012 14746 6016
rect 14682 5956 14686 6012
rect 14686 5956 14742 6012
rect 14742 5956 14746 6012
rect 14682 5952 14746 5956
rect 14762 6012 14826 6016
rect 14762 5956 14766 6012
rect 14766 5956 14822 6012
rect 14822 5956 14826 6012
rect 14762 5952 14826 5956
rect 19950 6012 20014 6016
rect 19950 5956 19954 6012
rect 19954 5956 20010 6012
rect 20010 5956 20014 6012
rect 19950 5952 20014 5956
rect 20030 6012 20094 6016
rect 20030 5956 20034 6012
rect 20034 5956 20090 6012
rect 20090 5956 20094 6012
rect 20030 5952 20094 5956
rect 20110 6012 20174 6016
rect 20110 5956 20114 6012
rect 20114 5956 20170 6012
rect 20170 5956 20174 6012
rect 20110 5952 20174 5956
rect 20190 6012 20254 6016
rect 20190 5956 20194 6012
rect 20194 5956 20250 6012
rect 20250 5956 20254 6012
rect 20190 5952 20254 5956
rect 19564 5672 19628 5676
rect 19564 5616 19614 5672
rect 19614 5616 19628 5672
rect 19564 5612 19628 5616
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 11808 5468 11872 5472
rect 11808 5412 11812 5468
rect 11812 5412 11868 5468
rect 11868 5412 11872 5468
rect 11808 5408 11872 5412
rect 11888 5468 11952 5472
rect 11888 5412 11892 5468
rect 11892 5412 11948 5468
rect 11948 5412 11952 5468
rect 11888 5408 11952 5412
rect 11968 5468 12032 5472
rect 11968 5412 11972 5468
rect 11972 5412 12028 5468
rect 12028 5412 12032 5468
rect 11968 5408 12032 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 17316 5468 17380 5472
rect 17316 5412 17320 5468
rect 17320 5412 17376 5468
rect 17376 5412 17380 5468
rect 17316 5408 17380 5412
rect 17396 5468 17460 5472
rect 17396 5412 17400 5468
rect 17400 5412 17456 5468
rect 17456 5412 17460 5468
rect 17396 5408 17460 5412
rect 17476 5468 17540 5472
rect 17476 5412 17480 5468
rect 17480 5412 17536 5468
rect 17536 5412 17540 5468
rect 17476 5408 17540 5412
rect 22664 5468 22728 5472
rect 22664 5412 22668 5468
rect 22668 5412 22724 5468
rect 22724 5412 22728 5468
rect 22664 5408 22728 5412
rect 22744 5468 22808 5472
rect 22744 5412 22748 5468
rect 22748 5412 22804 5468
rect 22804 5412 22808 5468
rect 22744 5408 22808 5412
rect 22824 5468 22888 5472
rect 22824 5412 22828 5468
rect 22828 5412 22884 5468
rect 22884 5412 22888 5468
rect 22824 5408 22888 5412
rect 22904 5468 22968 5472
rect 22904 5412 22908 5468
rect 22908 5412 22964 5468
rect 22964 5412 22968 5468
rect 22904 5408 22968 5412
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 9094 4924 9158 4928
rect 9094 4868 9098 4924
rect 9098 4868 9154 4924
rect 9154 4868 9158 4924
rect 9094 4864 9158 4868
rect 9174 4924 9238 4928
rect 9174 4868 9178 4924
rect 9178 4868 9234 4924
rect 9234 4868 9238 4924
rect 9174 4864 9238 4868
rect 9254 4924 9318 4928
rect 9254 4868 9258 4924
rect 9258 4868 9314 4924
rect 9314 4868 9318 4924
rect 9254 4864 9318 4868
rect 9334 4924 9398 4928
rect 9334 4868 9338 4924
rect 9338 4868 9394 4924
rect 9394 4868 9398 4924
rect 9334 4864 9398 4868
rect 14522 4924 14586 4928
rect 14522 4868 14526 4924
rect 14526 4868 14582 4924
rect 14582 4868 14586 4924
rect 14522 4864 14586 4868
rect 14602 4924 14666 4928
rect 14602 4868 14606 4924
rect 14606 4868 14662 4924
rect 14662 4868 14666 4924
rect 14602 4864 14666 4868
rect 14682 4924 14746 4928
rect 14682 4868 14686 4924
rect 14686 4868 14742 4924
rect 14742 4868 14746 4924
rect 14682 4864 14746 4868
rect 14762 4924 14826 4928
rect 14762 4868 14766 4924
rect 14766 4868 14822 4924
rect 14822 4868 14826 4924
rect 14762 4864 14826 4868
rect 19950 4924 20014 4928
rect 19950 4868 19954 4924
rect 19954 4868 20010 4924
rect 20010 4868 20014 4924
rect 19950 4864 20014 4868
rect 20030 4924 20094 4928
rect 20030 4868 20034 4924
rect 20034 4868 20090 4924
rect 20090 4868 20094 4924
rect 20030 4864 20094 4868
rect 20110 4924 20174 4928
rect 20110 4868 20114 4924
rect 20114 4868 20170 4924
rect 20170 4868 20174 4924
rect 20110 4864 20174 4868
rect 20190 4924 20254 4928
rect 20190 4868 20194 4924
rect 20194 4868 20250 4924
rect 20250 4868 20254 4924
rect 20190 4864 20254 4868
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 11808 4380 11872 4384
rect 11808 4324 11812 4380
rect 11812 4324 11868 4380
rect 11868 4324 11872 4380
rect 11808 4320 11872 4324
rect 11888 4380 11952 4384
rect 11888 4324 11892 4380
rect 11892 4324 11948 4380
rect 11948 4324 11952 4380
rect 11888 4320 11952 4324
rect 11968 4380 12032 4384
rect 11968 4324 11972 4380
rect 11972 4324 12028 4380
rect 12028 4324 12032 4380
rect 11968 4320 12032 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 17316 4380 17380 4384
rect 17316 4324 17320 4380
rect 17320 4324 17376 4380
rect 17376 4324 17380 4380
rect 17316 4320 17380 4324
rect 17396 4380 17460 4384
rect 17396 4324 17400 4380
rect 17400 4324 17456 4380
rect 17456 4324 17460 4380
rect 17396 4320 17460 4324
rect 17476 4380 17540 4384
rect 17476 4324 17480 4380
rect 17480 4324 17536 4380
rect 17536 4324 17540 4380
rect 17476 4320 17540 4324
rect 22664 4380 22728 4384
rect 22664 4324 22668 4380
rect 22668 4324 22724 4380
rect 22724 4324 22728 4380
rect 22664 4320 22728 4324
rect 22744 4380 22808 4384
rect 22744 4324 22748 4380
rect 22748 4324 22804 4380
rect 22804 4324 22808 4380
rect 22744 4320 22808 4324
rect 22824 4380 22888 4384
rect 22824 4324 22828 4380
rect 22828 4324 22884 4380
rect 22884 4324 22888 4380
rect 22824 4320 22888 4324
rect 22904 4380 22968 4384
rect 22904 4324 22908 4380
rect 22908 4324 22964 4380
rect 22964 4324 22968 4380
rect 22904 4320 22968 4324
rect 19564 3980 19628 4044
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 9094 3836 9158 3840
rect 9094 3780 9098 3836
rect 9098 3780 9154 3836
rect 9154 3780 9158 3836
rect 9094 3776 9158 3780
rect 9174 3836 9238 3840
rect 9174 3780 9178 3836
rect 9178 3780 9234 3836
rect 9234 3780 9238 3836
rect 9174 3776 9238 3780
rect 9254 3836 9318 3840
rect 9254 3780 9258 3836
rect 9258 3780 9314 3836
rect 9314 3780 9318 3836
rect 9254 3776 9318 3780
rect 9334 3836 9398 3840
rect 9334 3780 9338 3836
rect 9338 3780 9394 3836
rect 9394 3780 9398 3836
rect 9334 3776 9398 3780
rect 14522 3836 14586 3840
rect 14522 3780 14526 3836
rect 14526 3780 14582 3836
rect 14582 3780 14586 3836
rect 14522 3776 14586 3780
rect 14602 3836 14666 3840
rect 14602 3780 14606 3836
rect 14606 3780 14662 3836
rect 14662 3780 14666 3836
rect 14602 3776 14666 3780
rect 14682 3836 14746 3840
rect 14682 3780 14686 3836
rect 14686 3780 14742 3836
rect 14742 3780 14746 3836
rect 14682 3776 14746 3780
rect 14762 3836 14826 3840
rect 14762 3780 14766 3836
rect 14766 3780 14822 3836
rect 14822 3780 14826 3836
rect 14762 3776 14826 3780
rect 19950 3836 20014 3840
rect 19950 3780 19954 3836
rect 19954 3780 20010 3836
rect 20010 3780 20014 3836
rect 19950 3776 20014 3780
rect 20030 3836 20094 3840
rect 20030 3780 20034 3836
rect 20034 3780 20090 3836
rect 20090 3780 20094 3836
rect 20030 3776 20094 3780
rect 20110 3836 20174 3840
rect 20110 3780 20114 3836
rect 20114 3780 20170 3836
rect 20170 3780 20174 3836
rect 20110 3776 20174 3780
rect 20190 3836 20254 3840
rect 20190 3780 20194 3836
rect 20194 3780 20250 3836
rect 20250 3780 20254 3836
rect 20190 3776 20254 3780
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 11808 3292 11872 3296
rect 11808 3236 11812 3292
rect 11812 3236 11868 3292
rect 11868 3236 11872 3292
rect 11808 3232 11872 3236
rect 11888 3292 11952 3296
rect 11888 3236 11892 3292
rect 11892 3236 11948 3292
rect 11948 3236 11952 3292
rect 11888 3232 11952 3236
rect 11968 3292 12032 3296
rect 11968 3236 11972 3292
rect 11972 3236 12028 3292
rect 12028 3236 12032 3292
rect 11968 3232 12032 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 17316 3292 17380 3296
rect 17316 3236 17320 3292
rect 17320 3236 17376 3292
rect 17376 3236 17380 3292
rect 17316 3232 17380 3236
rect 17396 3292 17460 3296
rect 17396 3236 17400 3292
rect 17400 3236 17456 3292
rect 17456 3236 17460 3292
rect 17396 3232 17460 3236
rect 17476 3292 17540 3296
rect 17476 3236 17480 3292
rect 17480 3236 17536 3292
rect 17536 3236 17540 3292
rect 17476 3232 17540 3236
rect 22664 3292 22728 3296
rect 22664 3236 22668 3292
rect 22668 3236 22724 3292
rect 22724 3236 22728 3292
rect 22664 3232 22728 3236
rect 22744 3292 22808 3296
rect 22744 3236 22748 3292
rect 22748 3236 22804 3292
rect 22804 3236 22808 3292
rect 22744 3232 22808 3236
rect 22824 3292 22888 3296
rect 22824 3236 22828 3292
rect 22828 3236 22884 3292
rect 22884 3236 22888 3292
rect 22824 3232 22888 3236
rect 22904 3292 22968 3296
rect 22904 3236 22908 3292
rect 22908 3236 22964 3292
rect 22964 3236 22968 3292
rect 22904 3232 22968 3236
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 9094 2748 9158 2752
rect 9094 2692 9098 2748
rect 9098 2692 9154 2748
rect 9154 2692 9158 2748
rect 9094 2688 9158 2692
rect 9174 2748 9238 2752
rect 9174 2692 9178 2748
rect 9178 2692 9234 2748
rect 9234 2692 9238 2748
rect 9174 2688 9238 2692
rect 9254 2748 9318 2752
rect 9254 2692 9258 2748
rect 9258 2692 9314 2748
rect 9314 2692 9318 2748
rect 9254 2688 9318 2692
rect 9334 2748 9398 2752
rect 9334 2692 9338 2748
rect 9338 2692 9394 2748
rect 9394 2692 9398 2748
rect 9334 2688 9398 2692
rect 14522 2748 14586 2752
rect 14522 2692 14526 2748
rect 14526 2692 14582 2748
rect 14582 2692 14586 2748
rect 14522 2688 14586 2692
rect 14602 2748 14666 2752
rect 14602 2692 14606 2748
rect 14606 2692 14662 2748
rect 14662 2692 14666 2748
rect 14602 2688 14666 2692
rect 14682 2748 14746 2752
rect 14682 2692 14686 2748
rect 14686 2692 14742 2748
rect 14742 2692 14746 2748
rect 14682 2688 14746 2692
rect 14762 2748 14826 2752
rect 14762 2692 14766 2748
rect 14766 2692 14822 2748
rect 14822 2692 14826 2748
rect 14762 2688 14826 2692
rect 19950 2748 20014 2752
rect 19950 2692 19954 2748
rect 19954 2692 20010 2748
rect 20010 2692 20014 2748
rect 19950 2688 20014 2692
rect 20030 2748 20094 2752
rect 20030 2692 20034 2748
rect 20034 2692 20090 2748
rect 20090 2692 20094 2748
rect 20030 2688 20094 2692
rect 20110 2748 20174 2752
rect 20110 2692 20114 2748
rect 20114 2692 20170 2748
rect 20170 2692 20174 2748
rect 20110 2688 20174 2692
rect 20190 2748 20254 2752
rect 20190 2692 20194 2748
rect 20194 2692 20250 2748
rect 20250 2692 20254 2748
rect 20190 2688 20254 2692
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 11808 2204 11872 2208
rect 11808 2148 11812 2204
rect 11812 2148 11868 2204
rect 11868 2148 11872 2204
rect 11808 2144 11872 2148
rect 11888 2204 11952 2208
rect 11888 2148 11892 2204
rect 11892 2148 11948 2204
rect 11948 2148 11952 2204
rect 11888 2144 11952 2148
rect 11968 2204 12032 2208
rect 11968 2148 11972 2204
rect 11972 2148 12028 2204
rect 12028 2148 12032 2204
rect 11968 2144 12032 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 17316 2204 17380 2208
rect 17316 2148 17320 2204
rect 17320 2148 17376 2204
rect 17376 2148 17380 2204
rect 17316 2144 17380 2148
rect 17396 2204 17460 2208
rect 17396 2148 17400 2204
rect 17400 2148 17456 2204
rect 17456 2148 17460 2204
rect 17396 2144 17460 2148
rect 17476 2204 17540 2208
rect 17476 2148 17480 2204
rect 17480 2148 17536 2204
rect 17536 2148 17540 2204
rect 17476 2144 17540 2148
rect 22664 2204 22728 2208
rect 22664 2148 22668 2204
rect 22668 2148 22724 2204
rect 22724 2148 22728 2204
rect 22664 2144 22728 2148
rect 22744 2204 22808 2208
rect 22744 2148 22748 2204
rect 22748 2148 22804 2204
rect 22804 2148 22808 2204
rect 22744 2144 22808 2148
rect 22824 2204 22888 2208
rect 22824 2148 22828 2204
rect 22828 2148 22884 2204
rect 22884 2148 22888 2204
rect 22824 2144 22888 2148
rect 22904 2204 22968 2208
rect 22904 2148 22908 2204
rect 22908 2148 22964 2204
rect 22964 2148 22968 2204
rect 22904 2144 22968 2148
<< metal4 >>
rect 3658 21248 3978 21808
rect 3658 21184 3666 21248
rect 3730 21184 3746 21248
rect 3810 21184 3826 21248
rect 3890 21184 3906 21248
rect 3970 21184 3978 21248
rect 3658 20160 3978 21184
rect 3658 20096 3666 20160
rect 3730 20096 3746 20160
rect 3810 20096 3826 20160
rect 3890 20096 3906 20160
rect 3970 20096 3978 20160
rect 3658 19072 3978 20096
rect 3658 19008 3666 19072
rect 3730 19008 3746 19072
rect 3810 19008 3826 19072
rect 3890 19008 3906 19072
rect 3970 19008 3978 19072
rect 3658 17984 3978 19008
rect 3658 17920 3666 17984
rect 3730 17920 3746 17984
rect 3810 17920 3826 17984
rect 3890 17920 3906 17984
rect 3970 17920 3978 17984
rect 3658 16896 3978 17920
rect 3658 16832 3666 16896
rect 3730 16832 3746 16896
rect 3810 16832 3826 16896
rect 3890 16832 3906 16896
rect 3970 16832 3978 16896
rect 3658 15808 3978 16832
rect 3658 15744 3666 15808
rect 3730 15744 3746 15808
rect 3810 15744 3826 15808
rect 3890 15744 3906 15808
rect 3970 15744 3978 15808
rect 3658 14720 3978 15744
rect 3658 14656 3666 14720
rect 3730 14656 3746 14720
rect 3810 14656 3826 14720
rect 3890 14656 3906 14720
rect 3970 14656 3978 14720
rect 3658 13632 3978 14656
rect 3658 13568 3666 13632
rect 3730 13568 3746 13632
rect 3810 13568 3826 13632
rect 3890 13568 3906 13632
rect 3970 13568 3978 13632
rect 3658 12544 3978 13568
rect 3658 12480 3666 12544
rect 3730 12480 3746 12544
rect 3810 12480 3826 12544
rect 3890 12480 3906 12544
rect 3970 12480 3978 12544
rect 3658 11456 3978 12480
rect 3658 11392 3666 11456
rect 3730 11392 3746 11456
rect 3810 11392 3826 11456
rect 3890 11392 3906 11456
rect 3970 11392 3978 11456
rect 3658 10368 3978 11392
rect 3658 10304 3666 10368
rect 3730 10304 3746 10368
rect 3810 10304 3826 10368
rect 3890 10304 3906 10368
rect 3970 10304 3978 10368
rect 3658 9280 3978 10304
rect 3658 9216 3666 9280
rect 3730 9216 3746 9280
rect 3810 9216 3826 9280
rect 3890 9216 3906 9280
rect 3970 9216 3978 9280
rect 3658 8192 3978 9216
rect 3658 8128 3666 8192
rect 3730 8128 3746 8192
rect 3810 8128 3826 8192
rect 3890 8128 3906 8192
rect 3970 8128 3978 8192
rect 3658 7104 3978 8128
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6016 3978 7040
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4928 3978 5952
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 3840 3978 4864
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 2752 3978 3776
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 6372 21792 6692 21808
rect 6372 21728 6380 21792
rect 6444 21728 6460 21792
rect 6524 21728 6540 21792
rect 6604 21728 6620 21792
rect 6684 21728 6692 21792
rect 6372 20704 6692 21728
rect 6372 20640 6380 20704
rect 6444 20640 6460 20704
rect 6524 20640 6540 20704
rect 6604 20640 6620 20704
rect 6684 20640 6692 20704
rect 6372 19616 6692 20640
rect 6372 19552 6380 19616
rect 6444 19552 6460 19616
rect 6524 19552 6540 19616
rect 6604 19552 6620 19616
rect 6684 19552 6692 19616
rect 6372 18528 6692 19552
rect 6372 18464 6380 18528
rect 6444 18464 6460 18528
rect 6524 18464 6540 18528
rect 6604 18464 6620 18528
rect 6684 18464 6692 18528
rect 6372 17440 6692 18464
rect 6372 17376 6380 17440
rect 6444 17376 6460 17440
rect 6524 17376 6540 17440
rect 6604 17376 6620 17440
rect 6684 17376 6692 17440
rect 6372 16352 6692 17376
rect 6372 16288 6380 16352
rect 6444 16288 6460 16352
rect 6524 16288 6540 16352
rect 6604 16288 6620 16352
rect 6684 16288 6692 16352
rect 6372 15264 6692 16288
rect 6372 15200 6380 15264
rect 6444 15200 6460 15264
rect 6524 15200 6540 15264
rect 6604 15200 6620 15264
rect 6684 15200 6692 15264
rect 6372 14176 6692 15200
rect 6372 14112 6380 14176
rect 6444 14112 6460 14176
rect 6524 14112 6540 14176
rect 6604 14112 6620 14176
rect 6684 14112 6692 14176
rect 6372 13088 6692 14112
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 5472 6692 6496
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 9086 21248 9406 21808
rect 9086 21184 9094 21248
rect 9158 21184 9174 21248
rect 9238 21184 9254 21248
rect 9318 21184 9334 21248
rect 9398 21184 9406 21248
rect 9086 20160 9406 21184
rect 9086 20096 9094 20160
rect 9158 20096 9174 20160
rect 9238 20096 9254 20160
rect 9318 20096 9334 20160
rect 9398 20096 9406 20160
rect 9086 19072 9406 20096
rect 9086 19008 9094 19072
rect 9158 19008 9174 19072
rect 9238 19008 9254 19072
rect 9318 19008 9334 19072
rect 9398 19008 9406 19072
rect 9086 17984 9406 19008
rect 9086 17920 9094 17984
rect 9158 17920 9174 17984
rect 9238 17920 9254 17984
rect 9318 17920 9334 17984
rect 9398 17920 9406 17984
rect 9086 16896 9406 17920
rect 9086 16832 9094 16896
rect 9158 16832 9174 16896
rect 9238 16832 9254 16896
rect 9318 16832 9334 16896
rect 9398 16832 9406 16896
rect 9086 15808 9406 16832
rect 9086 15744 9094 15808
rect 9158 15744 9174 15808
rect 9238 15744 9254 15808
rect 9318 15744 9334 15808
rect 9398 15744 9406 15808
rect 9086 14720 9406 15744
rect 9086 14656 9094 14720
rect 9158 14656 9174 14720
rect 9238 14656 9254 14720
rect 9318 14656 9334 14720
rect 9398 14656 9406 14720
rect 9086 13632 9406 14656
rect 9086 13568 9094 13632
rect 9158 13568 9174 13632
rect 9238 13568 9254 13632
rect 9318 13568 9334 13632
rect 9398 13568 9406 13632
rect 9086 12544 9406 13568
rect 9086 12480 9094 12544
rect 9158 12480 9174 12544
rect 9238 12480 9254 12544
rect 9318 12480 9334 12544
rect 9398 12480 9406 12544
rect 9086 11456 9406 12480
rect 9086 11392 9094 11456
rect 9158 11392 9174 11456
rect 9238 11392 9254 11456
rect 9318 11392 9334 11456
rect 9398 11392 9406 11456
rect 9086 10368 9406 11392
rect 9086 10304 9094 10368
rect 9158 10304 9174 10368
rect 9238 10304 9254 10368
rect 9318 10304 9334 10368
rect 9398 10304 9406 10368
rect 9086 9280 9406 10304
rect 9086 9216 9094 9280
rect 9158 9216 9174 9280
rect 9238 9216 9254 9280
rect 9318 9216 9334 9280
rect 9398 9216 9406 9280
rect 9086 8192 9406 9216
rect 9086 8128 9094 8192
rect 9158 8128 9174 8192
rect 9238 8128 9254 8192
rect 9318 8128 9334 8192
rect 9398 8128 9406 8192
rect 9086 7104 9406 8128
rect 9086 7040 9094 7104
rect 9158 7040 9174 7104
rect 9238 7040 9254 7104
rect 9318 7040 9334 7104
rect 9398 7040 9406 7104
rect 9086 6016 9406 7040
rect 9086 5952 9094 6016
rect 9158 5952 9174 6016
rect 9238 5952 9254 6016
rect 9318 5952 9334 6016
rect 9398 5952 9406 6016
rect 9086 4928 9406 5952
rect 9086 4864 9094 4928
rect 9158 4864 9174 4928
rect 9238 4864 9254 4928
rect 9318 4864 9334 4928
rect 9398 4864 9406 4928
rect 9086 3840 9406 4864
rect 9086 3776 9094 3840
rect 9158 3776 9174 3840
rect 9238 3776 9254 3840
rect 9318 3776 9334 3840
rect 9398 3776 9406 3840
rect 9086 2752 9406 3776
rect 9086 2688 9094 2752
rect 9158 2688 9174 2752
rect 9238 2688 9254 2752
rect 9318 2688 9334 2752
rect 9398 2688 9406 2752
rect 9086 2128 9406 2688
rect 11800 21792 12120 21808
rect 11800 21728 11808 21792
rect 11872 21728 11888 21792
rect 11952 21728 11968 21792
rect 12032 21728 12048 21792
rect 12112 21728 12120 21792
rect 11800 20704 12120 21728
rect 11800 20640 11808 20704
rect 11872 20640 11888 20704
rect 11952 20640 11968 20704
rect 12032 20640 12048 20704
rect 12112 20640 12120 20704
rect 11800 19616 12120 20640
rect 11800 19552 11808 19616
rect 11872 19552 11888 19616
rect 11952 19552 11968 19616
rect 12032 19552 12048 19616
rect 12112 19552 12120 19616
rect 11800 18528 12120 19552
rect 11800 18464 11808 18528
rect 11872 18464 11888 18528
rect 11952 18464 11968 18528
rect 12032 18464 12048 18528
rect 12112 18464 12120 18528
rect 11800 17440 12120 18464
rect 11800 17376 11808 17440
rect 11872 17376 11888 17440
rect 11952 17376 11968 17440
rect 12032 17376 12048 17440
rect 12112 17376 12120 17440
rect 11800 16352 12120 17376
rect 11800 16288 11808 16352
rect 11872 16288 11888 16352
rect 11952 16288 11968 16352
rect 12032 16288 12048 16352
rect 12112 16288 12120 16352
rect 11800 15264 12120 16288
rect 11800 15200 11808 15264
rect 11872 15200 11888 15264
rect 11952 15200 11968 15264
rect 12032 15200 12048 15264
rect 12112 15200 12120 15264
rect 11800 14176 12120 15200
rect 11800 14112 11808 14176
rect 11872 14112 11888 14176
rect 11952 14112 11968 14176
rect 12032 14112 12048 14176
rect 12112 14112 12120 14176
rect 11800 13088 12120 14112
rect 11800 13024 11808 13088
rect 11872 13024 11888 13088
rect 11952 13024 11968 13088
rect 12032 13024 12048 13088
rect 12112 13024 12120 13088
rect 11800 12000 12120 13024
rect 11800 11936 11808 12000
rect 11872 11936 11888 12000
rect 11952 11936 11968 12000
rect 12032 11936 12048 12000
rect 12112 11936 12120 12000
rect 11800 10912 12120 11936
rect 11800 10848 11808 10912
rect 11872 10848 11888 10912
rect 11952 10848 11968 10912
rect 12032 10848 12048 10912
rect 12112 10848 12120 10912
rect 11800 9824 12120 10848
rect 11800 9760 11808 9824
rect 11872 9760 11888 9824
rect 11952 9760 11968 9824
rect 12032 9760 12048 9824
rect 12112 9760 12120 9824
rect 11800 8736 12120 9760
rect 11800 8672 11808 8736
rect 11872 8672 11888 8736
rect 11952 8672 11968 8736
rect 12032 8672 12048 8736
rect 12112 8672 12120 8736
rect 11800 7648 12120 8672
rect 11800 7584 11808 7648
rect 11872 7584 11888 7648
rect 11952 7584 11968 7648
rect 12032 7584 12048 7648
rect 12112 7584 12120 7648
rect 11800 6560 12120 7584
rect 11800 6496 11808 6560
rect 11872 6496 11888 6560
rect 11952 6496 11968 6560
rect 12032 6496 12048 6560
rect 12112 6496 12120 6560
rect 11800 5472 12120 6496
rect 11800 5408 11808 5472
rect 11872 5408 11888 5472
rect 11952 5408 11968 5472
rect 12032 5408 12048 5472
rect 12112 5408 12120 5472
rect 11800 4384 12120 5408
rect 11800 4320 11808 4384
rect 11872 4320 11888 4384
rect 11952 4320 11968 4384
rect 12032 4320 12048 4384
rect 12112 4320 12120 4384
rect 11800 3296 12120 4320
rect 11800 3232 11808 3296
rect 11872 3232 11888 3296
rect 11952 3232 11968 3296
rect 12032 3232 12048 3296
rect 12112 3232 12120 3296
rect 11800 2208 12120 3232
rect 11800 2144 11808 2208
rect 11872 2144 11888 2208
rect 11952 2144 11968 2208
rect 12032 2144 12048 2208
rect 12112 2144 12120 2208
rect 11800 2128 12120 2144
rect 14514 21248 14834 21808
rect 14514 21184 14522 21248
rect 14586 21184 14602 21248
rect 14666 21184 14682 21248
rect 14746 21184 14762 21248
rect 14826 21184 14834 21248
rect 14514 20160 14834 21184
rect 14514 20096 14522 20160
rect 14586 20096 14602 20160
rect 14666 20096 14682 20160
rect 14746 20096 14762 20160
rect 14826 20096 14834 20160
rect 14514 19072 14834 20096
rect 14514 19008 14522 19072
rect 14586 19008 14602 19072
rect 14666 19008 14682 19072
rect 14746 19008 14762 19072
rect 14826 19008 14834 19072
rect 14514 17984 14834 19008
rect 14514 17920 14522 17984
rect 14586 17920 14602 17984
rect 14666 17920 14682 17984
rect 14746 17920 14762 17984
rect 14826 17920 14834 17984
rect 14514 16896 14834 17920
rect 14514 16832 14522 16896
rect 14586 16832 14602 16896
rect 14666 16832 14682 16896
rect 14746 16832 14762 16896
rect 14826 16832 14834 16896
rect 14514 15808 14834 16832
rect 14514 15744 14522 15808
rect 14586 15744 14602 15808
rect 14666 15744 14682 15808
rect 14746 15744 14762 15808
rect 14826 15744 14834 15808
rect 14514 14720 14834 15744
rect 14514 14656 14522 14720
rect 14586 14656 14602 14720
rect 14666 14656 14682 14720
rect 14746 14656 14762 14720
rect 14826 14656 14834 14720
rect 14514 13632 14834 14656
rect 14514 13568 14522 13632
rect 14586 13568 14602 13632
rect 14666 13568 14682 13632
rect 14746 13568 14762 13632
rect 14826 13568 14834 13632
rect 14514 12544 14834 13568
rect 14514 12480 14522 12544
rect 14586 12480 14602 12544
rect 14666 12480 14682 12544
rect 14746 12480 14762 12544
rect 14826 12480 14834 12544
rect 14514 11456 14834 12480
rect 14514 11392 14522 11456
rect 14586 11392 14602 11456
rect 14666 11392 14682 11456
rect 14746 11392 14762 11456
rect 14826 11392 14834 11456
rect 14514 10368 14834 11392
rect 17228 21792 17548 21808
rect 17228 21728 17236 21792
rect 17300 21728 17316 21792
rect 17380 21728 17396 21792
rect 17460 21728 17476 21792
rect 17540 21728 17548 21792
rect 17228 20704 17548 21728
rect 17228 20640 17236 20704
rect 17300 20640 17316 20704
rect 17380 20640 17396 20704
rect 17460 20640 17476 20704
rect 17540 20640 17548 20704
rect 17228 19616 17548 20640
rect 17228 19552 17236 19616
rect 17300 19552 17316 19616
rect 17380 19552 17396 19616
rect 17460 19552 17476 19616
rect 17540 19552 17548 19616
rect 17228 18528 17548 19552
rect 17228 18464 17236 18528
rect 17300 18464 17316 18528
rect 17380 18464 17396 18528
rect 17460 18464 17476 18528
rect 17540 18464 17548 18528
rect 17228 17440 17548 18464
rect 17228 17376 17236 17440
rect 17300 17376 17316 17440
rect 17380 17376 17396 17440
rect 17460 17376 17476 17440
rect 17540 17376 17548 17440
rect 17228 16352 17548 17376
rect 17228 16288 17236 16352
rect 17300 16288 17316 16352
rect 17380 16288 17396 16352
rect 17460 16288 17476 16352
rect 17540 16288 17548 16352
rect 17228 15264 17548 16288
rect 17228 15200 17236 15264
rect 17300 15200 17316 15264
rect 17380 15200 17396 15264
rect 17460 15200 17476 15264
rect 17540 15200 17548 15264
rect 17228 14176 17548 15200
rect 17228 14112 17236 14176
rect 17300 14112 17316 14176
rect 17380 14112 17396 14176
rect 17460 14112 17476 14176
rect 17540 14112 17548 14176
rect 17228 13088 17548 14112
rect 17228 13024 17236 13088
rect 17300 13024 17316 13088
rect 17380 13024 17396 13088
rect 17460 13024 17476 13088
rect 17540 13024 17548 13088
rect 17228 12000 17548 13024
rect 17228 11936 17236 12000
rect 17300 11936 17316 12000
rect 17380 11936 17396 12000
rect 17460 11936 17476 12000
rect 17540 11936 17548 12000
rect 17228 10912 17548 11936
rect 17228 10848 17236 10912
rect 17300 10848 17316 10912
rect 17380 10848 17396 10912
rect 17460 10848 17476 10912
rect 17540 10848 17548 10912
rect 15147 10572 15213 10573
rect 15147 10508 15148 10572
rect 15212 10508 15213 10572
rect 15147 10507 15213 10508
rect 14514 10304 14522 10368
rect 14586 10304 14602 10368
rect 14666 10304 14682 10368
rect 14746 10304 14762 10368
rect 14826 10304 14834 10368
rect 14514 9280 14834 10304
rect 14514 9216 14522 9280
rect 14586 9216 14602 9280
rect 14666 9216 14682 9280
rect 14746 9216 14762 9280
rect 14826 9216 14834 9280
rect 14514 8192 14834 9216
rect 14514 8128 14522 8192
rect 14586 8128 14602 8192
rect 14666 8128 14682 8192
rect 14746 8128 14762 8192
rect 14826 8128 14834 8192
rect 14514 7104 14834 8128
rect 14514 7040 14522 7104
rect 14586 7040 14602 7104
rect 14666 7040 14682 7104
rect 14746 7040 14762 7104
rect 14826 7040 14834 7104
rect 14514 6016 14834 7040
rect 15150 6765 15210 10507
rect 17228 9824 17548 10848
rect 17228 9760 17236 9824
rect 17300 9760 17316 9824
rect 17380 9760 17396 9824
rect 17460 9760 17476 9824
rect 17540 9760 17548 9824
rect 17228 8736 17548 9760
rect 17228 8672 17236 8736
rect 17300 8672 17316 8736
rect 17380 8672 17396 8736
rect 17460 8672 17476 8736
rect 17540 8672 17548 8736
rect 17228 7648 17548 8672
rect 17228 7584 17236 7648
rect 17300 7584 17316 7648
rect 17380 7584 17396 7648
rect 17460 7584 17476 7648
rect 17540 7584 17548 7648
rect 15147 6764 15213 6765
rect 15147 6700 15148 6764
rect 15212 6700 15213 6764
rect 15147 6699 15213 6700
rect 14514 5952 14522 6016
rect 14586 5952 14602 6016
rect 14666 5952 14682 6016
rect 14746 5952 14762 6016
rect 14826 5952 14834 6016
rect 14514 4928 14834 5952
rect 14514 4864 14522 4928
rect 14586 4864 14602 4928
rect 14666 4864 14682 4928
rect 14746 4864 14762 4928
rect 14826 4864 14834 4928
rect 14514 3840 14834 4864
rect 14514 3776 14522 3840
rect 14586 3776 14602 3840
rect 14666 3776 14682 3840
rect 14746 3776 14762 3840
rect 14826 3776 14834 3840
rect 14514 2752 14834 3776
rect 14514 2688 14522 2752
rect 14586 2688 14602 2752
rect 14666 2688 14682 2752
rect 14746 2688 14762 2752
rect 14826 2688 14834 2752
rect 14514 2128 14834 2688
rect 17228 6560 17548 7584
rect 17228 6496 17236 6560
rect 17300 6496 17316 6560
rect 17380 6496 17396 6560
rect 17460 6496 17476 6560
rect 17540 6496 17548 6560
rect 17228 5472 17548 6496
rect 19942 21248 20262 21808
rect 19942 21184 19950 21248
rect 20014 21184 20030 21248
rect 20094 21184 20110 21248
rect 20174 21184 20190 21248
rect 20254 21184 20262 21248
rect 19942 20160 20262 21184
rect 19942 20096 19950 20160
rect 20014 20096 20030 20160
rect 20094 20096 20110 20160
rect 20174 20096 20190 20160
rect 20254 20096 20262 20160
rect 19942 19072 20262 20096
rect 19942 19008 19950 19072
rect 20014 19008 20030 19072
rect 20094 19008 20110 19072
rect 20174 19008 20190 19072
rect 20254 19008 20262 19072
rect 19942 17984 20262 19008
rect 19942 17920 19950 17984
rect 20014 17920 20030 17984
rect 20094 17920 20110 17984
rect 20174 17920 20190 17984
rect 20254 17920 20262 17984
rect 19942 16896 20262 17920
rect 19942 16832 19950 16896
rect 20014 16832 20030 16896
rect 20094 16832 20110 16896
rect 20174 16832 20190 16896
rect 20254 16832 20262 16896
rect 19942 15808 20262 16832
rect 19942 15744 19950 15808
rect 20014 15744 20030 15808
rect 20094 15744 20110 15808
rect 20174 15744 20190 15808
rect 20254 15744 20262 15808
rect 19942 14720 20262 15744
rect 19942 14656 19950 14720
rect 20014 14656 20030 14720
rect 20094 14656 20110 14720
rect 20174 14656 20190 14720
rect 20254 14656 20262 14720
rect 19942 13632 20262 14656
rect 19942 13568 19950 13632
rect 20014 13568 20030 13632
rect 20094 13568 20110 13632
rect 20174 13568 20190 13632
rect 20254 13568 20262 13632
rect 19942 12544 20262 13568
rect 19942 12480 19950 12544
rect 20014 12480 20030 12544
rect 20094 12480 20110 12544
rect 20174 12480 20190 12544
rect 20254 12480 20262 12544
rect 19942 11456 20262 12480
rect 19942 11392 19950 11456
rect 20014 11392 20030 11456
rect 20094 11392 20110 11456
rect 20174 11392 20190 11456
rect 20254 11392 20262 11456
rect 19942 10368 20262 11392
rect 19942 10304 19950 10368
rect 20014 10304 20030 10368
rect 20094 10304 20110 10368
rect 20174 10304 20190 10368
rect 20254 10304 20262 10368
rect 19942 9280 20262 10304
rect 19942 9216 19950 9280
rect 20014 9216 20030 9280
rect 20094 9216 20110 9280
rect 20174 9216 20190 9280
rect 20254 9216 20262 9280
rect 19942 8192 20262 9216
rect 19942 8128 19950 8192
rect 20014 8128 20030 8192
rect 20094 8128 20110 8192
rect 20174 8128 20190 8192
rect 20254 8128 20262 8192
rect 19942 7104 20262 8128
rect 19942 7040 19950 7104
rect 20014 7040 20030 7104
rect 20094 7040 20110 7104
rect 20174 7040 20190 7104
rect 20254 7040 20262 7104
rect 19942 6016 20262 7040
rect 19942 5952 19950 6016
rect 20014 5952 20030 6016
rect 20094 5952 20110 6016
rect 20174 5952 20190 6016
rect 20254 5952 20262 6016
rect 19563 5676 19629 5677
rect 19563 5612 19564 5676
rect 19628 5612 19629 5676
rect 19563 5611 19629 5612
rect 17228 5408 17236 5472
rect 17300 5408 17316 5472
rect 17380 5408 17396 5472
rect 17460 5408 17476 5472
rect 17540 5408 17548 5472
rect 17228 4384 17548 5408
rect 17228 4320 17236 4384
rect 17300 4320 17316 4384
rect 17380 4320 17396 4384
rect 17460 4320 17476 4384
rect 17540 4320 17548 4384
rect 17228 3296 17548 4320
rect 19566 4045 19626 5611
rect 19942 4928 20262 5952
rect 19942 4864 19950 4928
rect 20014 4864 20030 4928
rect 20094 4864 20110 4928
rect 20174 4864 20190 4928
rect 20254 4864 20262 4928
rect 19563 4044 19629 4045
rect 19563 3980 19564 4044
rect 19628 3980 19629 4044
rect 19563 3979 19629 3980
rect 17228 3232 17236 3296
rect 17300 3232 17316 3296
rect 17380 3232 17396 3296
rect 17460 3232 17476 3296
rect 17540 3232 17548 3296
rect 17228 2208 17548 3232
rect 17228 2144 17236 2208
rect 17300 2144 17316 2208
rect 17380 2144 17396 2208
rect 17460 2144 17476 2208
rect 17540 2144 17548 2208
rect 17228 2128 17548 2144
rect 19942 3840 20262 4864
rect 19942 3776 19950 3840
rect 20014 3776 20030 3840
rect 20094 3776 20110 3840
rect 20174 3776 20190 3840
rect 20254 3776 20262 3840
rect 19942 2752 20262 3776
rect 19942 2688 19950 2752
rect 20014 2688 20030 2752
rect 20094 2688 20110 2752
rect 20174 2688 20190 2752
rect 20254 2688 20262 2752
rect 19942 2128 20262 2688
rect 22656 21792 22976 21808
rect 22656 21728 22664 21792
rect 22728 21728 22744 21792
rect 22808 21728 22824 21792
rect 22888 21728 22904 21792
rect 22968 21728 22976 21792
rect 22656 20704 22976 21728
rect 22656 20640 22664 20704
rect 22728 20640 22744 20704
rect 22808 20640 22824 20704
rect 22888 20640 22904 20704
rect 22968 20640 22976 20704
rect 22656 19616 22976 20640
rect 22656 19552 22664 19616
rect 22728 19552 22744 19616
rect 22808 19552 22824 19616
rect 22888 19552 22904 19616
rect 22968 19552 22976 19616
rect 22656 18528 22976 19552
rect 22656 18464 22664 18528
rect 22728 18464 22744 18528
rect 22808 18464 22824 18528
rect 22888 18464 22904 18528
rect 22968 18464 22976 18528
rect 22656 17440 22976 18464
rect 22656 17376 22664 17440
rect 22728 17376 22744 17440
rect 22808 17376 22824 17440
rect 22888 17376 22904 17440
rect 22968 17376 22976 17440
rect 22656 16352 22976 17376
rect 22656 16288 22664 16352
rect 22728 16288 22744 16352
rect 22808 16288 22824 16352
rect 22888 16288 22904 16352
rect 22968 16288 22976 16352
rect 22656 15264 22976 16288
rect 22656 15200 22664 15264
rect 22728 15200 22744 15264
rect 22808 15200 22824 15264
rect 22888 15200 22904 15264
rect 22968 15200 22976 15264
rect 22656 14176 22976 15200
rect 22656 14112 22664 14176
rect 22728 14112 22744 14176
rect 22808 14112 22824 14176
rect 22888 14112 22904 14176
rect 22968 14112 22976 14176
rect 22656 13088 22976 14112
rect 22656 13024 22664 13088
rect 22728 13024 22744 13088
rect 22808 13024 22824 13088
rect 22888 13024 22904 13088
rect 22968 13024 22976 13088
rect 22656 12000 22976 13024
rect 22656 11936 22664 12000
rect 22728 11936 22744 12000
rect 22808 11936 22824 12000
rect 22888 11936 22904 12000
rect 22968 11936 22976 12000
rect 22656 10912 22976 11936
rect 22656 10848 22664 10912
rect 22728 10848 22744 10912
rect 22808 10848 22824 10912
rect 22888 10848 22904 10912
rect 22968 10848 22976 10912
rect 22656 9824 22976 10848
rect 22656 9760 22664 9824
rect 22728 9760 22744 9824
rect 22808 9760 22824 9824
rect 22888 9760 22904 9824
rect 22968 9760 22976 9824
rect 22656 8736 22976 9760
rect 22656 8672 22664 8736
rect 22728 8672 22744 8736
rect 22808 8672 22824 8736
rect 22888 8672 22904 8736
rect 22968 8672 22976 8736
rect 22656 7648 22976 8672
rect 22656 7584 22664 7648
rect 22728 7584 22744 7648
rect 22808 7584 22824 7648
rect 22888 7584 22904 7648
rect 22968 7584 22976 7648
rect 22656 6560 22976 7584
rect 22656 6496 22664 6560
rect 22728 6496 22744 6560
rect 22808 6496 22824 6560
rect 22888 6496 22904 6560
rect 22968 6496 22976 6560
rect 22656 5472 22976 6496
rect 22656 5408 22664 5472
rect 22728 5408 22744 5472
rect 22808 5408 22824 5472
rect 22888 5408 22904 5472
rect 22968 5408 22976 5472
rect 22656 4384 22976 5408
rect 22656 4320 22664 4384
rect 22728 4320 22744 4384
rect 22808 4320 22824 4384
rect 22888 4320 22904 4384
rect 22968 4320 22976 4384
rect 22656 3296 22976 4320
rect 22656 3232 22664 3296
rect 22728 3232 22744 3296
rect 22808 3232 22824 3296
rect 22888 3232 22904 3296
rect 22968 3232 22976 3296
rect 22656 2208 22976 3232
rect 22656 2144 22664 2208
rect 22728 2144 22744 2208
rect 22808 2144 22824 2208
rect 22888 2144 22904 2208
rect 22968 2144 22976 2208
rect 22656 2128 22976 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666464484
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1666464484
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A
timestamp 1666464484
transform -1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1666464484
transform -1 0 15272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666464484
transform -1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1666464484
transform -1 0 17848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__B
timestamp 1666464484
transform -1 0 21160 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1666464484
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1666464484
transform -1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1666464484
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1666464484
transform 1 0 4600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__C1
timestamp 1666464484
transform 1 0 5152 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__S
timestamp 1666464484
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__B1
timestamp 1666464484
transform 1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1666464484
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__D
timestamp 1666464484
transform 1 0 4968 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1666464484
transform -1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1666464484
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1666464484
transform 1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5152 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71
timestamp 1666464484
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1666464484
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1666464484
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93
timestamp 1666464484
transform 1 0 9660 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 1666464484
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666464484
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_120
timestamp 1666464484
transform 1 0 12144 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1666464484
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_132
timestamp 1666464484
transform 1 0 13248 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_149
timestamp 1666464484
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_154
timestamp 1666464484
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1666464484
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1666464484
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1666464484
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1666464484
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1666464484
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1666464484
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_122
timestamp 1666464484
transform 1 0 12328 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_135
timestamp 1666464484
transform 1 0 13524 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp 1666464484
transform 1 0 14260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1666464484
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1666464484
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_176
timestamp 1666464484
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_182
timestamp 1666464484
transform 1 0 17848 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1666464484
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_203
timestamp 1666464484
transform 1 0 19780 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1666464484
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1666464484
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_49
timestamp 1666464484
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1666464484
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1666464484
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1666464484
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_112
timestamp 1666464484
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_116
timestamp 1666464484
transform 1 0 11776 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1666464484
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1666464484
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_149
timestamp 1666464484
transform 1 0 14812 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1666464484
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp 1666464484
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1666464484
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666464484
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1666464484
transform 1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_212
timestamp 1666464484
transform 1 0 20608 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_218
timestamp 1666464484
transform 1 0 21160 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_230
timestamp 1666464484
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp 1666464484
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_30
timestamp 1666464484
transform 1 0 3864 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1666464484
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1666464484
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1666464484
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1666464484
transform 1 0 12420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_134
timestamp 1666464484
transform 1 0 13432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1666464484
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_151
timestamp 1666464484
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1666464484
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1666464484
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_204
timestamp 1666464484
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1666464484
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1666464484
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1666464484
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1666464484
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1666464484
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_151
timestamp 1666464484
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_155
timestamp 1666464484
transform 1 0 15364 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1666464484
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1666464484
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1666464484
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1666464484
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_185
timestamp 1666464484
transform 1 0 18124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_202
timestamp 1666464484
transform 1 0 19688 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_214
timestamp 1666464484
transform 1 0 20792 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_226
timestamp 1666464484
transform 1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_232
timestamp 1666464484
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1666464484
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1666464484
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1666464484
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1666464484
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1666464484
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_68
timestamp 1666464484
transform 1 0 7360 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1666464484
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1666464484
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1666464484
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp 1666464484
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_140
timestamp 1666464484
transform 1 0 13984 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_150
timestamp 1666464484
transform 1 0 14904 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1666464484
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_173
timestamp 1666464484
transform 1 0 17020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_182
timestamp 1666464484
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1666464484
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1666464484
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1666464484
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_113
timestamp 1666464484
transform 1 0 11500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1666464484
transform 1 0 12328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1666464484
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_152
timestamp 1666464484
transform 1 0 15088 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_167
timestamp 1666464484
transform 1 0 16468 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_174
timestamp 1666464484
transform 1 0 17112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1666464484
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1666464484
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_219
timestamp 1666464484
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_231
timestamp 1666464484
transform 1 0 22356 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_21
timestamp 1666464484
transform 1 0 3036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_28
timestamp 1666464484
transform 1 0 3680 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1666464484
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1666464484
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_65
timestamp 1666464484
transform 1 0 7084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_71
timestamp 1666464484
transform 1 0 7636 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_89
timestamp 1666464484
transform 1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1666464484
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1666464484
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_145
timestamp 1666464484
transform 1 0 14444 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1666464484
transform 1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1666464484
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_179
timestamp 1666464484
transform 1 0 17572 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_187
timestamp 1666464484
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_197
timestamp 1666464484
transform 1 0 19228 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1666464484
transform 1 0 20424 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1666464484
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1666464484
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_44
timestamp 1666464484
transform 1 0 5152 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_72
timestamp 1666464484
transform 1 0 7728 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1666464484
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1666464484
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_110
timestamp 1666464484
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_122
timestamp 1666464484
transform 1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_128
timestamp 1666464484
transform 1 0 12880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_146
timestamp 1666464484
transform 1 0 14536 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1666464484
transform 1 0 15272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_161
timestamp 1666464484
transform 1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_168
timestamp 1666464484
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1666464484
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1666464484
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_206
timestamp 1666464484
transform 1 0 20056 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_218
timestamp 1666464484
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp 1666464484
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1666464484
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_36
timestamp 1666464484
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1666464484
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1666464484
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_68
timestamp 1666464484
transform 1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_72
timestamp 1666464484
transform 1 0 7728 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1666464484
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_142
timestamp 1666464484
transform 1 0 14168 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_150
timestamp 1666464484
transform 1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1666464484
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1666464484
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1666464484
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_195
timestamp 1666464484
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_203
timestamp 1666464484
transform 1 0 19780 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_210
timestamp 1666464484
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1666464484
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1666464484
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1666464484
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1666464484
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1666464484
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_114
timestamp 1666464484
transform 1 0 11592 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1666464484
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1666464484
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1666464484
transform 1 0 14628 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1666464484
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_171
timestamp 1666464484
transform 1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_184
timestamp 1666464484
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1666464484
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_203
timestamp 1666464484
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_210
timestamp 1666464484
transform 1 0 20424 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_222
timestamp 1666464484
transform 1 0 21528 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp 1666464484
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1666464484
transform 1 0 2116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_28
timestamp 1666464484
transform 1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_35
timestamp 1666464484
transform 1 0 4324 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1666464484
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1666464484
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_85
timestamp 1666464484
transform 1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1666464484
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1666464484
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_143
timestamp 1666464484
transform 1 0 14260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_152
timestamp 1666464484
transform 1 0 15088 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_158
timestamp 1666464484
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1666464484
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1666464484
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1666464484
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1666464484
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_210
timestamp 1666464484
transform 1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_47
timestamp 1666464484
transform 1 0 5428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_59
timestamp 1666464484
transform 1 0 6532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_114
timestamp 1666464484
transform 1 0 11592 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_129
timestamp 1666464484
transform 1 0 12972 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1666464484
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_172
timestamp 1666464484
transform 1 0 16928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_176
timestamp 1666464484
transform 1 0 17296 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1666464484
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_188
timestamp 1666464484
transform 1 0 18400 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_204
timestamp 1666464484
transform 1 0 19872 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_216
timestamp 1666464484
transform 1 0 20976 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1666464484
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_232
timestamp 1666464484
transform 1 0 22448 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_21
timestamp 1666464484
transform 1 0 3036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1666464484
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1666464484
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_77
timestamp 1666464484
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_94
timestamp 1666464484
transform 1 0 9752 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1666464484
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1666464484
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_148
timestamp 1666464484
transform 1 0 14720 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1666464484
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_177
timestamp 1666464484
transform 1 0 17388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_189
timestamp 1666464484
transform 1 0 18492 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_201
timestamp 1666464484
transform 1 0 19596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1666464484
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1666464484
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1666464484
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1666464484
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_71
timestamp 1666464484
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_114
timestamp 1666464484
transform 1 0 11592 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_126
timestamp 1666464484
transform 1 0 12696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1666464484
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_151
timestamp 1666464484
transform 1 0 14996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1666464484
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1666464484
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1666464484
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_21
timestamp 1666464484
transform 1 0 3036 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_41
timestamp 1666464484
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1666464484
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1666464484
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_86
timestamp 1666464484
transform 1 0 9016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1666464484
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_120
timestamp 1666464484
transform 1 0 12144 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1666464484
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1666464484
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1666464484
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_11
timestamp 1666464484
transform 1 0 2116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1666464484
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_38
timestamp 1666464484
transform 1 0 4600 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_45
timestamp 1666464484
transform 1 0 5244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1666464484
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1666464484
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_73
timestamp 1666464484
transform 1 0 7820 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1666464484
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1666464484
transform 1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1666464484
transform 1 0 11408 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1666464484
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1666464484
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_146
timestamp 1666464484
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_158
timestamp 1666464484
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_170
timestamp 1666464484
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_182
timestamp 1666464484
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1666464484
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1666464484
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_21
timestamp 1666464484
transform 1 0 3036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_35
timestamp 1666464484
transform 1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1666464484
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1666464484
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_70
timestamp 1666464484
transform 1 0 7544 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1666464484
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_97
timestamp 1666464484
transform 1 0 10028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1666464484
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_122
timestamp 1666464484
transform 1 0 12328 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_134
timestamp 1666464484
transform 1 0 13432 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1666464484
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_151
timestamp 1666464484
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1666464484
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1666464484
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1666464484
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1666464484
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_39
timestamp 1666464484
transform 1 0 4692 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_43
timestamp 1666464484
transform 1 0 5060 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_61
timestamp 1666464484
transform 1 0 6716 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_72
timestamp 1666464484
transform 1 0 7728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1666464484
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_94
timestamp 1666464484
transform 1 0 9752 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_103
timestamp 1666464484
transform 1 0 10580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_116
timestamp 1666464484
transform 1 0 11776 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_122
timestamp 1666464484
transform 1 0 12328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_151
timestamp 1666464484
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_163
timestamp 1666464484
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_175
timestamp 1666464484
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1666464484
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1666464484
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1666464484
transform 1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_23
timestamp 1666464484
transform 1 0 3220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1666464484
transform 1 0 4324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1666464484
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1666464484
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_76
timestamp 1666464484
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_84
timestamp 1666464484
transform 1 0 8832 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1666464484
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_101
timestamp 1666464484
transform 1 0 10396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1666464484
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_127
timestamp 1666464484
transform 1 0 12788 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1666464484
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_145
timestamp 1666464484
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1666464484
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1666464484
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_20
timestamp 1666464484
transform 1 0 2944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1666464484
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1666464484
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_46
timestamp 1666464484
transform 1 0 5336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_54
timestamp 1666464484
transform 1 0 6072 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_58
timestamp 1666464484
transform 1 0 6440 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1666464484
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1666464484
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1666464484
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_107
timestamp 1666464484
transform 1 0 10948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_120
timestamp 1666464484
transform 1 0 12144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1666464484
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_131
timestamp 1666464484
transform 1 0 13156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1666464484
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_12
timestamp 1666464484
transform 1 0 2208 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_63
timestamp 1666464484
transform 1 0 6900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1666464484
transform 1 0 8004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_88
timestamp 1666464484
transform 1 0 9200 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1666464484
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1666464484
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1666464484
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1666464484
transform 1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1666464484
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_38
timestamp 1666464484
transform 1 0 4600 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_47
timestamp 1666464484
transform 1 0 5428 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_59
timestamp 1666464484
transform 1 0 6532 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_67
timestamp 1666464484
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_91
timestamp 1666464484
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_98
timestamp 1666464484
transform 1 0 10120 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1666464484
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1666464484
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1666464484
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1666464484
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_17
timestamp 1666464484
transform 1 0 2668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1666464484
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_43
timestamp 1666464484
transform 1 0 5060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1666464484
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1666464484
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_77
timestamp 1666464484
transform 1 0 8188 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1666464484
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1666464484
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_48
timestamp 1666464484
transform 1 0 5520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1666464484
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_69
timestamp 1666464484
transform 1 0 7452 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_74
timestamp 1666464484
transform 1 0 7912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1666464484
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_45
timestamp 1666464484
transform 1 0 5244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 1666464484
transform 1 0 5612 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1666464484
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1666464484
transform 1 0 6716 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_65
timestamp 1666464484
transform 1 0 7084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_77
timestamp 1666464484
transform 1 0 8188 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_89
timestamp 1666464484
transform 1 0 9292 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_101
timestamp 1666464484
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1666464484
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1666464484
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1666464484
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1666464484
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_13
timestamp 1666464484
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_25
timestamp 1666464484
transform 1 0 3404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_37
timestamp 1666464484
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1666464484
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_29
timestamp 1666464484
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_41
timestamp 1666464484
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1666464484
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_85
timestamp 1666464484
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_97
timestamp 1666464484
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1666464484
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_141
timestamp 1666464484
transform 1 0 14076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_153
timestamp 1666464484
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1666464484
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_197
timestamp 1666464484
transform 1 0 19228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_209
timestamp 1666464484
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1666464484
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 22816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 22816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 22816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 22816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 22816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 22816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 22816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7452 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4416 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4324 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1666464484
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5152 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14352 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13524 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 1666464484
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_2  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12420 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _235_
timestamp 1666464484
transform 1 0 11868 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11684 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _238_
timestamp 1666464484
transform 1 0 11684 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5612 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12788 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13984 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1666464484
transform -1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _244_
timestamp 1666464484
transform -1 0 13800 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1666464484
transform -1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1666464484
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_4  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 17020 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_1  _249_
timestamp 1666464484
transform 1 0 16376 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15548 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _251_
timestamp 1666464484
transform -1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _252_
timestamp 1666464484
transform 1 0 17296 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _253_
timestamp 1666464484
transform -1 0 13524 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _254_
timestamp 1666464484
transform -1 0 13524 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _255_
timestamp 1666464484
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15364 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _257_
timestamp 1666464484
transform -1 0 15180 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _258_
timestamp 1666464484
transform 1 0 15456 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp 1666464484
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1666464484
transform -1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15456 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _265_
timestamp 1666464484
transform -1 0 17848 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1666464484
transform -1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1666464484
transform -1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _268_
timestamp 1666464484
transform -1 0 19872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _269_
timestamp 1666464484
transform -1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _270_
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _271_
timestamp 1666464484
transform 1 0 16008 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16652 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15732 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _274_
timestamp 1666464484
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1666464484
transform -1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1666464484
transform 1 0 14628 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _277_
timestamp 1666464484
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _278_
timestamp 1666464484
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _279_
timestamp 1666464484
transform 1 0 18400 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1666464484
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _281_
timestamp 1666464484
transform 1 0 19412 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19688 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18584 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _285_
timestamp 1666464484
transform 1 0 16836 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14628 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 1666464484
transform -1 0 17664 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _290_
timestamp 1666464484
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1666464484
transform -1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _292_
timestamp 1666464484
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 15088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13616 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _296_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12880 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _297_
timestamp 1666464484
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _298_
timestamp 1666464484
transform -1 0 18400 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _299_
timestamp 1666464484
transform 1 0 17572 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _300_
timestamp 1666464484
transform 1 0 18400 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _301_
timestamp 1666464484
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _302_
timestamp 1666464484
transform 1 0 17296 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1666464484
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _304_
timestamp 1666464484
transform -1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _305_
timestamp 1666464484
transform 1 0 16836 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _306_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19228 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _307_
timestamp 1666464484
transform -1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _308_
timestamp 1666464484
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18952 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _310_
timestamp 1666464484
transform 1 0 18400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _311_
timestamp 1666464484
transform 1 0 17388 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _312_
timestamp 1666464484
transform 1 0 19412 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _313_
timestamp 1666464484
transform -1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _314_
timestamp 1666464484
transform 1 0 19872 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _315_
timestamp 1666464484
transform 1 0 20608 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _316_
timestamp 1666464484
transform 1 0 20056 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _317_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19228 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _318_
timestamp 1666464484
transform 1 0 18216 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _319_
timestamp 1666464484
transform -1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _320_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _321_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 19228 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1666464484
transform 1 0 14076 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _323_
timestamp 1666464484
transform -1 0 15916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 13800 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _325_
timestamp 1666464484
transform 1 0 15824 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1666464484
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _327_
timestamp 1666464484
transform 1 0 15364 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _328_
timestamp 1666464484
transform 1 0 12696 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _329_
timestamp 1666464484
transform 1 0 12880 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _330_
timestamp 1666464484
transform -1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _331_
timestamp 1666464484
transform 1 0 14260 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _332_
timestamp 1666464484
transform 1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _333_
timestamp 1666464484
transform -1 0 2300 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _334_
timestamp 1666464484
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 1666464484
transform -1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14168 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _337_
timestamp 1666464484
transform -1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _339_
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _341_
timestamp 1666464484
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _342_
timestamp 1666464484
transform -1 0 14996 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 14996 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _344_
timestamp 1666464484
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp 1666464484
transform 1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _346_
timestamp 1666464484
transform 1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _347_
timestamp 1666464484
transform 1 0 11684 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1666464484
transform -1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _349_
timestamp 1666464484
transform 1 0 11776 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _350_
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _351_
timestamp 1666464484
transform -1 0 14996 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp 1666464484
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _353_
timestamp 1666464484
transform 1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _354_
timestamp 1666464484
transform 1 0 6532 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _355_
timestamp 1666464484
transform 1 0 11500 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _356_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _357_
timestamp 1666464484
transform -1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _358_
timestamp 1666464484
transform 1 0 3036 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _359_
timestamp 1666464484
transform 1 0 3956 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_4  _360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6716 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1666464484
transform 1 0 3956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _362_
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _363_
timestamp 1666464484
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _364_
timestamp 1666464484
transform -1 0 8556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _365_
timestamp 1666464484
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _366_
timestamp 1666464484
transform -1 0 8648 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _367_
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _368_
timestamp 1666464484
transform -1 0 10120 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _369_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7544 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _370_
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1666464484
transform -1 0 2668 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1666464484
transform 1 0 4968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _373_
timestamp 1666464484
transform -1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _374_
timestamp 1666464484
transform -1 0 8188 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _375_
timestamp 1666464484
transform -1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _376_
timestamp 1666464484
transform -1 0 5888 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _377_
timestamp 1666464484
transform 1 0 4692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1666464484
transform 1 0 1840 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1666464484
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _380_
timestamp 1666464484
transform -1 0 10120 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1666464484
transform 1 0 8924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _382_
timestamp 1666464484
transform 1 0 9108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _383_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1666464484
transform 1 0 3036 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1666464484
transform -1 0 3496 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _386_
timestamp 1666464484
transform -1 0 4232 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _387_
timestamp 1666464484
transform -1 0 6348 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _388_
timestamp 1666464484
transform 1 0 5704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _389_
timestamp 1666464484
transform -1 0 5520 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1666464484
transform 1 0 4232 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1666464484
transform 1 0 2760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _392_
timestamp 1666464484
transform -1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8648 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _394_
timestamp 1666464484
transform 1 0 6624 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _395_
timestamp 1666464484
transform -1 0 6900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1666464484
transform 1 0 6532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1666464484
transform 1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10028 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _400_
timestamp 1666464484
transform 1 0 6716 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _401_
timestamp 1666464484
transform -1 0 6440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _402_
timestamp 1666464484
transform -1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _403_
timestamp 1666464484
transform -1 0 7728 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _405_
timestamp 1666464484
transform -1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _406_
timestamp 1666464484
transform -1 0 3220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _407_
timestamp 1666464484
transform -1 0 4324 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _408_
timestamp 1666464484
transform -1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1666464484
transform 1 0 4784 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1666464484
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _411_
timestamp 1666464484
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _412_
timestamp 1666464484
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _413_
timestamp 1666464484
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _414_
timestamp 1666464484
transform -1 0 7636 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _415_
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _416_
timestamp 1666464484
transform -1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _417_
timestamp 1666464484
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _418_
timestamp 1666464484
transform 1 0 6072 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _419_
timestamp 1666464484
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _420_
timestamp 1666464484
transform 1 0 4784 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _421_
timestamp 1666464484
transform -1 0 3496 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _422_
timestamp 1666464484
transform 1 0 3956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _423_
timestamp 1666464484
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _424_
timestamp 1666464484
transform -1 0 5612 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _425_
timestamp 1666464484
transform -1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _426_
timestamp 1666464484
transform 1 0 3404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _427_
timestamp 1666464484
transform 1 0 2944 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _428_
timestamp 1666464484
transform 1 0 2668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _429_
timestamp 1666464484
transform -1 0 4784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _430_
timestamp 1666464484
transform -1 0 13800 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _431_
timestamp 1666464484
transform -1 0 10948 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _432_
timestamp 1666464484
transform 1 0 8372 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1666464484
transform -1 0 8464 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _434_
timestamp 1666464484
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp 1666464484
transform 1 0 6716 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _436_
timestamp 1666464484
transform -1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _437_
timestamp 1666464484
transform -1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _438_
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _439_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10028 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _440_
timestamp 1666464484
transform 1 0 9108 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9752 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _442_
timestamp 1666464484
transform 1 0 9752 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _443_
timestamp 1666464484
transform 1 0 7176 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _444_
timestamp 1666464484
transform -1 0 9292 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _445_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9292 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _446_
timestamp 1666464484
transform 1 0 6532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _447_
timestamp 1666464484
transform 1 0 10120 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _448_
timestamp 1666464484
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _449_
timestamp 1666464484
transform 1 0 9936 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp 1666464484
transform 1 0 9752 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1666464484
transform 1 0 10120 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _452_
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _453_
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1666464484
transform 1 0 9752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1666464484
transform 1 0 9936 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1666464484
transform -1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1666464484
transform 1 0 1564 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1666464484
transform -1 0 3036 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1666464484
transform 1 0 1564 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1666464484
transform 1 0 3956 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1666464484
transform 1 0 2208 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1666464484
transform 1 0 3956 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1666464484
transform 1 0 4324 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1666464484
transform 1 0 3404 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1666464484
transform 1 0 1564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1666464484
transform -1 0 9292 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1666464484
transform 1 0 6992 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1666464484
transform 1 0 4600 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1666464484
transform 1 0 4140 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1666464484
transform 1 0 2392 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1666464484
transform 1 0 1564 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1666464484
transform 1 0 1564 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _475_
timestamp 1666464484
transform 1 0 4600 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _476_
timestamp 1666464484
transform 1 0 7176 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _477_
timestamp 1666464484
transform 1 0 6164 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _478_
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _479_
timestamp 1666464484
transform -1 0 8924 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _480_
timestamp 1666464484
transform 1 0 5152 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5888 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1666464484
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1666464484
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1666464484
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1666464484
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 19668 800 19908 0 FreeSans 960 0 0 0 OP
port 0 nsew signal tristate
flabel metal3 s 0 3892 800 4132 0 FreeSans 960 0 0 0 clk
port 1 nsew signal input
flabel metal3 s 0 11780 800 12020 0 FreeSans 960 0 0 0 rst
port 2 nsew signal input
flabel metal4 s 3658 2128 3978 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 9086 2128 9406 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 14514 2128 14834 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 19942 2128 20262 21808 0 FreeSans 1920 90 0 0 vccd1
port 3 nsew power bidirectional
flabel metal4 s 6372 2128 6692 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 11800 2128 12120 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 17228 2128 17548 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
flabel metal4 s 22656 2128 22976 21808 0 FreeSans 1920 90 0 0 vssd1
port 4 nsew ground bidirectional
rlabel metal1 11960 21216 11960 21216 0 vccd1
rlabel via1 12040 21760 12040 21760 0 vssd1
rlabel metal2 2714 10642 2714 10642 0 LFSR\[0\]
rlabel metal2 2530 14144 2530 14144 0 LFSR\[1\]
rlabel viali 5211 14314 5211 14314 0 LFSR\[2\]
rlabel metal1 3910 13906 3910 13906 0 LFSR\[3\]
rlabel metal1 5428 12818 5428 12818 0 LFSR\[4\]
rlabel metal2 6900 12954 6900 12954 0 LFSR\[5\]
rlabel metal1 5060 11526 5060 11526 0 LFSR\[6\]
rlabel metal2 2162 19635 2162 19635 0 OP
rlabel metal1 2070 11050 2070 11050 0 OP_reg
rlabel via1 12650 12971 12650 12971 0 PC\[0\]
rlabel metal1 14122 7310 14122 7310 0 PC\[1\]
rlabel metal1 15916 2346 15916 2346 0 PC\[2\]
rlabel metal1 14582 4624 14582 4624 0 PC\[3\]
rlabel metal1 13386 7888 13386 7888 0 PC\[4\]
rlabel metal2 11178 3230 11178 3230 0 PC\[5\]
rlabel metal1 14651 8602 14651 8602 0 _000_
rlabel metal2 11270 6970 11270 6970 0 _001_
rlabel metal2 17434 7463 17434 7463 0 _002_
rlabel metal2 18630 5576 18630 5576 0 _003_
rlabel metal1 12742 6392 12742 6392 0 _004_
rlabel metal1 9430 5780 9430 5780 0 _005_
rlabel metal1 12581 8806 12581 8806 0 _006_
rlabel metal2 12558 10234 12558 10234 0 _007_
rlabel metal1 11035 11118 11035 11118 0 _008_
rlabel metal1 10989 10710 10989 10710 0 _009_
rlabel metal1 17158 5746 17158 5746 0 _010_
rlabel metal2 16422 6052 16422 6052 0 _011_
rlabel metal1 16606 4522 16606 4522 0 _012_
rlabel metal1 14398 5678 14398 5678 0 _013_
rlabel metal2 18906 7344 18906 7344 0 _014_
rlabel metal1 12834 6698 12834 6698 0 _015_
rlabel metal1 9384 12614 9384 12614 0 _016_
rlabel via1 1881 10642 1881 10642 0 _017_
rlabel metal2 4462 10472 4462 10472 0 _018_
rlabel metal1 1927 9622 1927 9622 0 _019_
rlabel metal2 4232 10676 4232 10676 0 _020_
rlabel metal1 2376 8534 2376 8534 0 _021_
rlabel metal1 4319 9622 4319 9622 0 _022_
rlabel metal1 5193 10030 5193 10030 0 _023_
rlabel metal1 3618 10710 3618 10710 0 _024_
rlabel metal2 1978 7650 1978 7650 0 _025_
rlabel metal1 6435 4522 6435 4522 0 _026_
rlabel metal1 9062 2618 9062 2618 0 _027_
rlabel metal1 7212 3502 7212 3502 0 _028_
rlabel metal2 6118 3910 6118 3910 0 _029_
rlabel metal2 4830 3298 4830 3298 0 _030_
rlabel metal1 2893 4114 2893 4114 0 _031_
rlabel metal1 2663 5202 2663 5202 0 _032_
rlabel metal2 2714 6086 2714 6086 0 _033_
rlabel metal1 4814 6358 4814 6358 0 _034_
rlabel metal1 7953 8942 7953 8942 0 _035_
rlabel metal1 6240 9962 6240 9962 0 _036_
rlabel metal1 6987 10710 6987 10710 0 _037_
rlabel metal1 8704 8466 8704 8466 0 _038_
rlabel metal1 12144 2618 12144 2618 0 _039_
rlabel metal1 18676 4998 18676 4998 0 _040_
rlabel metal1 19642 3672 19642 3672 0 _041_
rlabel metal1 14444 4182 14444 4182 0 _042_
rlabel metal1 14214 6766 14214 6766 0 _043_
rlabel metal2 15042 6154 15042 6154 0 _044_
rlabel metal2 12466 13056 12466 13056 0 _045_
rlabel metal1 12558 12784 12558 12784 0 _046_
rlabel metal1 16767 12886 16767 12886 0 _047_
rlabel metal2 15778 4046 15778 4046 0 _048_
rlabel metal1 17020 3570 17020 3570 0 _049_
rlabel metal1 16146 3434 16146 3434 0 _050_
rlabel metal1 17572 3434 17572 3434 0 _051_
rlabel metal1 13570 3570 13570 3570 0 _052_
rlabel metal1 13156 2414 13156 2414 0 _053_
rlabel metal1 18630 2414 18630 2414 0 _054_
rlabel metal1 14766 4624 14766 4624 0 _055_
rlabel metal1 14444 2890 14444 2890 0 _056_
rlabel metal2 15870 4216 15870 4216 0 _057_
rlabel metal1 17158 2414 17158 2414 0 _058_
rlabel metal1 17434 2618 17434 2618 0 _059_
rlabel metal2 16054 5984 16054 5984 0 _060_
rlabel metal1 17204 4114 17204 4114 0 _061_
rlabel metal1 17250 2278 17250 2278 0 _062_
rlabel metal2 18722 7106 18722 7106 0 _063_
rlabel metal2 15226 7174 15226 7174 0 _064_
rlabel via1 17810 7786 17810 7786 0 _065_
rlabel metal1 15962 7344 15962 7344 0 _066_
rlabel metal1 16744 7514 16744 7514 0 _067_
rlabel metal1 16376 9078 16376 9078 0 _068_
rlabel metal1 16652 8466 16652 8466 0 _069_
rlabel metal1 20332 5678 20332 5678 0 _070_
rlabel metal2 14030 7956 14030 7956 0 _071_
rlabel metal2 15686 8160 15686 8160 0 _072_
rlabel metal1 18814 8500 18814 8500 0 _073_
rlabel metal1 17250 6256 17250 6256 0 _074_
rlabel metal2 18998 8670 18998 8670 0 _075_
rlabel metal1 19136 2278 19136 2278 0 _076_
rlabel metal1 19734 8058 19734 8058 0 _077_
rlabel metal1 19274 8432 19274 8432 0 _078_
rlabel metal1 17986 8398 17986 8398 0 _079_
rlabel metal1 13386 7310 13386 7310 0 _080_
rlabel metal2 13294 7548 13294 7548 0 _081_
rlabel metal1 16100 7922 16100 7922 0 _082_
rlabel metal2 15226 8194 15226 8194 0 _083_
rlabel metal1 14536 5746 14536 5746 0 _084_
rlabel metal2 18538 3604 18538 3604 0 _085_
rlabel metal1 18584 4794 18584 4794 0 _086_
rlabel metal1 14858 3706 14858 3706 0 _087_
rlabel metal1 14214 5882 14214 5882 0 _088_
rlabel metal2 13386 7820 13386 7820 0 _089_
rlabel metal2 18078 8772 18078 8772 0 _090_
rlabel metal2 18630 8228 18630 8228 0 _091_
rlabel metal1 18906 7412 18906 7412 0 _092_
rlabel metal1 18078 7378 18078 7378 0 _093_
rlabel metal1 17112 5882 17112 5882 0 _094_
rlabel metal1 18354 4250 18354 4250 0 _095_
rlabel metal1 19550 4046 19550 4046 0 _096_
rlabel metal2 17986 5576 17986 5576 0 _097_
rlabel metal1 17572 6426 17572 6426 0 _098_
rlabel metal2 20562 3706 20562 3706 0 _099_
rlabel metal1 19182 2618 19182 2618 0 _100_
rlabel metal1 18814 2992 18814 2992 0 _101_
rlabel metal2 18906 3196 18906 3196 0 _102_
rlabel metal1 18354 3162 18354 3162 0 _103_
rlabel metal1 19412 5202 19412 5202 0 _104_
rlabel metal2 19550 5372 19550 5372 0 _105_
rlabel metal2 20378 6698 20378 6698 0 _106_
rlabel metal1 20286 5270 20286 5270 0 _107_
rlabel metal2 19826 5712 19826 5712 0 _108_
rlabel metal2 19274 5780 19274 5780 0 _109_
rlabel metal1 18906 5338 18906 5338 0 _110_
rlabel metal1 19734 5882 19734 5882 0 _111_
rlabel metal2 19458 6086 19458 6086 0 _112_
rlabel metal1 14076 5338 14076 5338 0 _113_
rlabel metal2 14030 6494 14030 6494 0 _114_
rlabel metal1 13432 6290 13432 6290 0 _115_
rlabel metal2 13294 5984 13294 5984 0 _116_
rlabel metal1 13294 6222 13294 6222 0 _117_
rlabel metal1 14352 6358 14352 6358 0 _118_
rlabel metal1 12834 5338 12834 5338 0 _119_
rlabel metal1 12926 5576 12926 5576 0 _120_
rlabel metal1 14260 4794 14260 4794 0 _121_
rlabel metal1 1932 19346 1932 19346 0 _122_
rlabel metal1 14674 10064 14674 10064 0 _123_
rlabel metal1 13846 9554 13846 9554 0 _124_
rlabel metal1 10948 12818 10948 12818 0 _125_
rlabel metal1 13570 12750 13570 12750 0 _126_
rlabel metal2 12926 9146 12926 9146 0 _127_
rlabel metal1 14352 11322 14352 11322 0 _128_
rlabel metal1 14674 11866 14674 11866 0 _129_
rlabel metal1 14306 10710 14306 10710 0 _130_
rlabel metal1 12972 10642 12972 10642 0 _131_
rlabel metal1 10718 13396 10718 13396 0 _132_
rlabel metal1 11500 11866 11500 11866 0 _133_
rlabel metal1 12006 11220 12006 11220 0 _134_
rlabel metal2 14306 9554 14306 9554 0 _135_
rlabel metal1 14122 9894 14122 9894 0 _136_
rlabel metal2 12098 10438 12098 10438 0 _137_
rlabel metal1 4048 2346 4048 2346 0 _138_
rlabel metal1 10350 12750 10350 12750 0 _139_
rlabel metal1 9476 12818 9476 12818 0 _140_
rlabel metal1 3772 12410 3772 12410 0 _141_
rlabel metal1 5106 12070 5106 12070 0 _142_
rlabel metal1 2208 11594 2208 11594 0 _143_
rlabel metal1 2254 11764 2254 11764 0 _144_
rlabel metal1 1794 11152 1794 11152 0 _145_
rlabel metal2 5198 15742 5198 15742 0 _146_
rlabel metal1 8372 15674 8372 15674 0 _147_
rlabel metal1 7866 15436 7866 15436 0 _148_
rlabel metal2 7774 14994 7774 14994 0 _149_
rlabel metal2 7590 14926 7590 14926 0 _150_
rlabel metal1 5198 13294 5198 13294 0 _151_
rlabel metal2 2162 12716 2162 12716 0 _152_
rlabel metal2 2622 11628 2622 11628 0 _153_
rlabel metal2 7038 15674 7038 15674 0 _154_
rlabel metal1 7360 15130 7360 15130 0 _155_
rlabel metal1 5014 14416 5014 14416 0 _156_
rlabel metal2 4922 14586 4922 14586 0 _157_
rlabel metal2 2346 14756 2346 14756 0 _158_
rlabel metal2 2162 14348 2162 14348 0 _159_
rlabel metal1 9338 14994 9338 14994 0 _160_
rlabel metal1 8970 13838 8970 13838 0 _161_
rlabel metal1 9430 14586 9430 14586 0 _162_
rlabel via2 3542 14909 3542 14909 0 _163_
rlabel metal2 2990 14620 2990 14620 0 _164_
rlabel metal1 3726 14382 3726 14382 0 _165_
rlabel metal2 5290 15742 5290 15742 0 _166_
rlabel metal1 5520 15470 5520 15470 0 _167_
rlabel metal1 4830 15130 4830 15130 0 _168_
rlabel metal2 3266 14416 3266 14416 0 _169_
rlabel metal2 2070 14212 2070 14212 0 _170_
rlabel metal2 6762 13294 6762 13294 0 _171_
rlabel metal1 6670 13838 6670 13838 0 _172_
rlabel metal1 7084 12954 7084 12954 0 _173_
rlabel metal1 5888 12954 5888 12954 0 _174_
rlabel metal1 4646 12614 4646 12614 0 _175_
rlabel metal1 7222 15028 7222 15028 0 _176_
rlabel metal1 6624 13294 6624 13294 0 _177_
rlabel metal1 6900 13158 6900 13158 0 _178_
rlabel metal1 6670 11866 6670 11866 0 _179_
rlabel metal2 4094 14348 4094 14348 0 _180_
rlabel metal1 2944 11322 2944 11322 0 _181_
rlabel metal1 3726 12750 3726 12750 0 _182_
rlabel metal2 4278 12240 4278 12240 0 _183_
rlabel metal1 2461 7378 2461 7378 0 _184_
rlabel metal1 9338 2448 9338 2448 0 _185_
rlabel metal1 7268 2618 7268 2618 0 _186_
rlabel metal1 7728 4114 7728 4114 0 _187_
rlabel metal1 6026 2618 6026 2618 0 _188_
rlabel metal1 5060 2618 5060 2618 0 _189_
rlabel metal1 3128 3706 3128 3706 0 _190_
rlabel metal1 3634 4726 3634 4726 0 _191_
rlabel metal1 3174 5644 3174 5644 0 _192_
rlabel metal1 3588 5202 3588 5202 0 _193_
rlabel metal2 2898 6154 2898 6154 0 _194_
rlabel metal1 11546 12614 11546 12614 0 _195_
rlabel metal1 9706 13430 9706 13430 0 _196_
rlabel metal1 7314 11220 7314 11220 0 _197_
rlabel metal2 6486 11492 6486 11492 0 _198_
rlabel metal2 5842 11322 5842 11322 0 _199_
rlabel metal2 7774 11628 7774 11628 0 _200_
rlabel metal2 9430 11934 9430 11934 0 _201_
rlabel metal1 4876 6766 4876 6766 0 _202_
rlabel metal1 6394 3026 6394 3026 0 _203_
rlabel metal1 5474 2414 5474 2414 0 _204_
rlabel metal1 3680 2618 3680 2618 0 _205_
rlabel metal1 4738 6732 4738 6732 0 _206_
rlabel metal1 4600 6766 4600 6766 0 _207_
rlabel metal2 4462 7548 4462 7548 0 _208_
rlabel metal2 12374 13056 12374 13056 0 _209_
rlabel metal1 14352 12818 14352 12818 0 _210_
rlabel metal1 14582 10778 14582 10778 0 _211_
rlabel metal2 14214 13056 14214 13056 0 _212_
rlabel metal1 14352 12614 14352 12614 0 _213_
rlabel metal1 10994 11764 10994 11764 0 _214_
rlabel metal1 12834 12206 12834 12206 0 _215_
rlabel metal1 15594 2414 15594 2414 0 _216_
rlabel metal1 13432 3706 13432 3706 0 _217_
rlabel metal1 11546 2346 11546 2346 0 _218_
rlabel metal2 11730 2618 11730 2618 0 _219_
rlabel metal2 5934 5304 5934 5304 0 clk
rlabel metal1 6118 3094 6118 3094 0 clknet_0_clk
rlabel metal2 2714 3332 2714 3332 0 clknet_2_0__leaf_clk
rlabel metal1 1932 8398 1932 8398 0 clknet_2_1__leaf_clk
rlabel metal2 6026 5168 6026 5168 0 clknet_2_2__leaf_clk
rlabel metal2 6210 10336 6210 10336 0 clknet_2_3__leaf_clk
rlabel metal1 7406 2346 7406 2346 0 clock_div\[0\]
rlabel metal1 7260 2278 7260 2278 0 clock_div\[1\]
rlabel metal1 8096 2414 8096 2414 0 clock_div\[2\]
rlabel metal2 6578 3740 6578 3740 0 clock_div\[3\]
rlabel metal1 4876 2482 4876 2482 0 clock_div\[4\]
rlabel metal1 3864 2414 3864 2414 0 clock_div\[5\]
rlabel metal1 3910 5100 3910 5100 0 clock_div\[6\]
rlabel metal1 3358 6800 3358 6800 0 clock_div\[7\]
rlabel metal1 5612 6426 5612 6426 0 clock_div\[8\]
rlabel metal1 2070 12852 2070 12852 0 just_inc
rlabel metal1 13018 13294 13018 13294 0 just_rst
rlabel metal1 17296 2346 17296 2346 0 net1
rlabel metal2 4094 7990 4094 7990 0 prev_clk_div
rlabel metal2 13386 10098 13386 10098 0 rhythm_LFSR\[0\]
rlabel metal1 13708 10778 13708 10778 0 rhythm_LFSR\[1\]
rlabel metal2 13938 11832 13938 11832 0 rhythm_LFSR\[2\]
rlabel metal1 13570 11696 13570 11696 0 rhythm_LFSR\[3\]
rlabel metal1 3082 13158 3082 13158 0 rst
rlabel metal2 8970 9894 8970 9894 0 tempo_LFSR\[0\]
rlabel metal1 9292 11526 9292 11526 0 tempo_LFSR\[1\]
rlabel metal2 8418 10948 8418 10948 0 tempo_LFSR\[2\]
rlabel metal1 7590 11050 7590 11050 0 tempo_LFSR\[3\]
rlabel metal1 14490 11084 14490 11084 0 tune_ROM\[0\]
rlabel metal2 15226 10591 15226 10591 0 tune_ROM\[1\]
rlabel metal1 10074 14450 10074 14450 0 tune_ROM\[2\]
rlabel metal1 8648 14382 8648 14382 0 tune_ROM\[3\]
rlabel metal1 6394 16082 6394 16082 0 tune_ROM\[4\]
rlabel metal1 9108 13158 9108 13158 0 tune_ROM\[5\]
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
