magic
tech sky130B
magscale 1 2
timestamp 1674824011
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 14 1980 29334 27792
<< metal2 >>
rect 1306 29200 1362 30000
rect 3790 29200 3846 30000
rect 6274 29200 6330 30000
rect 8758 29200 8814 30000
rect 11242 29200 11298 30000
rect 13726 29200 13782 30000
rect 16210 29200 16266 30000
rect 18694 29200 18750 30000
rect 21178 29200 21234 30000
rect 23662 29200 23718 30000
rect 26146 29200 26202 30000
rect 28630 29200 28686 30000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3882 0 3938 800
rect 4986 0 5042 800
rect 6090 0 6146 800
rect 7194 0 7250 800
rect 8298 0 8354 800
rect 9402 0 9458 800
rect 10506 0 10562 800
rect 11610 0 11666 800
rect 12714 0 12770 800
rect 13818 0 13874 800
rect 14922 0 14978 800
rect 16026 0 16082 800
rect 17130 0 17186 800
rect 18234 0 18290 800
rect 19338 0 19394 800
rect 20442 0 20498 800
rect 21546 0 21602 800
rect 22650 0 22706 800
rect 23754 0 23810 800
rect 24858 0 24914 800
rect 25962 0 26018 800
rect 27066 0 27122 800
rect 28170 0 28226 800
rect 29274 0 29330 800
<< obsm2 >>
rect 20 29144 1250 29322
rect 1418 29144 3734 29322
rect 3902 29144 6218 29322
rect 6386 29144 8702 29322
rect 8870 29144 11186 29322
rect 11354 29144 13670 29322
rect 13838 29144 16154 29322
rect 16322 29144 18638 29322
rect 18806 29144 21122 29322
rect 21290 29144 23606 29322
rect 23774 29144 26090 29322
rect 26258 29144 28574 29322
rect 28742 29144 29328 29322
rect 20 856 29328 29144
rect 20 734 514 856
rect 682 734 1618 856
rect 1786 734 2722 856
rect 2890 734 3826 856
rect 3994 734 4930 856
rect 5098 734 6034 856
rect 6202 734 7138 856
rect 7306 734 8242 856
rect 8410 734 9346 856
rect 9514 734 10450 856
rect 10618 734 11554 856
rect 11722 734 12658 856
rect 12826 734 13762 856
rect 13930 734 14866 856
rect 15034 734 15970 856
rect 16138 734 17074 856
rect 17242 734 18178 856
rect 18346 734 19282 856
rect 19450 734 20386 856
rect 20554 734 21490 856
rect 21658 734 22594 856
rect 22762 734 23698 856
rect 23866 734 24802 856
rect 24970 734 25906 856
rect 26074 734 27010 856
rect 27178 734 28114 856
rect 28282 734 29218 856
<< metal3 >>
rect 29200 14832 30000 14952
<< obsm3 >>
rect 1853 15032 29200 27777
rect 1853 14752 29120 15032
rect 1853 2143 29200 14752
<< metal4 >>
rect 4417 2128 4737 27792
rect 7890 2128 8210 27792
rect 11363 2128 11683 27792
rect 14836 2128 15156 27792
rect 18309 2128 18629 27792
rect 21782 2128 22102 27792
rect 25255 2128 25575 27792
rect 28728 2128 29048 27792
<< obsm4 >>
rect 4107 3707 4337 26349
rect 4817 3707 7810 26349
rect 8290 3707 11283 26349
rect 11763 3707 14756 26349
rect 15236 3707 18229 26349
rect 18709 3707 19629 26349
<< labels >>
rlabel metal2 s 1306 29200 1362 30000 6 clk
port 1 nsew signal input
rlabel metal2 s 6274 29200 6330 30000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 8758 29200 8814 30000 6 io_in[1]
port 3 nsew signal input
rlabel metal2 s 11242 29200 11298 30000 6 io_in[2]
port 4 nsew signal input
rlabel metal2 s 13726 29200 13782 30000 6 io_in[3]
port 5 nsew signal input
rlabel metal2 s 16210 29200 16266 30000 6 io_in[4]
port 6 nsew signal input
rlabel metal2 s 18694 29200 18750 30000 6 io_in[5]
port 7 nsew signal input
rlabel metal2 s 21178 29200 21234 30000 6 io_in[6]
port 8 nsew signal input
rlabel metal2 s 23662 29200 23718 30000 6 io_in[7]
port 9 nsew signal input
rlabel metal2 s 26146 29200 26202 30000 6 io_in[8]
port 10 nsew signal input
rlabel metal2 s 28630 29200 28686 30000 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 29200 14832 30000 14952 6 io_oeb
port 12 nsew signal output
rlabel metal2 s 570 0 626 800 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 23754 0 23810 800 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 io_out[2]
port 32 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 io_out[3]
port 33 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 io_out[4]
port 34 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 io_out[5]
port 35 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 io_out[6]
port 36 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 io_out[7]
port 37 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 io_out[8]
port 38 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 io_out[9]
port 39 nsew signal output
rlabel metal2 s 3790 29200 3846 30000 6 rst
port 40 nsew signal input
rlabel metal4 s 4417 2128 4737 27792 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 7890 2128 8210 27792 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 14836 2128 15156 27792 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 21782 2128 22102 27792 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 28728 2128 29048 27792 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2885152
string GDS_FILE /media/lucah/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS5401/runs/23_01_27_13_50/results/signoff/tholin_avalonsemi_5401.magic.gds
string GDS_START 584214
<< end >>

