// This is the unpowered netlist.
module multiplexer (design_clk_o,
    dso_tune,
    oeb_6502,
    oeb_as1802,
    oeb_as2650,
    oeb_as5401,
    oeb_mc14500,
    rst_6502,
    rst_LCD,
    rst_as1802,
    rst_as2650,
    rst_as5401,
    rst_counter,
    rst_diceroll,
    rst_mc14500,
    rst_tbb1143,
    rst_tune,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    dsi_all,
    dso_6502,
    dso_LCD,
    dso_as1802,
    dso_as2650,
    dso_as5401,
    dso_counter,
    dso_diceroll,
    dso_mc14500,
    dso_multiplier,
    dso_tbb1143,
    io_in,
    io_oeb,
    io_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output design_clk_o;
 input dso_tune;
 input oeb_6502;
 input oeb_as1802;
 input oeb_as2650;
 input oeb_as5401;
 input oeb_mc14500;
 output rst_6502;
 output rst_LCD;
 output rst_as1802;
 output rst_as2650;
 output rst_as5401;
 output rst_counter;
 output rst_diceroll;
 output rst_mc14500;
 output rst_tbb1143;
 output rst_tune;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [26:0] dsi_all;
 input [26:0] dso_6502;
 input [7:0] dso_LCD;
 input [26:0] dso_as1802;
 input [26:0] dso_as2650;
 input [26:0] dso_as5401;
 input [11:0] dso_counter;
 input [7:0] dso_diceroll;
 input [8:0] dso_mc14500;
 input [7:0] dso_multiplier;
 input [7:0] dso_tbb1143;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire \design_addr[0] ;
 wire \design_addr[1] ;
 wire \design_addr[2] ;
 wire \design_addr[3] ;
 wire net374;
 wire clknet_0_wb_clk_i;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net358;
 wire net368;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire wb_clk_override;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[2] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire \wb_design_addr_override[0] ;
 wire \wb_design_addr_override[1] ;
 wire \wb_design_addr_override[2] ;
 wire \wb_design_addr_override[3] ;
 wire wb_feedback_delay;
 wire \wb_io_override[0] ;
 wire \wb_io_override[10] ;
 wire \wb_io_override[11] ;
 wire \wb_io_override[12] ;
 wire \wb_io_override[13] ;
 wire \wb_io_override[14] ;
 wire \wb_io_override[15] ;
 wire \wb_io_override[16] ;
 wire \wb_io_override[17] ;
 wire \wb_io_override[18] ;
 wire \wb_io_override[19] ;
 wire \wb_io_override[1] ;
 wire \wb_io_override[20] ;
 wire \wb_io_override[21] ;
 wire \wb_io_override[22] ;
 wire \wb_io_override[23] ;
 wire \wb_io_override[24] ;
 wire \wb_io_override[25] ;
 wire \wb_io_override[26] ;
 wire \wb_io_override[2] ;
 wire \wb_io_override[3] ;
 wire \wb_io_override[4] ;
 wire \wb_io_override[5] ;
 wire \wb_io_override[6] ;
 wire \wb_io_override[7] ;
 wire \wb_io_override[8] ;
 wire \wb_io_override[9] ;
 wire wb_override;
 wire wb_rst_override;
 wire wb_single_step;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_0_net235;
 wire clknet_1_0__leaf_net235;
 wire clknet_1_1__leaf_net235;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;

 sky130_fd_sc_hd__mux2_4 _0574_ (.A0(net195),
    .A1(wb_rst_override),
    .S(wb_override),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_4 _0575_ (.A(\design_addr[1] ),
    .X(_0222_));
 sky130_fd_sc_hd__clkinv_2 _0576_ (.A(\design_addr[0] ),
    .Y(_0223_));
 sky130_fd_sc_hd__or2_1 _0577_ (.A(\design_addr[3] ),
    .B(\design_addr[2] ),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_4 _0578_ (.A(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__nor3_4 _0579_ (.A(_0222_),
    .B(_0223_),
    .C(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__clkbuf_4 _0580_ (.A(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_4 _0581_ (.A(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__or2b_1 _0582_ (.A(_0221_),
    .B_N(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _0583_ (.A(_0229_),
    .X(net321));
 sky130_fd_sc_hd__buf_2 _0584_ (.A(\design_addr[0] ),
    .X(_0230_));
 sky130_fd_sc_hd__nor3b_1 _0585_ (.A(_0230_),
    .B(_0225_),
    .C_N(\design_addr[1] ),
    .Y(_0231_));
 sky130_fd_sc_hd__clkbuf_4 _0586_ (.A(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__or2b_1 _0587_ (.A(_0221_),
    .B_N(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_1 _0588_ (.A(_0233_),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 _0589_ (.A(\design_addr[3] ),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_2 _0590_ (.A(\design_addr[2] ),
    .X(_0235_));
 sky130_fd_sc_hd__and4bb_1 _0591_ (.A_N(_0234_),
    .B_N(_0235_),
    .C(_0222_),
    .D(_0230_),
    .X(_0236_));
 sky130_fd_sc_hd__clkbuf_4 _0592_ (.A(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__or2b_1 _0593_ (.A(_0221_),
    .B_N(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _0594_ (.A(_0238_),
    .X(net318));
 sky130_fd_sc_hd__or2b_1 _0595_ (.A(_0234_),
    .B_N(_0235_),
    .X(_0239_));
 sky130_fd_sc_hd__or4_1 _0596_ (.A(_0222_),
    .B(_0230_),
    .C(_0221_),
    .D(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0240_),
    .X(net324));
 sky130_fd_sc_hd__and4bb_2 _0598_ (.A_N(_0222_),
    .B_N(_0234_),
    .C(_0235_),
    .D(_0230_),
    .X(_0241_));
 sky130_fd_sc_hd__clkbuf_4 _0599_ (.A(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__or2b_1 _0600_ (.A(_0221_),
    .B_N(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_1 _0601_ (.A(_0243_),
    .X(net322));
 sky130_fd_sc_hd__and4bb_1 _0602_ (.A_N(\design_addr[0] ),
    .B_N(_0234_),
    .C(_0235_),
    .D(\design_addr[1] ),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_4 _0603_ (.A(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__or2b_1 _0604_ (.A(_0221_),
    .B_N(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_1 _0605_ (.A(_0246_),
    .X(net325));
 sky130_fd_sc_hd__and4b_1 _0606_ (.A_N(_0234_),
    .B(_0235_),
    .C(\design_addr[1] ),
    .D(\design_addr[0] ),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_4 _0607_ (.A(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__clkbuf_4 _0608_ (.A(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_4 _0609_ (.A(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__or2b_1 _0610_ (.A(_0221_),
    .B_N(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_1 _0611_ (.A(_0251_),
    .X(net320));
 sky130_fd_sc_hd__or3b_2 _0612_ (.A(_0222_),
    .B(_0235_),
    .C_N(_0234_),
    .X(_0252_));
 sky130_fd_sc_hd__or3_1 _0613_ (.A(_0230_),
    .B(_0221_),
    .C(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0614_ (.A(_0253_),
    .X(net317));
 sky130_fd_sc_hd__or3_1 _0615_ (.A(_0223_),
    .B(_0221_),
    .C(_0252_),
    .X(_0254_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0254_),
    .X(net319));
 sky130_fd_sc_hd__and4bb_1 _0617_ (.A_N(\design_addr[0] ),
    .B_N(_0235_),
    .C(_0234_),
    .D(\design_addr[1] ),
    .X(_0255_));
 sky130_fd_sc_hd__or2b_1 _0618_ (.A(_0221_),
    .B_N(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_1 _0619_ (.A(_0256_),
    .X(net326));
 sky130_fd_sc_hd__nor4b_4 _0620_ (.A(\design_addr[1] ),
    .B(\design_addr[0] ),
    .C(\design_addr[2] ),
    .D_N(\design_addr[3] ),
    .Y(_0257_));
 sky130_fd_sc_hd__and4bb_2 _0621_ (.A_N(\design_addr[1] ),
    .B_N(_0235_),
    .C(_0234_),
    .D(\design_addr[0] ),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_2 _0622_ (.A1(net196),
    .A2(_0257_),
    .B1(_0258_),
    .B2(net197),
    .X(_0259_));
 sky130_fd_sc_hd__a211o_1 _0623_ (.A1(net198),
    .A2(_0249_),
    .B1(net199),
    .C1(_0223_),
    .X(_0260_));
 sky130_fd_sc_hd__nor2_1 _0624_ (.A(_0222_),
    .B(_0225_),
    .Y(_0261_));
 sky130_fd_sc_hd__a211o_1 _0625_ (.A1(net198),
    .A2(_0247_),
    .B1(_0259_),
    .C1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__buf_4 _0626_ (.A(_0262_),
    .X(net270));
 sky130_fd_sc_hd__nor2_1 _0627_ (.A(_0230_),
    .B(_0239_),
    .Y(_0263_));
 sky130_fd_sc_hd__o22ai_4 _0628_ (.A1(_0259_),
    .A2(_0260_),
    .B1(net270),
    .B2(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__clkinv_2 _0629_ (.A(_0264_),
    .Y(net266));
 sky130_fd_sc_hd__or2_1 _0630_ (.A(_0232_),
    .B(net266),
    .X(_0265_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0631_ (.A(_0265_),
    .X(net263));
 sky130_fd_sc_hd__nor3_1 _0632_ (.A(_0222_),
    .B(_0230_),
    .C(_0239_),
    .Y(_0266_));
 sky130_fd_sc_hd__clkbuf_4 _0633_ (.A(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__or2_1 _0634_ (.A(_0245_),
    .B(net270),
    .X(_0268_));
 sky130_fd_sc_hd__buf_2 _0635_ (.A(_0268_),
    .X(net268));
 sky130_fd_sc_hd__a21o_1 _0636_ (.A1(net200),
    .A2(_0267_),
    .B1(net268),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_2 _0637_ (.A(_0269_),
    .X(net267));
 sky130_fd_sc_hd__o21ai_4 _0638_ (.A1(_0223_),
    .A2(_0225_),
    .B1(_0252_),
    .Y(net272));
 sky130_fd_sc_hd__clkbuf_4 _0639_ (.A(_0258_),
    .X(_0270_));
 sky130_fd_sc_hd__buf_2 _0640_ (.A(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__clkbuf_4 _0641_ (.A(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_1 _0642_ (.A(_0237_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _0643_ (.A(_0273_),
    .Y(net274));
 sky130_fd_sc_hd__nor2_1 _0644_ (.A(_0242_),
    .B(net274),
    .Y(_0274_));
 sky130_fd_sc_hd__clkinv_2 _0645_ (.A(_0274_),
    .Y(net275));
 sky130_fd_sc_hd__or3_1 _0646_ (.A(_0237_),
    .B(_0267_),
    .C(_0241_),
    .X(_0275_));
 sky130_fd_sc_hd__buf_2 _0647_ (.A(_0275_),
    .X(net276));
 sky130_fd_sc_hd__or2_1 _0648_ (.A(_0245_),
    .B(net276),
    .X(_0276_));
 sky130_fd_sc_hd__buf_2 _0649_ (.A(_0276_),
    .X(net278));
 sky130_fd_sc_hd__nor3_4 _0650_ (.A(_0222_),
    .B(_0230_),
    .C(_0225_),
    .Y(_0277_));
 sky130_fd_sc_hd__or2_1 _0651_ (.A(net278),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_2 _0652_ (.A(_0278_),
    .X(net289));
 sky130_fd_sc_hd__and2_1 _0653_ (.A(net162),
    .B(_0255_),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_2 _0654_ (.A(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__a221o_1 _0655_ (.A1(net117),
    .A2(_0242_),
    .B1(_0250_),
    .B2(net63),
    .C1(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__buf_2 _0656_ (.A(_0257_),
    .X(_0282_));
 sky130_fd_sc_hd__a22o_1 _0657_ (.A1(net28),
    .A2(_0237_),
    .B1(_0282_),
    .B2(net1),
    .X(_0283_));
 sky130_fd_sc_hd__a221o_1 _0658_ (.A1(net90),
    .A2(_0228_),
    .B1(_0272_),
    .B2(net36),
    .C1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _0659_ (.A(_0281_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_2 _0660_ (.A(_0285_),
    .X(net290));
 sky130_fd_sc_hd__a22o_1 _0661_ (.A1(net101),
    .A2(_0228_),
    .B1(_0272_),
    .B2(net47),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _0662_ (.A(_0257_),
    .X(_0287_));
 sky130_fd_sc_hd__a221o_1 _0663_ (.A1(net129),
    .A2(_0232_),
    .B1(_0250_),
    .B2(net74),
    .C1(_0280_),
    .X(_0288_));
 sky130_fd_sc_hd__a221o_1 _0664_ (.A1(net29),
    .A2(_0237_),
    .B1(_0287_),
    .B2(net12),
    .C1(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__a211o_2 _0665_ (.A1(net120),
    .A2(_0242_),
    .B1(_0286_),
    .C1(_0289_),
    .X(net291));
 sky130_fd_sc_hd__a21o_1 _0666_ (.A1(_0222_),
    .A2(_0230_),
    .B1(_0235_),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_2 _0667_ (.A1(net162),
    .A2(_0255_),
    .B1(_0290_),
    .B2(_0234_),
    .X(_0291_));
 sky130_fd_sc_hd__a221o_1 _0668_ (.A1(net130),
    .A2(_0232_),
    .B1(_0250_),
    .B2(net82),
    .C1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__a22o_1 _0669_ (.A1(net109),
    .A2(_0228_),
    .B1(_0237_),
    .B2(net30),
    .X(_0293_));
 sky130_fd_sc_hd__a221o_1 _0670_ (.A1(net121),
    .A2(_0242_),
    .B1(_0272_),
    .B2(net55),
    .C1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__a211o_2 _0671_ (.A1(net20),
    .A2(_0287_),
    .B1(_0292_),
    .C1(_0294_),
    .X(net292));
 sky130_fd_sc_hd__a221o_1 _0672_ (.A1(net131),
    .A2(_0232_),
    .B1(_0272_),
    .B2(net56),
    .C1(_0291_),
    .X(_0295_));
 sky130_fd_sc_hd__a22o_1 _0673_ (.A1(net122),
    .A2(_0242_),
    .B1(_0249_),
    .B2(net83),
    .X(_0296_));
 sky130_fd_sc_hd__a221o_1 _0674_ (.A1(net110),
    .A2(_0228_),
    .B1(_0237_),
    .B2(net31),
    .C1(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__a211o_2 _0675_ (.A1(net21),
    .A2(_0287_),
    .B1(_0295_),
    .C1(_0297_),
    .X(net293));
 sky130_fd_sc_hd__a22o_1 _0676_ (.A1(net111),
    .A2(_0227_),
    .B1(_0287_),
    .B2(net22),
    .X(_0298_));
 sky130_fd_sc_hd__a221o_1 _0677_ (.A1(net32),
    .A2(_0237_),
    .B1(_0267_),
    .B2(net137),
    .C1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__a221o_1 _0678_ (.A1(net132),
    .A2(_0232_),
    .B1(_0249_),
    .B2(net84),
    .C1(_0279_),
    .X(_0300_));
 sky130_fd_sc_hd__a221o_1 _0679_ (.A1(net123),
    .A2(_0242_),
    .B1(_0272_),
    .B2(net57),
    .C1(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _0680_ (.A(_0299_),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_2 _0681_ (.A(_0302_),
    .X(net294));
 sky130_fd_sc_hd__a22o_1 _0682_ (.A1(net112),
    .A2(_0226_),
    .B1(_0282_),
    .B2(net23),
    .X(_0303_));
 sky130_fd_sc_hd__a221o_1 _0683_ (.A1(net33),
    .A2(_0237_),
    .B1(_0242_),
    .B2(net124),
    .C1(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__a22o_1 _0684_ (.A1(net138),
    .A2(_0267_),
    .B1(_0272_),
    .B2(net58),
    .X(_0305_));
 sky130_fd_sc_hd__a221o_1 _0685_ (.A1(net133),
    .A2(_0232_),
    .B1(_0249_),
    .B2(net85),
    .C1(_0279_),
    .X(_0306_));
 sky130_fd_sc_hd__or3_1 _0686_ (.A(_0304_),
    .B(_0305_),
    .C(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0687_ (.A(_0307_),
    .X(net295));
 sky130_fd_sc_hd__a22o_1 _0688_ (.A1(net34),
    .A2(_0237_),
    .B1(_0267_),
    .B2(net139),
    .X(_0308_));
 sky130_fd_sc_hd__a221o_1 _0689_ (.A1(net134),
    .A2(_0232_),
    .B1(_0271_),
    .B2(net59),
    .C1(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _0690_ (.A1(net113),
    .A2(_0227_),
    .B1(_0242_),
    .B2(net125),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _0691_ (.A1(net154),
    .A2(_0245_),
    .B1(_0282_),
    .B2(net24),
    .X(_0311_));
 sky130_fd_sc_hd__a211o_1 _0692_ (.A1(net86),
    .A2(_0249_),
    .B1(_0291_),
    .C1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__or3_1 _0693_ (.A(_0309_),
    .B(_0310_),
    .C(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_2 _0694_ (.A(_0313_),
    .X(net296));
 sky130_fd_sc_hd__a22o_1 _0695_ (.A1(net155),
    .A2(_0245_),
    .B1(_0257_),
    .B2(net25),
    .X(_0314_));
 sky130_fd_sc_hd__a221o_1 _0696_ (.A1(net140),
    .A2(_0267_),
    .B1(_0271_),
    .B2(net60),
    .C1(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__a22o_1 _0697_ (.A1(net35),
    .A2(_0236_),
    .B1(_0241_),
    .B2(net126),
    .X(_0316_));
 sky130_fd_sc_hd__a22o_1 _0698_ (.A1(net114),
    .A2(_0226_),
    .B1(_0231_),
    .B2(net135),
    .X(_0317_));
 sky130_fd_sc_hd__a211o_1 _0699_ (.A1(net87),
    .A2(_0249_),
    .B1(_0316_),
    .C1(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__or3_1 _0700_ (.A(_0280_),
    .B(_0315_),
    .C(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_2 _0701_ (.A(_0319_),
    .X(net297));
 sky130_fd_sc_hd__a22o_1 _0702_ (.A1(net127),
    .A2(_0241_),
    .B1(_0245_),
    .B2(net156),
    .X(_0320_));
 sky130_fd_sc_hd__a221o_1 _0703_ (.A1(net141),
    .A2(_0267_),
    .B1(_0249_),
    .B2(net88),
    .C1(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__a221o_1 _0704_ (.A1(net136),
    .A2(_0232_),
    .B1(_0287_),
    .B2(net26),
    .C1(_0291_),
    .X(_0322_));
 sky130_fd_sc_hd__a211o_1 _0705_ (.A1(net115),
    .A2(_0228_),
    .B1(_0321_),
    .C1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__a221o_2 _0706_ (.A1(net61),
    .A2(_0272_),
    .B1(_0277_),
    .B2(net146),
    .C1(_0323_),
    .X(net298));
 sky130_fd_sc_hd__a22o_1 _0707_ (.A1(net116),
    .A2(_0226_),
    .B1(_0270_),
    .B2(net62),
    .X(_0324_));
 sky130_fd_sc_hd__a221o_1 _0708_ (.A1(net142),
    .A2(_0267_),
    .B1(_0277_),
    .B2(net147),
    .C1(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__a221o_1 _0709_ (.A1(net157),
    .A2(_0245_),
    .B1(_0248_),
    .B2(net89),
    .C1(_0279_),
    .X(_0326_));
 sky130_fd_sc_hd__a221o_1 _0710_ (.A1(net128),
    .A2(_0241_),
    .B1(_0287_),
    .B2(net27),
    .C1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _0711_ (.A(_0325_),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_2 _0712_ (.A(_0328_),
    .X(net299));
 sky130_fd_sc_hd__a22o_1 _0713_ (.A1(net143),
    .A2(_0267_),
    .B1(_0241_),
    .B2(net118),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _0714_ (.A(_0232_),
    .B(_0279_),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _0715_ (.A1(net91),
    .A2(_0226_),
    .B1(_0277_),
    .B2(net148),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_1 _0716_ (.A1(net158),
    .A2(_0244_),
    .B1(_0247_),
    .B2(net64),
    .X(_0332_));
 sky130_fd_sc_hd__a221o_1 _0717_ (.A1(net2),
    .A2(_0282_),
    .B1(_0270_),
    .B2(net37),
    .C1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__or4_1 _0718_ (.A(_0329_),
    .B(_0330_),
    .C(_0331_),
    .D(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_2 _0719_ (.A(_0334_),
    .X(net300));
 sky130_fd_sc_hd__a22o_1 _0720_ (.A1(net3),
    .A2(_0257_),
    .B1(_0277_),
    .B2(net149),
    .X(_0335_));
 sky130_fd_sc_hd__a221o_1 _0721_ (.A1(net144),
    .A2(_0267_),
    .B1(_0242_),
    .B2(net119),
    .C1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__a221o_1 _0722_ (.A1(net159),
    .A2(_0245_),
    .B1(_0248_),
    .B2(net65),
    .C1(_0279_),
    .X(_0337_));
 sky130_fd_sc_hd__a221o_1 _0723_ (.A1(net92),
    .A2(_0227_),
    .B1(_0271_),
    .B2(net38),
    .C1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _0724_ (.A(_0336_),
    .B(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0725_ (.A(_0339_),
    .X(net301));
 sky130_fd_sc_hd__a22o_1 _0726_ (.A1(net145),
    .A2(_0266_),
    .B1(_0277_),
    .B2(net150),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _0727_ (.A(_0231_),
    .B(_0291_),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _0728_ (.A1(net160),
    .A2(_0245_),
    .B1(_0282_),
    .B2(net4),
    .X(_0342_));
 sky130_fd_sc_hd__a2111o_1 _0729_ (.A1(net39),
    .A2(_0271_),
    .B1(_0340_),
    .C1(_0341_),
    .D1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__a221o_2 _0730_ (.A1(net93),
    .A2(_0228_),
    .B1(_0250_),
    .B2(net66),
    .C1(_0343_),
    .X(net302));
 sky130_fd_sc_hd__a22o_1 _0731_ (.A1(net161),
    .A2(_0245_),
    .B1(_0277_),
    .B2(net151),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_1 _0732_ (.A1(net94),
    .A2(_0226_),
    .B1(_0282_),
    .B2(net5),
    .X(_0345_));
 sky130_fd_sc_hd__a221o_1 _0733_ (.A1(net67),
    .A2(_0248_),
    .B1(_0270_),
    .B2(net40),
    .C1(_0291_),
    .X(_0346_));
 sky130_fd_sc_hd__or3_1 _0734_ (.A(_0344_),
    .B(_0345_),
    .C(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_2 _0735_ (.A(_0347_),
    .X(net303));
 sky130_fd_sc_hd__a22o_1 _0736_ (.A1(net95),
    .A2(_0226_),
    .B1(_0277_),
    .B2(net152),
    .X(_0348_));
 sky130_fd_sc_hd__a221o_1 _0737_ (.A1(net6),
    .A2(_0287_),
    .B1(_0272_),
    .B2(net41),
    .C1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__a211o_2 _0738_ (.A1(net68),
    .A2(_0250_),
    .B1(_0330_),
    .C1(_0349_),
    .X(net304));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(net96),
    .A2(_0228_),
    .B1(_0287_),
    .B2(net7),
    .X(_0350_));
 sky130_fd_sc_hd__a221o_1 _0740_ (.A1(net42),
    .A2(_0272_),
    .B1(_0277_),
    .B2(net153),
    .C1(_0280_),
    .X(_0351_));
 sky130_fd_sc_hd__a211o_2 _0741_ (.A1(net69),
    .A2(_0250_),
    .B1(_0350_),
    .C1(_0351_),
    .X(net305));
 sky130_fd_sc_hd__a22o_1 _0742_ (.A1(net97),
    .A2(_0226_),
    .B1(_0248_),
    .B2(net70),
    .X(_0352_));
 sky130_fd_sc_hd__a221o_1 _0743_ (.A1(net8),
    .A2(_0282_),
    .B1(_0271_),
    .B2(net43),
    .C1(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _0744_ (.A(_0341_),
    .B(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_2 _0745_ (.A(_0354_),
    .X(net306));
 sky130_fd_sc_hd__a22o_1 _0746_ (.A1(net9),
    .A2(_0257_),
    .B1(_0270_),
    .B2(net44),
    .X(_0355_));
 sky130_fd_sc_hd__a221o_1 _0747_ (.A1(net98),
    .A2(_0227_),
    .B1(_0249_),
    .B2(net71),
    .C1(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _0748_ (.A(_0280_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_2 _0749_ (.A(_0357_),
    .X(net307));
 sky130_fd_sc_hd__a22o_1 _0750_ (.A1(net72),
    .A2(_0248_),
    .B1(_0270_),
    .B2(net45),
    .X(_0358_));
 sky130_fd_sc_hd__a221o_1 _0751_ (.A1(net99),
    .A2(_0227_),
    .B1(_0282_),
    .B2(net10),
    .C1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _0752_ (.A(_0341_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_2 _0753_ (.A(_0360_),
    .X(net308));
 sky130_fd_sc_hd__a22o_1 _0754_ (.A1(net11),
    .A2(_0257_),
    .B1(_0270_),
    .B2(net46),
    .X(_0361_));
 sky130_fd_sc_hd__a221o_1 _0755_ (.A1(net100),
    .A2(_0227_),
    .B1(_0249_),
    .B2(net73),
    .C1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__or2_1 _0756_ (.A(_0280_),
    .B(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_2 _0757_ (.A(_0363_),
    .X(net309));
 sky130_fd_sc_hd__a22o_1 _0758_ (.A1(net102),
    .A2(_0226_),
    .B1(_0270_),
    .B2(net48),
    .X(_0364_));
 sky130_fd_sc_hd__a221o_1 _0759_ (.A1(net75),
    .A2(_0248_),
    .B1(_0282_),
    .B2(net13),
    .C1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or2_1 _0760_ (.A(_0330_),
    .B(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_2 _0761_ (.A(_0366_),
    .X(net310));
 sky130_fd_sc_hd__a22o_1 _0762_ (.A1(net14),
    .A2(_0257_),
    .B1(_0270_),
    .B2(net49),
    .X(_0367_));
 sky130_fd_sc_hd__a221o_1 _0763_ (.A1(net103),
    .A2(_0227_),
    .B1(_0248_),
    .B2(net76),
    .C1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__or2_1 _0764_ (.A(_0280_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_2 _0765_ (.A(_0369_),
    .X(net311));
 sky130_fd_sc_hd__a22o_1 _0766_ (.A1(net77),
    .A2(_0248_),
    .B1(_0257_),
    .B2(net15),
    .X(_0370_));
 sky130_fd_sc_hd__a221o_1 _0767_ (.A1(net104),
    .A2(_0227_),
    .B1(_0271_),
    .B2(net50),
    .C1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _0768_ (.A(_0341_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_2 _0769_ (.A(_0372_),
    .X(net312));
 sky130_fd_sc_hd__a22o_1 _0770_ (.A1(net16),
    .A2(_0257_),
    .B1(_0270_),
    .B2(net51),
    .X(_0373_));
 sky130_fd_sc_hd__a221o_1 _0771_ (.A1(net105),
    .A2(_0226_),
    .B1(_0248_),
    .B2(net78),
    .C1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _0772_ (.A(_0280_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_2 _0773_ (.A(_0375_),
    .X(net313));
 sky130_fd_sc_hd__a22o_1 _0774_ (.A1(net106),
    .A2(_0227_),
    .B1(_0271_),
    .B2(net52),
    .X(_0376_));
 sky130_fd_sc_hd__a221o_1 _0775_ (.A1(net79),
    .A2(_0250_),
    .B1(_0287_),
    .B2(net17),
    .C1(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(_0330_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_2 _0777_ (.A(_0378_),
    .X(net314));
 sky130_fd_sc_hd__a22o_1 _0778_ (.A1(net18),
    .A2(_0287_),
    .B1(_0271_),
    .B2(net53),
    .X(_0379_));
 sky130_fd_sc_hd__a221o_1 _0779_ (.A1(net107),
    .A2(_0228_),
    .B1(_0250_),
    .B2(net80),
    .C1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__or2_1 _0780_ (.A(_0280_),
    .B(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_2 _0781_ (.A(_0381_),
    .X(net315));
 sky130_fd_sc_hd__a22o_1 _0782_ (.A1(net19),
    .A2(_0282_),
    .B1(_0271_),
    .B2(net54),
    .X(_0382_));
 sky130_fd_sc_hd__a221o_1 _0783_ (.A1(net108),
    .A2(_0228_),
    .B1(_0250_),
    .B2(net81),
    .C1(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__or2_1 _0784_ (.A(_0280_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_2 _0785_ (.A(_0384_),
    .X(net316));
 sky130_fd_sc_hd__mux2_2 _0786_ (.A0(clknet_3_0__leaf_wb_clk_i),
    .A1(wb_clk_override),
    .S(wb_single_step),
    .X(_0385_));
 sky130_fd_sc_hd__buf_2 _0787_ (.A(wb_override),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_2 _0788_ (.A0(net163),
    .A1(_0385_),
    .S(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_1 _0789_ (.A(_0387_),
    .X(net235));
 sky130_fd_sc_hd__buf_2 _0790_ (.A(_0386_),
    .X(_0388_));
 sky130_fd_sc_hd__buf_2 _0791_ (.A(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__and2b_1 _0792_ (.A_N(_0388_),
    .B(net164),
    .X(_0390_));
 sky130_fd_sc_hd__a31o_1 _0793_ (.A1(_0389_),
    .A2(\wb_io_override[0] ),
    .A3(net263),
    .B1(_0390_),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 _0794_ (.A(_0386_),
    .X(_0391_));
 sky130_fd_sc_hd__and2b_1 _0795_ (.A_N(_0391_),
    .B(net165),
    .X(_0392_));
 sky130_fd_sc_hd__a31o_1 _0796_ (.A1(_0389_),
    .A2(\wb_io_override[1] ),
    .A3(net266),
    .B1(_0392_),
    .X(net247));
 sky130_fd_sc_hd__and2b_1 _0797_ (.A_N(_0391_),
    .B(net166),
    .X(_0393_));
 sky130_fd_sc_hd__a31o_1 _0798_ (.A1(_0389_),
    .A2(\wb_io_override[2] ),
    .A3(net266),
    .B1(_0393_),
    .X(net255));
 sky130_fd_sc_hd__and2b_1 _0799_ (.A_N(_0391_),
    .B(net167),
    .X(_0394_));
 sky130_fd_sc_hd__a31o_1 _0800_ (.A1(_0389_),
    .A2(\wb_io_override[3] ),
    .A3(net266),
    .B1(_0394_),
    .X(net256));
 sky130_fd_sc_hd__and2b_1 _0801_ (.A_N(_0391_),
    .B(net168),
    .X(_0395_));
 sky130_fd_sc_hd__a31o_1 _0802_ (.A1(_0389_),
    .A2(\wb_io_override[4] ),
    .A3(net267),
    .B1(_0395_),
    .X(net257));
 sky130_fd_sc_hd__and2b_1 _0803_ (.A_N(_0391_),
    .B(net169),
    .X(_0396_));
 sky130_fd_sc_hd__a31o_1 _0804_ (.A1(_0389_),
    .A2(\wb_io_override[5] ),
    .A3(net268),
    .B1(_0396_),
    .X(net258));
 sky130_fd_sc_hd__and2b_1 _0805_ (.A_N(_0391_),
    .B(net170),
    .X(_0397_));
 sky130_fd_sc_hd__a31o_1 _0806_ (.A1(_0389_),
    .A2(\wb_io_override[6] ),
    .A3(net270),
    .B1(_0397_),
    .X(net259));
 sky130_fd_sc_hd__and2b_1 _0807_ (.A_N(_0391_),
    .B(net171),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_1 _0808_ (.A1(_0389_),
    .A2(\wb_io_override[7] ),
    .A3(net270),
    .B1(_0398_),
    .X(net260));
 sky130_fd_sc_hd__and2b_1 _0809_ (.A_N(_0391_),
    .B(net172),
    .X(_0399_));
 sky130_fd_sc_hd__a31o_1 _0810_ (.A1(_0389_),
    .A2(\wb_io_override[8] ),
    .A3(net272),
    .B1(_0399_),
    .X(net261));
 sky130_fd_sc_hd__and2b_1 _0811_ (.A_N(_0391_),
    .B(net173),
    .X(_0400_));
 sky130_fd_sc_hd__a31o_1 _0812_ (.A1(_0389_),
    .A2(\wb_io_override[9] ),
    .A3(net272),
    .B1(_0400_),
    .X(net262));
 sky130_fd_sc_hd__buf_2 _0813_ (.A(_0388_),
    .X(_0401_));
 sky130_fd_sc_hd__and2b_1 _0814_ (.A_N(_0391_),
    .B(net174),
    .X(_0402_));
 sky130_fd_sc_hd__a31o_1 _0815_ (.A1(_0401_),
    .A2(\wb_io_override[10] ),
    .A3(net274),
    .B1(_0402_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 _0816_ (.A(wb_override),
    .X(_0403_));
 sky130_fd_sc_hd__and2b_1 _0817_ (.A_N(_0403_),
    .B(net175),
    .X(_0404_));
 sky130_fd_sc_hd__a31o_1 _0818_ (.A1(_0401_),
    .A2(\wb_io_override[11] ),
    .A3(net274),
    .B1(_0404_),
    .X(net238));
 sky130_fd_sc_hd__and2b_1 _0819_ (.A_N(_0403_),
    .B(net176),
    .X(_0405_));
 sky130_fd_sc_hd__a31o_1 _0820_ (.A1(_0401_),
    .A2(\wb_io_override[12] ),
    .A3(net275),
    .B1(_0405_),
    .X(net239));
 sky130_fd_sc_hd__and2b_1 _0821_ (.A_N(_0403_),
    .B(net177),
    .X(_0406_));
 sky130_fd_sc_hd__a31o_1 _0822_ (.A1(_0401_),
    .A2(\wb_io_override[13] ),
    .A3(net276),
    .B1(_0406_),
    .X(net240));
 sky130_fd_sc_hd__and2b_1 _0823_ (.A_N(_0403_),
    .B(net178),
    .X(_0407_));
 sky130_fd_sc_hd__a31o_1 _0824_ (.A1(_0401_),
    .A2(\wb_io_override[14] ),
    .A3(net278),
    .B1(_0407_),
    .X(net241));
 sky130_fd_sc_hd__and2b_1 _0825_ (.A_N(_0403_),
    .B(net179),
    .X(_0408_));
 sky130_fd_sc_hd__a31o_1 _0826_ (.A1(_0401_),
    .A2(\wb_io_override[15] ),
    .A3(net278),
    .B1(_0408_),
    .X(net242));
 sky130_fd_sc_hd__and2b_1 _0827_ (.A_N(_0403_),
    .B(net180),
    .X(_0409_));
 sky130_fd_sc_hd__a31o_1 _0828_ (.A1(_0401_),
    .A2(\wb_io_override[16] ),
    .A3(net356),
    .B1(_0409_),
    .X(net243));
 sky130_fd_sc_hd__and2b_1 _0829_ (.A_N(_0403_),
    .B(net181),
    .X(_0410_));
 sky130_fd_sc_hd__a31o_1 _0830_ (.A1(_0401_),
    .A2(\wb_io_override[17] ),
    .A3(net356),
    .B1(_0410_),
    .X(net244));
 sky130_fd_sc_hd__and2b_1 _0831_ (.A_N(_0403_),
    .B(net182),
    .X(_0411_));
 sky130_fd_sc_hd__a31o_1 _0832_ (.A1(_0401_),
    .A2(\wb_io_override[18] ),
    .A3(net356),
    .B1(_0411_),
    .X(net245));
 sky130_fd_sc_hd__and2b_1 _0833_ (.A_N(_0403_),
    .B(net183),
    .X(_0412_));
 sky130_fd_sc_hd__a31o_1 _0834_ (.A1(_0401_),
    .A2(\wb_io_override[19] ),
    .A3(net356),
    .B1(_0412_),
    .X(net246));
 sky130_fd_sc_hd__and2b_1 _0835_ (.A_N(_0403_),
    .B(net184),
    .X(_0413_));
 sky130_fd_sc_hd__a31o_1 _0836_ (.A1(_0388_),
    .A2(\wb_io_override[20] ),
    .A3(net356),
    .B1(_0413_),
    .X(net248));
 sky130_fd_sc_hd__and2b_1 _0837_ (.A_N(_0386_),
    .B(net185),
    .X(_0414_));
 sky130_fd_sc_hd__a31o_1 _0838_ (.A1(_0388_),
    .A2(\wb_io_override[21] ),
    .A3(net356),
    .B1(_0414_),
    .X(net249));
 sky130_fd_sc_hd__and2b_1 _0839_ (.A_N(_0386_),
    .B(net186),
    .X(_0415_));
 sky130_fd_sc_hd__a31o_1 _0840_ (.A1(_0388_),
    .A2(\wb_io_override[22] ),
    .A3(net356),
    .B1(_0415_),
    .X(net250));
 sky130_fd_sc_hd__and2b_1 _0841_ (.A_N(_0386_),
    .B(net187),
    .X(_0416_));
 sky130_fd_sc_hd__a31o_1 _0842_ (.A1(_0388_),
    .A2(\wb_io_override[23] ),
    .A3(net356),
    .B1(_0416_),
    .X(net251));
 sky130_fd_sc_hd__and2b_1 _0843_ (.A_N(_0386_),
    .B(net188),
    .X(_0417_));
 sky130_fd_sc_hd__a31o_1 _0844_ (.A1(_0388_),
    .A2(\wb_io_override[24] ),
    .A3(net356),
    .B1(_0417_),
    .X(net252));
 sky130_fd_sc_hd__and2b_1 _0845_ (.A_N(_0386_),
    .B(net189),
    .X(_0418_));
 sky130_fd_sc_hd__a31o_1 _0846_ (.A1(_0388_),
    .A2(\wb_io_override[25] ),
    .A3(_0278_),
    .B1(_0418_),
    .X(net253));
 sky130_fd_sc_hd__and2b_1 _0847_ (.A_N(_0386_),
    .B(net190),
    .X(_0419_));
 sky130_fd_sc_hd__a31o_1 _0848_ (.A1(_0388_),
    .A2(\wb_io_override[26] ),
    .A3(_0278_),
    .B1(_0419_),
    .X(net254));
 sky130_fd_sc_hd__or2b_1 _0849_ (.A(net234),
    .B_N(net202),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(net203),
    .B(net204),
    .Y(_0421_));
 sky130_fd_sc_hd__nand2_1 _0851_ (.A(net233),
    .B(net205),
    .Y(_0422_));
 sky130_fd_sc_hd__a21o_1 _0852_ (.A1(_0420_),
    .A2(_0421_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__buf_2 _0853_ (.A(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_2 _0854_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__and2_1 _0855_ (.A(net328),
    .B(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_4 _0856_ (.A(net204),
    .X(_0427_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__clkinv_2 _0858_ (.A(_0423_),
    .Y(_0429_));
 sky130_fd_sc_hd__buf_2 _0859_ (.A(net203),
    .X(_0430_));
 sky130_fd_sc_hd__inv_2 _0860_ (.A(net203),
    .Y(_0431_));
 sky130_fd_sc_hd__buf_2 _0861_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__a21o_1 _0862_ (.A1(\wb_counter[0] ),
    .A2(_0432_),
    .B1(_0427_),
    .X(_0433_));
 sky130_fd_sc_hd__a31o_1 _0863_ (.A1(_0430_),
    .A2(_0264_),
    .A3(net290),
    .B1(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o211a_1 _0864_ (.A1(_0386_),
    .A2(_0428_),
    .B1(_0429_),
    .C1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__clkinv_2 _0865_ (.A(net201),
    .Y(_0436_));
 sky130_fd_sc_hd__clkbuf_2 _0866_ (.A(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__o21a_1 _0867_ (.A1(_0426_),
    .A2(_0435_),
    .B1(_0437_),
    .X(_0000_));
 sky130_fd_sc_hd__and4_1 _0868_ (.A(_0430_),
    .B(_0428_),
    .C(_0264_),
    .D(net291),
    .X(_0438_));
 sky130_fd_sc_hd__a221o_1 _0869_ (.A1(wb_rst_override),
    .A2(_0427_),
    .B1(_0421_),
    .B2(\wb_counter[1] ),
    .C1(_0425_),
    .X(_0439_));
 sky130_fd_sc_hd__o221a_1 _0870_ (.A1(net339),
    .A2(_0429_),
    .B1(_0438_),
    .B2(_0439_),
    .C1(_0437_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(net347),
    .B(_0425_),
    .X(_0440_));
 sky130_fd_sc_hd__a21o_1 _0872_ (.A1(\wb_counter[2] ),
    .A2(_0432_),
    .B1(_0427_),
    .X(_0441_));
 sky130_fd_sc_hd__a31o_1 _0873_ (.A1(_0430_),
    .A2(_0264_),
    .A3(net292),
    .B1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__o211a_1 _0874_ (.A1(\wb_design_addr_override[0] ),
    .A2(_0428_),
    .B1(_0429_),
    .C1(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__o21a_1 _0875_ (.A1(_0440_),
    .A2(_0443_),
    .B1(_0437_),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _0876_ (.A(net348),
    .B(_0425_),
    .X(_0444_));
 sky130_fd_sc_hd__a21o_1 _0877_ (.A1(\wb_counter[3] ),
    .A2(_0432_),
    .B1(_0427_),
    .X(_0445_));
 sky130_fd_sc_hd__a31o_1 _0878_ (.A1(_0430_),
    .A2(_0264_),
    .A3(net293),
    .B1(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__o211a_1 _0879_ (.A1(\wb_design_addr_override[1] ),
    .A2(_0428_),
    .B1(_0429_),
    .C1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__o21a_1 _0880_ (.A1(_0444_),
    .A2(_0447_),
    .B1(_0437_),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_1 _0881_ (.A(_0432_),
    .B(net267),
    .Y(_0448_));
 sky130_fd_sc_hd__or2_1 _0882_ (.A(_0427_),
    .B(_0424_),
    .X(_0449_));
 sky130_fd_sc_hd__a221o_1 _0883_ (.A1(\wb_counter[4] ),
    .A2(_0432_),
    .B1(net294),
    .B2(_0448_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_4 _0884_ (.A(_0436_),
    .X(_0451_));
 sky130_fd_sc_hd__o21a_1 _0885_ (.A1(net349),
    .A2(_0429_),
    .B1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__o311a_1 _0886_ (.A1(\wb_design_addr_override[2] ),
    .A2(_0428_),
    .A3(_0425_),
    .B1(_0450_),
    .C1(_0452_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _0887_ (.A(net350),
    .B(_0425_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _0888_ (.A(_0432_),
    .B(net268),
    .Y(_0454_));
 sky130_fd_sc_hd__a221o_1 _0889_ (.A1(\wb_counter[5] ),
    .A2(_0432_),
    .B1(net295),
    .B2(_0454_),
    .C1(_0427_),
    .X(_0455_));
 sky130_fd_sc_hd__o211a_1 _0890_ (.A1(\wb_design_addr_override[3] ),
    .A2(_0428_),
    .B1(_0429_),
    .C1(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__o21a_1 _0891_ (.A1(_0453_),
    .A2(_0456_),
    .B1(_0437_),
    .X(_0005_));
 sky130_fd_sc_hd__nor2_1 _0892_ (.A(_0431_),
    .B(net270),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _0893_ (.A(net412),
    .Y(_0458_));
 sky130_fd_sc_hd__o2bb2a_1 _0894_ (.A1_N(net296),
    .A2_N(_0457_),
    .B1(_0458_),
    .B2(_0430_),
    .X(_0459_));
 sky130_fd_sc_hd__o2bb2a_1 _0895_ (.A1_N(net351),
    .A2_N(_0425_),
    .B1(_0449_),
    .B2(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _0896_ (.A(net201),
    .B(_0460_),
    .Y(_0006_));
 sky130_fd_sc_hd__nor2_2 _0897_ (.A(_0427_),
    .B(_0423_),
    .Y(_0461_));
 sky130_fd_sc_hd__buf_2 _0898_ (.A(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _0899_ (.A1(\wb_counter[7] ),
    .A2(_0432_),
    .B1(net297),
    .B2(_0457_),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _0900_ (.A1(net352),
    .A2(_0425_),
    .B1(_0462_),
    .B2(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _0901_ (.A(_0437_),
    .B(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0902_ (.A(_0465_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _0903_ (.A(_0431_),
    .B(net272),
    .Y(_0466_));
 sky130_fd_sc_hd__a22oi_1 _0904_ (.A1(\wb_counter[8] ),
    .A2(_0432_),
    .B1(net298),
    .B2(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__o2bb2a_1 _0905_ (.A1_N(net353),
    .A2_N(_0425_),
    .B1(_0449_),
    .B2(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_1 _0906_ (.A(net201),
    .B(_0468_),
    .Y(_0008_));
 sky130_fd_sc_hd__buf_2 _0907_ (.A(_0424_),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _0908_ (.A1(\wb_counter[9] ),
    .A2(_0431_),
    .B1(net299),
    .B2(_0466_),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _0909_ (.A1(net354),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__and2_1 _0910_ (.A(_0437_),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0472_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _0912_ (.A(\wb_counter[10] ),
    .B(_0431_),
    .X(_0473_));
 sky130_fd_sc_hd__a31o_1 _0913_ (.A1(_0430_),
    .A2(_0273_),
    .A3(net300),
    .B1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _0914_ (.A1(net329),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__and2_1 _0915_ (.A(_0437_),
    .B(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _0916_ (.A(_0476_),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(\wb_counter[11] ),
    .B(_0431_),
    .X(_0477_));
 sky130_fd_sc_hd__a31o_1 _0918_ (.A1(_0430_),
    .A2(_0273_),
    .A3(net301),
    .B1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _0919_ (.A1(net330),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__and2_1 _0920_ (.A(_0437_),
    .B(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0480_),
    .X(_0011_));
 sky130_fd_sc_hd__a21o_1 _0922_ (.A1(_0274_),
    .A2(net302),
    .B1(_0432_),
    .X(_0481_));
 sky130_fd_sc_hd__or2_1 _0923_ (.A(\wb_counter[12] ),
    .B(_0430_),
    .X(_0482_));
 sky130_fd_sc_hd__a32o_1 _0924_ (.A1(_0461_),
    .A2(_0481_),
    .A3(_0482_),
    .B1(_0425_),
    .B2(net331),
    .X(_0483_));
 sky130_fd_sc_hd__and2_1 _0925_ (.A(_0437_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _0926_ (.A(_0484_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_2 _0927_ (.A(_0436_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(\wb_counter[13] ),
    .A1(net303),
    .S(_0430_),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _0929_ (.A1(net332),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__and2_1 _0930_ (.A(_0485_),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _0931_ (.A(_0488_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _0932_ (.A(net203),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(\wb_counter[14] ),
    .A1(net304),
    .S(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _0934_ (.A1(net333),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__and2_1 _0935_ (.A(_0485_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _0936_ (.A(_0492_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(\wb_counter[15] ),
    .A1(net305),
    .S(_0489_),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _0938_ (.A1(net334),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _0939_ (.A(_0485_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _0940_ (.A(_0495_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0941_ (.A0(\wb_counter[16] ),
    .A1(net306),
    .S(_0489_),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _0942_ (.A1(net335),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__and2_1 _0943_ (.A(_0485_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _0944_ (.A(_0498_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0945_ (.A0(\wb_counter[17] ),
    .A1(net307),
    .S(_0489_),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _0946_ (.A1(net336),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__and2_1 _0947_ (.A(_0485_),
    .B(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _0948_ (.A(_0501_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(\wb_counter[18] ),
    .A1(net308),
    .S(_0489_),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _0950_ (.A1(net337),
    .A2(_0469_),
    .B1(_0462_),
    .B2(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(_0485_),
    .B(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _0952_ (.A(_0504_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(\wb_counter[19] ),
    .A1(net309),
    .S(_0489_),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _0954_ (.A1(net338),
    .A2(_0469_),
    .B1(_0461_),
    .B2(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(_0485_),
    .B(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _0956_ (.A(_0507_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0957_ (.A0(\wb_counter[20] ),
    .A1(net310),
    .S(_0489_),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_1 _0958_ (.A1(net340),
    .A2(_0424_),
    .B1(_0461_),
    .B2(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__and2_1 _0959_ (.A(_0485_),
    .B(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__clkbuf_1 _0960_ (.A(_0510_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(\wb_counter[21] ),
    .A1(net311),
    .S(_0489_),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _0962_ (.A1(net341),
    .A2(_0424_),
    .B1(_0461_),
    .B2(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__and2_1 _0963_ (.A(_0485_),
    .B(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__clkbuf_1 _0964_ (.A(_0513_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(\wb_counter[22] ),
    .A1(net312),
    .S(_0489_),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _0966_ (.A1(net342),
    .A2(_0424_),
    .B1(_0461_),
    .B2(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__and2_1 _0967_ (.A(_0485_),
    .B(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _0968_ (.A(_0516_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_2 _0969_ (.A(_0436_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(\wb_counter[23] ),
    .A1(net313),
    .S(_0489_),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _0971_ (.A1(net343),
    .A2(_0424_),
    .B1(_0461_),
    .B2(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__and2_1 _0972_ (.A(_0517_),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _0973_ (.A(_0520_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _0974_ (.A(_0430_),
    .B(_0428_),
    .C(_0429_),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _0975_ (.A1(net344),
    .A2(_0424_),
    .B1(_0521_),
    .B2(net314),
    .X(_0522_));
 sky130_fd_sc_hd__and2_1 _0976_ (.A(_0517_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0523_),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_1 _0978_ (.A1(net345),
    .A2(_0424_),
    .B1(_0521_),
    .B2(net315),
    .X(_0524_));
 sky130_fd_sc_hd__and2_1 _0979_ (.A(_0517_),
    .B(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(_0525_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _0981_ (.A1(net346),
    .A2(_0424_),
    .B1(_0521_),
    .B2(net316),
    .X(_0526_));
 sky130_fd_sc_hd__and2_1 _0982_ (.A(_0517_),
    .B(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0527_),
    .X(_0026_));
 sky130_fd_sc_hd__xnor2_1 _0984_ (.A(net410),
    .B(net201),
    .Y(_0027_));
 sky130_fd_sc_hd__nand2_1 _0985_ (.A(net410),
    .B(_0451_),
    .Y(_0528_));
 sky130_fd_sc_hd__xnor2_1 _0986_ (.A(net408),
    .B(_0528_),
    .Y(_0028_));
 sky130_fd_sc_hd__and4b_1 _0987_ (.A_N(net201),
    .B(net410),
    .C(net408),
    .D(net438),
    .X(_0529_));
 sky130_fd_sc_hd__a31o_1 _0988_ (.A1(net408),
    .A2(net410),
    .A3(_0436_),
    .B1(net438),
    .X(_0530_));
 sky130_fd_sc_hd__and2b_1 _0989_ (.A_N(_0529_),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(_0531_),
    .X(_0029_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(net430),
    .B(_0529_),
    .Y(_0532_));
 sky130_fd_sc_hd__or2_1 _0992_ (.A(net430),
    .B(_0529_),
    .X(_0533_));
 sky130_fd_sc_hd__and2_1 _0993_ (.A(net431),
    .B(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(net432),
    .X(_0030_));
 sky130_fd_sc_hd__xnor2_1 _0995_ (.A(net403),
    .B(_0532_),
    .Y(_0031_));
 sky130_fd_sc_hd__and4_1 _0996_ (.A(net436),
    .B(net403),
    .C(net430),
    .D(_0529_),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_2 _0997_ (.A(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__a31o_1 _0998_ (.A1(net403),
    .A2(net430),
    .A3(_0529_),
    .B1(net436),
    .X(_0537_));
 sky130_fd_sc_hd__and2b_1 _0999_ (.A_N(_0536_),
    .B(net437),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(_0538_),
    .X(_0032_));
 sky130_fd_sc_hd__xnor2_1 _1001_ (.A(net413),
    .B(_0536_),
    .Y(_0033_));
 sky130_fd_sc_hd__and2_1 _1002_ (.A(net405),
    .B(net412),
    .X(_0539_));
 sky130_fd_sc_hd__and2_1 _1003_ (.A(_0536_),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__a21oi_1 _1004_ (.A1(\wb_counter[6] ),
    .A2(_0536_),
    .B1(net405),
    .Y(_0541_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(_0540_),
    .B(net406),
    .Y(_0034_));
 sky130_fd_sc_hd__xor2_1 _1006_ (.A(net401),
    .B(_0540_),
    .X(_0035_));
 sky130_fd_sc_hd__and2_1 _1007_ (.A(net433),
    .B(net401),
    .X(_0542_));
 sky130_fd_sc_hd__and3_1 _1008_ (.A(_0536_),
    .B(_0539_),
    .C(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a31o_1 _1009_ (.A1(net401),
    .A2(_0536_),
    .A3(_0539_),
    .B1(net433),
    .X(_0544_));
 sky130_fd_sc_hd__and2b_1 _1010_ (.A_N(_0543_),
    .B(net434),
    .X(_0545_));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(net435),
    .X(_0036_));
 sky130_fd_sc_hd__and4_1 _1012_ (.A(net392),
    .B(_0536_),
    .C(_0539_),
    .D(_0542_),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(net392),
    .B(_0543_),
    .Y(_0547_));
 sky130_fd_sc_hd__nor2_1 _1014_ (.A(_0546_),
    .B(net393),
    .Y(_0037_));
 sky130_fd_sc_hd__xor2_1 _1015_ (.A(net399),
    .B(_0546_),
    .X(_0038_));
 sky130_fd_sc_hd__nand2_1 _1016_ (.A(net399),
    .B(_0546_),
    .Y(_0548_));
 sky130_fd_sc_hd__xnor2_1 _1017_ (.A(net388),
    .B(_0548_),
    .Y(_0039_));
 sky130_fd_sc_hd__and4_1 _1018_ (.A(net421),
    .B(net388),
    .C(net399),
    .D(_0546_),
    .X(_0549_));
 sky130_fd_sc_hd__a31o_1 _1019_ (.A1(net388),
    .A2(net399),
    .A3(_0546_),
    .B1(net421),
    .X(_0550_));
 sky130_fd_sc_hd__and2b_1 _1020_ (.A_N(_0549_),
    .B(net422),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(_0551_),
    .X(_0040_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(net429),
    .B(_0549_),
    .Y(_0552_));
 sky130_fd_sc_hd__or2_1 _1023_ (.A(net429),
    .B(_0549_),
    .X(_0553_));
 sky130_fd_sc_hd__and2_1 _1024_ (.A(_0552_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(_0554_),
    .X(_0041_));
 sky130_fd_sc_hd__xnor2_1 _1026_ (.A(net397),
    .B(_0552_),
    .Y(_0042_));
 sky130_fd_sc_hd__and4_1 _1027_ (.A(net423),
    .B(net397),
    .C(\wb_counter[14] ),
    .D(_0549_),
    .X(_0555_));
 sky130_fd_sc_hd__a31o_1 _1028_ (.A1(net397),
    .A2(\wb_counter[14] ),
    .A3(_0549_),
    .B1(net423),
    .X(_0556_));
 sky130_fd_sc_hd__and2b_1 _1029_ (.A_N(_0555_),
    .B(net424),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(net425),
    .X(_0043_));
 sky130_fd_sc_hd__nand2_1 _1031_ (.A(net415),
    .B(_0555_),
    .Y(_0558_));
 sky130_fd_sc_hd__or2_1 _1032_ (.A(net415),
    .B(_0555_),
    .X(_0559_));
 sky130_fd_sc_hd__and2_1 _1033_ (.A(net416),
    .B(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(net417),
    .X(_0044_));
 sky130_fd_sc_hd__xnor2_1 _1035_ (.A(net386),
    .B(_0558_),
    .Y(_0045_));
 sky130_fd_sc_hd__and4_1 _1036_ (.A(net426),
    .B(net386),
    .C(net415),
    .D(_0555_),
    .X(_0561_));
 sky130_fd_sc_hd__a31o_1 _1037_ (.A1(net386),
    .A2(net415),
    .A3(_0555_),
    .B1(net426),
    .X(_0562_));
 sky130_fd_sc_hd__and2b_1 _1038_ (.A_N(_0561_),
    .B(net427),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _1039_ (.A(net428),
    .X(_0046_));
 sky130_fd_sc_hd__xor2_1 _1040_ (.A(net395),
    .B(_0561_),
    .X(_0047_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(net395),
    .B(_0561_),
    .Y(_0564_));
 sky130_fd_sc_hd__xnor2_1 _1042_ (.A(net390),
    .B(_0564_),
    .Y(_0048_));
 sky130_fd_sc_hd__and4_1 _1043_ (.A(net418),
    .B(net390),
    .C(net395),
    .D(_0561_),
    .X(_0565_));
 sky130_fd_sc_hd__a31o_1 _1044_ (.A1(net390),
    .A2(net395),
    .A3(_0561_),
    .B1(net418),
    .X(_0566_));
 sky130_fd_sc_hd__and2b_1 _1045_ (.A_N(_0565_),
    .B(net419),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _1046_ (.A(net420),
    .X(_0049_));
 sky130_fd_sc_hd__xor2_1 _1047_ (.A(net384),
    .B(_0565_),
    .X(_0050_));
 sky130_fd_sc_hd__and3_2 _1048_ (.A(net233),
    .B(net205),
    .C(net234),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_2 _1049_ (.A(_0427_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(net217),
    .A1(wb_rst_override),
    .S(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__and2_1 _1051_ (.A(_0517_),
    .B(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _1052_ (.A(_0571_),
    .X(_0051_));
 sky130_fd_sc_hd__nor2_1 _1053_ (.A(net201),
    .B(_0569_),
    .Y(_0572_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(wb_clk_override),
    .A1(net226),
    .S(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__clkbuf_1 _1055_ (.A(_0573_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(net206),
    .A1(wb_override),
    .S(_0569_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _1057_ (.A(_0517_),
    .B(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _1058_ (.A(_0117_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1059_ (.A0(net227),
    .A1(\wb_design_addr_override[0] ),
    .S(_0569_),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _1060_ (.A(_0517_),
    .B(_0118_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0119_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1062_ (.A0(net228),
    .A1(\wb_design_addr_override[1] ),
    .S(_0569_),
    .X(_0120_));
 sky130_fd_sc_hd__and2_1 _1063_ (.A(_0517_),
    .B(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_1 _1064_ (.A(_0121_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1065_ (.A0(net229),
    .A1(\wb_design_addr_override[2] ),
    .S(_0569_),
    .X(_0122_));
 sky130_fd_sc_hd__and2_1 _1066_ (.A(_0517_),
    .B(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_1 _1067_ (.A(_0123_),
    .X(_0056_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(\wb_design_addr_override[3] ),
    .Y(_0124_));
 sky130_fd_sc_hd__a21oi_1 _1069_ (.A1(_0124_),
    .A2(_0569_),
    .B1(net201),
    .Y(_0125_));
 sky130_fd_sc_hd__o21a_1 _1070_ (.A1(net230),
    .A2(_0569_),
    .B1(_0125_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1071_ (.A0(wb_single_step),
    .A1(net225),
    .S(_0572_),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _1072_ (.A(_0126_),
    .X(_0058_));
 sky130_fd_sc_hd__nor2_1 _1073_ (.A(net201),
    .B(_0422_),
    .Y(_0059_));
 sky130_fd_sc_hd__and3_1 _1074_ (.A(net202),
    .B(_0421_),
    .C(_0568_),
    .X(_0127_));
 sky130_fd_sc_hd__buf_2 _1075_ (.A(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_4 _1076_ (.A(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1077_ (.A0(\wb_counter[0] ),
    .A1(net206),
    .S(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__and2_1 _1078_ (.A(_0517_),
    .B(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _1079_ (.A(_0131_),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_2 _1080_ (.A(_0436_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1081_ (.A0(\wb_counter[1] ),
    .A1(net217),
    .S(_0129_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_1 _1082_ (.A(_0132_),
    .B(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _1083_ (.A(_0134_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(\wb_counter[2] ),
    .A1(net225),
    .S(_0129_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_1 _1085_ (.A(_0132_),
    .B(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _1086_ (.A(_0136_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1087_ (.A0(\wb_counter[3] ),
    .A1(net226),
    .S(_0129_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_1 _1088_ (.A(_0132_),
    .B(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _1089_ (.A(_0138_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(\wb_counter[4] ),
    .A1(net227),
    .S(_0129_),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _1091_ (.A(_0132_),
    .B(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _1092_ (.A(_0140_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1093_ (.A0(\wb_counter[5] ),
    .A1(net228),
    .S(_0129_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _1094_ (.A(_0132_),
    .B(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _1095_ (.A(_0142_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(\wb_counter[6] ),
    .A1(net229),
    .S(_0129_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _1097_ (.A(_0132_),
    .B(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _1098_ (.A(_0144_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1099_ (.A0(\wb_counter[7] ),
    .A1(net230),
    .S(_0129_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _1100_ (.A(_0132_),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _1101_ (.A(_0146_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1102_ (.A0(\wb_counter[8] ),
    .A1(net231),
    .S(_0129_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_1 _1103_ (.A(_0132_),
    .B(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _1104_ (.A(_0148_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1105_ (.A0(\wb_counter[9] ),
    .A1(net232),
    .S(_0129_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _1106_ (.A(_0132_),
    .B(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _1107_ (.A(_0150_),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_4 _1108_ (.A(_0128_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _1109_ (.A0(\wb_counter[10] ),
    .A1(net207),
    .S(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_1 _1110_ (.A(_0132_),
    .B(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _1111_ (.A(_0153_),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_2 _1112_ (.A(_0436_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1113_ (.A0(\wb_counter[11] ),
    .A1(net208),
    .S(_0151_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _1114_ (.A(_0154_),
    .B(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _1115_ (.A(_0156_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1116_ (.A0(\wb_counter[12] ),
    .A1(net209),
    .S(_0151_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _1117_ (.A(_0154_),
    .B(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _1118_ (.A(_0158_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(\wb_counter[13] ),
    .A1(net210),
    .S(_0151_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _1120_ (.A(_0154_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _1121_ (.A(_0160_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1122_ (.A0(\wb_counter[14] ),
    .A1(net211),
    .S(_0151_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _1123_ (.A(_0154_),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _1124_ (.A(_0162_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1125_ (.A0(\wb_counter[15] ),
    .A1(net212),
    .S(_0151_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _1126_ (.A(_0154_),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _1127_ (.A(_0164_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(\wb_counter[16] ),
    .A1(net213),
    .S(_0151_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_1 _1129_ (.A(_0154_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _1130_ (.A(_0166_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1131_ (.A0(\wb_counter[17] ),
    .A1(net214),
    .S(_0151_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _1132_ (.A(_0154_),
    .B(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _1133_ (.A(_0168_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1134_ (.A0(\wb_counter[18] ),
    .A1(net215),
    .S(_0151_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _1135_ (.A(_0154_),
    .B(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _1136_ (.A(_0170_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1137_ (.A0(\wb_counter[19] ),
    .A1(net216),
    .S(_0151_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _1138_ (.A(_0154_),
    .B(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _1139_ (.A(_0172_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _1140_ (.A0(\wb_counter[20] ),
    .A1(net218),
    .S(_0128_),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _1141_ (.A(_0154_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_1 _1142_ (.A(_0174_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1143_ (.A0(\wb_counter[21] ),
    .A1(net219),
    .S(_0128_),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _1144_ (.A(_0451_),
    .B(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__clkbuf_1 _1145_ (.A(_0176_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(\wb_counter[22] ),
    .A1(net220),
    .S(_0128_),
    .X(_0177_));
 sky130_fd_sc_hd__and2_1 _1147_ (.A(_0451_),
    .B(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_1 _1148_ (.A(_0178_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _1149_ (.A0(\wb_counter[23] ),
    .A1(net221),
    .S(_0128_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_1 _1150_ (.A(_0451_),
    .B(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__clkbuf_1 _1151_ (.A(_0180_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _1152_ (.A(_0451_),
    .B(wb_feedback_delay),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _1153_ (.A(_0181_),
    .X(_0084_));
 sky130_fd_sc_hd__or4b_1 _1154_ (.A(_0431_),
    .B(_0427_),
    .C(net201),
    .D_N(_0568_),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_4 _1155_ (.A(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_4 _1156_ (.A(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _1157_ (.A0(net206),
    .A1(\wb_io_override[0] ),
    .S(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_1 _1158_ (.A(_0185_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(net217),
    .A1(\wb_io_override[1] ),
    .S(_0184_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _1160_ (.A(_0186_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _1161_ (.A0(net225),
    .A1(\wb_io_override[2] ),
    .S(_0184_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _1162_ (.A(_0187_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1163_ (.A0(net226),
    .A1(\wb_io_override[3] ),
    .S(_0184_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _1164_ (.A(_0188_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1165_ (.A0(net227),
    .A1(\wb_io_override[4] ),
    .S(_0184_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _1166_ (.A(_0189_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1167_ (.A0(net228),
    .A1(\wb_io_override[5] ),
    .S(_0184_),
    .X(_0190_));
 sky130_fd_sc_hd__clkbuf_1 _1168_ (.A(_0190_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1169_ (.A0(net229),
    .A1(\wb_io_override[6] ),
    .S(_0184_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _1170_ (.A(_0191_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _1171_ (.A0(net230),
    .A1(\wb_io_override[7] ),
    .S(_0184_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _1172_ (.A(_0192_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1173_ (.A0(net231),
    .A1(\wb_io_override[8] ),
    .S(_0184_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _1174_ (.A(_0193_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(net232),
    .A1(\wb_io_override[9] ),
    .S(_0184_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _1176_ (.A(_0194_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _1177_ (.A(_0183_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(net207),
    .A1(\wb_io_override[10] ),
    .S(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _1179_ (.A(_0196_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(net208),
    .A1(\wb_io_override[11] ),
    .S(_0195_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _1181_ (.A(_0197_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(net209),
    .A1(\wb_io_override[12] ),
    .S(_0195_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _1183_ (.A(_0198_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(net210),
    .A1(\wb_io_override[13] ),
    .S(_0195_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _1185_ (.A(_0199_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _1186_ (.A0(net211),
    .A1(\wb_io_override[14] ),
    .S(_0195_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _1187_ (.A(_0200_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(net212),
    .A1(\wb_io_override[15] ),
    .S(_0195_),
    .X(_0201_));
 sky130_fd_sc_hd__clkbuf_1 _1189_ (.A(_0201_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(net213),
    .A1(\wb_io_override[16] ),
    .S(_0195_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _1191_ (.A(_0202_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1192_ (.A0(net214),
    .A1(\wb_io_override[17] ),
    .S(_0195_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _1193_ (.A(_0203_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1194_ (.A0(net215),
    .A1(\wb_io_override[18] ),
    .S(_0195_),
    .X(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _1195_ (.A(_0204_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _1196_ (.A0(net216),
    .A1(\wb_io_override[19] ),
    .S(_0195_),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _1197_ (.A(_0205_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1198_ (.A0(net218),
    .A1(\wb_io_override[20] ),
    .S(_0183_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _1199_ (.A(_0206_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(net219),
    .A1(\wb_io_override[21] ),
    .S(_0183_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _1201_ (.A(_0207_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1202_ (.A0(net220),
    .A1(\wb_io_override[22] ),
    .S(_0183_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _1203_ (.A(_0208_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _1204_ (.A0(net221),
    .A1(\wb_io_override[23] ),
    .S(_0183_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _1205_ (.A(_0209_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1206_ (.A0(net222),
    .A1(\wb_io_override[24] ),
    .S(_0183_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _1207_ (.A(_0210_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1208_ (.A0(net223),
    .A1(\wb_io_override[25] ),
    .S(_0183_),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _1209_ (.A(_0211_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(net224),
    .A1(\wb_io_override[26] ),
    .S(_0183_),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _1211_ (.A(_0212_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _1212_ (.A0(net191),
    .A1(\wb_design_addr_override[0] ),
    .S(wb_override),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(_0230_),
    .A1(_0213_),
    .S(_0451_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _1214_ (.A(_0214_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1215_ (.A0(net192),
    .A1(\wb_design_addr_override[1] ),
    .S(wb_override),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _1216_ (.A0(_0222_),
    .A1(_0215_),
    .S(_0451_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _1217_ (.A(_0216_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1218_ (.A0(net193),
    .A1(\wb_design_addr_override[2] ),
    .S(wb_override),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1219_ (.A0(_0235_),
    .A1(_0217_),
    .S(_0451_),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _1220_ (.A(_0218_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1221_ (.A0(net194),
    .A1(\wb_design_addr_override[3] ),
    .S(wb_override),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(_0234_),
    .A1(_0219_),
    .S(_0451_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _1223_ (.A(_0220_),
    .X(_0115_));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0000_),
    .Q(net328));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0001_),
    .Q(net339));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0002_),
    .Q(net347));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0003_),
    .Q(net348));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0004_),
    .Q(net349));
 sky130_fd_sc_hd__dfxtp_1 _1229_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0005_),
    .Q(net350));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0006_),
    .Q(net351));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0007_),
    .Q(net352));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0008_),
    .Q(net353));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0009_),
    .Q(net354));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0010_),
    .Q(net329));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0011_),
    .Q(net330));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0012_),
    .Q(net331));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0013_),
    .Q(net332));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0014_),
    .Q(net333));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0015_),
    .Q(net334));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0016_),
    .Q(net335));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0017_),
    .Q(net336));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0018_),
    .Q(net337));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0019_),
    .Q(net338));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0020_),
    .Q(net340));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0021_),
    .Q(net341));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_0022_),
    .Q(net342));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0023_),
    .Q(net343));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0024_),
    .Q(net344));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0025_),
    .Q(net345));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0026_),
    .Q(net346));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_1_0__leaf_net235),
    .D(net411),
    .Q(\wb_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_1_0__leaf_net235),
    .D(net409),
    .Q(\wb_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_1_0__leaf_net235),
    .D(_0029_),
    .Q(\wb_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_1_0__leaf_net235),
    .D(_0030_),
    .Q(\wb_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_1_0__leaf_net235),
    .D(net404),
    .Q(\wb_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_1_0__leaf_net235),
    .D(_0032_),
    .Q(\wb_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_1_0__leaf_net235),
    .D(net414),
    .Q(\wb_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_1_0__leaf_net235),
    .D(net407),
    .Q(\wb_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_1_0__leaf_net235),
    .D(net402),
    .Q(\wb_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_1_0__leaf_net235),
    .D(_0036_),
    .Q(\wb_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_1_1__leaf_net235),
    .D(net394),
    .Q(\wb_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_1_1__leaf_net235),
    .D(net400),
    .Q(\wb_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_1_1__leaf_net235),
    .D(net389),
    .Q(\wb_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_1_1__leaf_net235),
    .D(_0040_),
    .Q(\wb_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_1_1__leaf_net235),
    .D(_0041_),
    .Q(\wb_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_1_1__leaf_net235),
    .D(net398),
    .Q(\wb_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_1_1__leaf_net235),
    .D(_0043_),
    .Q(\wb_counter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_1_1__leaf_net235),
    .D(_0044_),
    .Q(\wb_counter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_1_1__leaf_net235),
    .D(net387),
    .Q(\wb_counter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_1_1__leaf_net235),
    .D(_0046_),
    .Q(\wb_counter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_1_1__leaf_net235),
    .D(net396),
    .Q(\wb_counter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_1_1__leaf_net235),
    .D(net391),
    .Q(\wb_counter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_1_1__leaf_net235),
    .D(_0049_),
    .Q(\wb_counter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_1_1__leaf_net235),
    .D(net385),
    .Q(\wb_counter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0051_),
    .Q(wb_rst_override));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0052_),
    .Q(wb_clk_override));
 sky130_fd_sc_hd__dfxtp_2 _1277_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0053_),
    .Q(wb_override));
 sky130_fd_sc_hd__dfxtp_1 _1278_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0054_),
    .Q(\wb_design_addr_override[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0055_),
    .Q(\wb_design_addr_override[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0056_),
    .Q(\wb_design_addr_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0057_),
    .Q(\wb_design_addr_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0058_),
    .Q(wb_single_step));
 sky130_fd_sc_hd__dfxtp_1 _1283_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0059_),
    .Q(wb_feedback_delay));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0060_),
    .Q(\wb_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0061_),
    .Q(\wb_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0062_),
    .Q(\wb_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0063_),
    .Q(\wb_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0064_),
    .Q(\wb_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_0065_),
    .Q(\wb_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0066_),
    .Q(\wb_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0067_),
    .Q(\wb_counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0068_),
    .Q(\wb_counter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0069_),
    .Q(\wb_counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0070_),
    .Q(\wb_counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1295_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0071_),
    .Q(\wb_counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0072_),
    .Q(\wb_counter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0073_),
    .Q(\wb_counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1298_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0074_),
    .Q(\wb_counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0075_),
    .Q(\wb_counter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0076_),
    .Q(\wb_counter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0077_),
    .Q(\wb_counter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0078_),
    .Q(\wb_counter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0079_),
    .Q(\wb_counter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0080_),
    .Q(\wb_counter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_0081_),
    .Q(\wb_counter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0082_),
    .Q(\wb_counter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_0083_),
    .Q(\wb_counter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_0084_),
    .Q(net327));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0085_),
    .Q(\wb_io_override[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0086_),
    .Q(\wb_io_override[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0087_),
    .Q(\wb_io_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0088_),
    .Q(\wb_io_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0089_),
    .Q(\wb_io_override[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0090_),
    .Q(\wb_io_override[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0091_),
    .Q(\wb_io_override[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0092_),
    .Q(\wb_io_override[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0093_),
    .Q(\wb_io_override[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0094_),
    .Q(\wb_io_override[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1319_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0095_),
    .Q(\wb_io_override[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0096_),
    .Q(\wb_io_override[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1321_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0097_),
    .Q(\wb_io_override[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1322_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0098_),
    .Q(\wb_io_override[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0099_),
    .Q(\wb_io_override[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0100_),
    .Q(\wb_io_override[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1325_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0101_),
    .Q(\wb_io_override[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1326_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_0102_),
    .Q(\wb_io_override[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1327_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0103_),
    .Q(\wb_io_override[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1328_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0104_),
    .Q(\wb_io_override[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1329_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0105_),
    .Q(\wb_io_override[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1330_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0106_),
    .Q(\wb_io_override[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1331_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0107_),
    .Q(\wb_io_override[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1332_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0108_),
    .Q(\wb_io_override[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1333_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0109_),
    .Q(\wb_io_override[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1334_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_0110_),
    .Q(\wb_io_override[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1335_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0111_),
    .Q(\wb_io_override[26] ));
 sky130_fd_sc_hd__dfxtp_2 _1336_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0112_),
    .Q(\design_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1337_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0113_),
    .Q(\design_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1338_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0114_),
    .Q(\design_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1339_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_0115_),
    .Q(\design_addr[3] ));
 sky130_fd_sc_hd__conb_1 multiplexer_374 (.HI(net374));
 sky130_fd_sc_hd__conb_1 multiplexer_375 (.HI(net375));
 sky130_fd_sc_hd__conb_1 multiplexer_376 (.HI(net376));
 sky130_fd_sc_hd__conb_1 multiplexer_377 (.HI(net377));
 sky130_fd_sc_hd__conb_1 multiplexer_378 (.HI(net378));
 sky130_fd_sc_hd__conb_1 multiplexer_379 (.HI(net379));
 sky130_fd_sc_hd__conb_1 multiplexer_380 (.HI(net380));
 sky130_fd_sc_hd__conb_1 multiplexer_381 (.HI(net381));
 sky130_fd_sc_hd__conb_1 multiplexer_382 (.HI(net382));
 sky130_fd_sc_hd__conb_1 multiplexer_383 (.HI(net383));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 multiplexer_358 (.LO(net358));
 sky130_fd_sc_hd__conb_1 multiplexer_359 (.LO(net359));
 sky130_fd_sc_hd__conb_1 multiplexer_360 (.LO(net360));
 sky130_fd_sc_hd__conb_1 multiplexer_361 (.LO(net361));
 sky130_fd_sc_hd__conb_1 multiplexer_362 (.LO(net362));
 sky130_fd_sc_hd__conb_1 multiplexer_363 (.LO(net363));
 sky130_fd_sc_hd__conb_1 multiplexer_364 (.LO(net364));
 sky130_fd_sc_hd__conb_1 multiplexer_365 (.LO(net365));
 sky130_fd_sc_hd__conb_1 multiplexer_366 (.LO(net366));
 sky130_fd_sc_hd__conb_1 multiplexer_367 (.LO(net367));
 sky130_fd_sc_hd__conb_1 multiplexer_368 (.LO(net368));
 sky130_fd_sc_hd__conb_1 multiplexer_369 (.LO(net369));
 sky130_fd_sc_hd__conb_1 multiplexer_370 (.LO(net370));
 sky130_fd_sc_hd__conb_1 multiplexer_371 (.LO(net371));
 sky130_fd_sc_hd__conb_1 multiplexer_372 (.LO(net372));
 sky130_fd_sc_hd__conb_1 multiplexer_373 (.HI(net373));
 sky130_fd_sc_hd__clkbuf_1 _1367_ (.A(net266),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 _1368_ (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 _1369_ (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _1370_ (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 _1371_ (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _1372_ (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 _1373_ (.A(net355),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 _1374_ (.A(net355),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 _1375_ (.A(net355),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 _1376_ (.A(net355),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 _1377_ (.A(net355),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 _1378_ (.A(net355),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 _1379_ (.A(net355),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 _1380_ (.A(net355),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 _1381_ (.A(net355),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 _1382_ (.A(net355),
    .X(net288));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(dso_6502[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(dso_6502[10]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(dso_6502[11]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(dso_6502[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(dso_6502[13]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(dso_6502[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(dso_6502[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(dso_6502[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(dso_6502[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(dso_6502[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(dso_6502[19]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(dso_6502[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(dso_6502[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(dso_6502[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(dso_6502[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(dso_6502[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(dso_6502[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(dso_6502[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(dso_6502[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(dso_6502[2]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(dso_6502[3]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(dso_6502[4]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(dso_6502[5]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(dso_6502[6]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(dso_6502[7]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(dso_6502[8]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(dso_6502[9]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(dso_LCD[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(dso_LCD[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(dso_LCD[2]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(dso_LCD[3]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(dso_LCD[4]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(dso_LCD[5]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(dso_LCD[6]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(dso_LCD[7]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(dso_as1802[0]),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(dso_as1802[10]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(dso_as1802[11]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(dso_as1802[12]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(dso_as1802[13]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(dso_as1802[14]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(dso_as1802[15]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(dso_as1802[16]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(dso_as1802[17]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(dso_as1802[18]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(dso_as1802[19]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(dso_as1802[1]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(dso_as1802[20]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(dso_as1802[21]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(dso_as1802[22]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(dso_as1802[23]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(dso_as1802[24]),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 input53 (.A(dso_as1802[25]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(dso_as1802[26]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(dso_as1802[2]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(dso_as1802[3]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(dso_as1802[4]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(dso_as1802[5]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(dso_as1802[6]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(dso_as1802[7]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(dso_as1802[8]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(dso_as1802[9]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(dso_as2650[0]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(dso_as2650[10]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(dso_as2650[11]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(dso_as2650[12]),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 input67 (.A(dso_as2650[13]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(dso_as2650[14]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(dso_as2650[15]),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 input70 (.A(dso_as2650[16]),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(dso_as2650[17]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(dso_as2650[18]),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 input73 (.A(dso_as2650[19]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(dso_as2650[1]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(dso_as2650[20]),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(dso_as2650[21]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(dso_as2650[22]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(dso_as2650[23]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(dso_as2650[24]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(dso_as2650[25]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(dso_as2650[26]),
    .X(net81));
 sky130_fd_sc_hd__dlymetal6s2s_1 input82 (.A(dso_as2650[2]),
    .X(net82));
 sky130_fd_sc_hd__dlymetal6s2s_1 input83 (.A(dso_as2650[3]),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 input84 (.A(dso_as2650[4]),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(dso_as2650[5]),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 input86 (.A(dso_as2650[6]),
    .X(net86));
 sky130_fd_sc_hd__dlymetal6s2s_1 input87 (.A(dso_as2650[7]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(dso_as2650[8]),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(dso_as2650[9]),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(dso_as5401[0]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(dso_as5401[10]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(dso_as5401[11]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(dso_as5401[12]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(dso_as5401[13]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(dso_as5401[14]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(dso_as5401[15]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(dso_as5401[16]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(dso_as5401[17]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(dso_as5401[18]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(dso_as5401[19]),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 input101 (.A(dso_as5401[1]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(dso_as5401[20]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(dso_as5401[21]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(dso_as5401[22]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(dso_as5401[23]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(dso_as5401[24]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(dso_as5401[25]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(dso_as5401[26]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(dso_as5401[2]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(dso_as5401[3]),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 input111 (.A(dso_as5401[4]),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 input112 (.A(dso_as5401[5]),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 input113 (.A(dso_as5401[6]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(dso_as5401[7]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(dso_as5401[8]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(dso_as5401[9]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(dso_counter[0]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(dso_counter[10]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(dso_counter[11]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(dso_counter[1]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(dso_counter[2]),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(dso_counter[3]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(dso_counter[4]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(dso_counter[5]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(dso_counter[6]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(dso_counter[7]),
    .X(net126));
 sky130_fd_sc_hd__buf_2 input127 (.A(dso_counter[8]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(dso_counter[9]),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 input129 (.A(dso_diceroll[0]),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(dso_diceroll[1]),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 input131 (.A(dso_diceroll[2]),
    .X(net131));
 sky130_fd_sc_hd__dlymetal6s2s_1 input132 (.A(dso_diceroll[3]),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 input133 (.A(dso_diceroll[4]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(dso_diceroll[5]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(dso_diceroll[6]),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input136 (.A(dso_diceroll[7]),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(dso_mc14500[0]),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 input138 (.A(dso_mc14500[1]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(dso_mc14500[2]),
    .X(net139));
 sky130_fd_sc_hd__dlymetal6s2s_1 input140 (.A(dso_mc14500[3]),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 input141 (.A(dso_mc14500[4]),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 input142 (.A(dso_mc14500[5]),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 input143 (.A(dso_mc14500[6]),
    .X(net143));
 sky130_fd_sc_hd__dlymetal6s2s_1 input144 (.A(dso_mc14500[7]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(dso_mc14500[8]),
    .X(net145));
 sky130_fd_sc_hd__dlymetal6s2s_1 input146 (.A(dso_multiplier[0]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(dso_multiplier[1]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(dso_multiplier[2]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(dso_multiplier[3]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(dso_multiplier[4]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(dso_multiplier[5]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(dso_multiplier[6]),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 input153 (.A(dso_multiplier[7]),
    .X(net153));
 sky130_fd_sc_hd__dlymetal6s2s_1 input154 (.A(dso_tbb1143[0]),
    .X(net154));
 sky130_fd_sc_hd__dlymetal6s2s_1 input155 (.A(dso_tbb1143[1]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 input156 (.A(dso_tbb1143[2]),
    .X(net156));
 sky130_fd_sc_hd__dlymetal6s2s_1 input157 (.A(dso_tbb1143[3]),
    .X(net157));
 sky130_fd_sc_hd__dlymetal6s2s_1 input158 (.A(dso_tbb1143[4]),
    .X(net158));
 sky130_fd_sc_hd__dlymetal6s2s_1 input159 (.A(dso_tbb1143[5]),
    .X(net159));
 sky130_fd_sc_hd__dlymetal6s2s_1 input160 (.A(dso_tbb1143[6]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(dso_tbb1143[7]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(dso_tune),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(io_in[10]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(io_in[11]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(io_in[12]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(io_in[13]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(io_in[14]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(io_in[15]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(io_in[16]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(io_in[17]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(io_in[18]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(io_in[19]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(io_in[20]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(io_in[21]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(io_in[22]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(io_in[23]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(io_in[24]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(io_in[25]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(io_in[26]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(io_in[27]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(io_in[28]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(io_in[29]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(io_in[30]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(io_in[31]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(io_in[32]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(io_in[33]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(io_in[34]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(io_in[35]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(io_in[36]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(io_in[37]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(io_in[5]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(io_in[6]),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 input193 (.A(io_in[7]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(io_in[8]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(io_in[9]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(oeb_6502),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(oeb_as1802),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(oeb_as2650),
    .X(net198));
 sky130_fd_sc_hd__dlymetal6s2s_1 input199 (.A(oeb_as5401),
    .X(net199));
 sky130_fd_sc_hd__dlymetal6s2s_1 input200 (.A(oeb_mc14500),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 input201 (.A(wb_rst_i),
    .X(net201));
 sky130_fd_sc_hd__dlymetal6s2s_1 input202 (.A(wbs_adr_i[21]),
    .X(net202));
 sky130_fd_sc_hd__buf_2 input203 (.A(wbs_adr_i[22]),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 input204 (.A(wbs_adr_i[23]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(wbs_cyc_i),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input206 (.A(wbs_dat_i[0]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(wbs_dat_i[10]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 input208 (.A(wbs_dat_i[11]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(wbs_dat_i[12]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(wbs_dat_i[13]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(wbs_dat_i[14]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(wbs_dat_i[15]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(wbs_dat_i[16]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(wbs_dat_i[17]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 input215 (.A(wbs_dat_i[18]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 input216 (.A(wbs_dat_i[19]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(wbs_dat_i[1]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 input218 (.A(wbs_dat_i[20]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 input219 (.A(wbs_dat_i[21]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input220 (.A(wbs_dat_i[22]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_2 input221 (.A(wbs_dat_i[23]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 input222 (.A(wbs_dat_i[24]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(wbs_dat_i[25]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 input224 (.A(wbs_dat_i[26]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(wbs_dat_i[2]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(wbs_dat_i[3]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(wbs_dat_i[4]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(wbs_dat_i[5]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 input229 (.A(wbs_dat_i[6]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 input230 (.A(wbs_dat_i[7]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 input231 (.A(wbs_dat_i[8]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 input232 (.A(wbs_dat_i[9]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(wbs_stb_i),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(wbs_we_i),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(clknet_1_1__leaf_net235),
    .X(design_clk_o));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(dsi_all[0]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(dsi_all[10]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(dsi_all[11]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(dsi_all[12]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(dsi_all[13]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(dsi_all[14]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(dsi_all[15]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(dsi_all[16]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(dsi_all[17]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(dsi_all[18]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(dsi_all[19]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(dsi_all[1]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(dsi_all[20]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(dsi_all[21]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(dsi_all[22]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(dsi_all[23]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(dsi_all[24]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(dsi_all[25]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(dsi_all[26]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(dsi_all[2]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(dsi_all[3]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(dsi_all[4]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(dsi_all[5]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net259),
    .X(dsi_all[6]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net260),
    .X(dsi_all[7]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .X(dsi_all[8]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .X(dsi_all[9]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .X(io_oeb[11]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(io_oeb[12]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(io_oeb[13]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(io_oeb[14]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(io_oeb[15]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(io_oeb[16]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(io_oeb[17]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(io_oeb[18]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(io_oeb[19]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(io_oeb[20]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(io_oeb[21]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(io_oeb[22]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(io_oeb[23]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(io_oeb[24]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(io_oeb[25]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(io_oeb[26]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(io_oeb[27]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(io_oeb[28]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(io_oeb[29]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(io_oeb[30]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(io_oeb[31]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(io_oeb[32]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(io_oeb[33]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(io_oeb[34]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(io_oeb[35]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(io_oeb[36]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(io_oeb[37]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net299),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net303),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net304),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(io_out[35]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(rst_6502));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .X(rst_LCD));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .X(rst_as1802));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .X(rst_as2650));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(rst_as5401));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(rst_counter));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(rst_diceroll));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(rst_mc14500));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(rst_tbb1143));
 sky130_fd_sc_hd__buf_2 output326 (.A(net326),
    .X(rst_tune));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net348),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output351 (.A(net351),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 fanout356 (.A(net289),
    .X(net356));
 sky130_fd_sc_hd__conb_1 multiplexer_357 (.LO(net357));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_net235 (.A(net235),
    .X(clknet_0_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_net235 (.A(clknet_0_net235),
    .X(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_net235 (.A(clknet_0_net235),
    .X(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\wb_counter[23] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0050_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\wb_counter[18] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0045_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\wb_counter[12] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0039_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\wb_counter[21] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0048_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\wb_counter[10] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0547_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0037_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\wb_counter[20] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0047_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\wb_counter[15] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0042_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\wb_counter[11] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0038_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\wb_counter[8] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0035_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\wb_counter[4] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0031_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\wb_counter[7] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0541_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0034_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\wb_counter[1] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0028_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\wb_counter[0] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0027_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\wb_counter[6] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0458_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0033_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\wb_counter[17] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0558_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0560_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\wb_counter[22] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0566_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0567_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\wb_counter[13] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0550_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\wb_counter[16] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0556_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0557_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\wb_counter[19] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0562_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0563_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\wb_counter[14] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\wb_counter[3] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0532_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0534_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\wb_counter[9] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0544_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0545_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\wb_counter[5] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0537_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\wb_counter[2] ),
    .X(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__S (.DIODE(_0129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__B (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__B (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__C (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A2 (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__A (.DIODE(_0226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A2 (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__A (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__A2 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__B_N (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__A (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A2 (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__A (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__B_N (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__B1 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__B1 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__B_N (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__B1 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__B1 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B1 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A2 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A2 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A2 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__A2 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__A2 (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0644__A (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__B_N (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A2 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__A2 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__A2 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A2 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__B1 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__A2 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A2 (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__A (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__A (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__B_N (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__A2 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A2 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__A2 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A2 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__B1 (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__A (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A2 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A2 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__A2 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__A2 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__A2 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__A2 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__B1 (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__B_N (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__A2 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__B1 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__A2 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A2 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__A2 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__A2 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__B1 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__A2 (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__A (.DIODE(_0258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__B1 (.DIODE(_0258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__A1 (.DIODE(_0259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__B1 (.DIODE(_0259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A2 (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A2 (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__C (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A2 (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__A (.DIODE(_0264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__B1 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__B1 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__B (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__A2 (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__B1 (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__A (.DIODE(_0270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A2 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__B1 (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__A (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__A2 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__A2 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__B1 (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__B (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__B1 (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__B (.DIODE(_0277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__C1 (.DIODE(_0308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__C1 (.DIODE(_0355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__C1 (.DIODE(_0361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__C1 (.DIODE(_0367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__C1 (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A1 (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__A_N (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A_N (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A_N (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__A_N (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__A_N (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__A_N (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__A (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__S (.DIODE(_0386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0958__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__B (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__S (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__B (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__A1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A1 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__S (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__S (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__S (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__S (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__B1 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__A2 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__A2 (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__A (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A_N (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__D_N (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__C (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(dso_6502[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(dso_6502[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(dso_6502[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(dso_6502[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(dso_6502[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(dso_6502[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(dso_6502[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(dso_6502[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(dso_6502[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(dso_6502[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(dso_6502[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(dso_6502[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(dso_6502[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(dso_6502[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(dso_6502[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(dso_6502[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(dso_6502[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(dso_6502[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(dso_6502[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(dso_6502[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(dso_6502[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(dso_6502[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(dso_6502[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(dso_6502[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(dso_6502[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(dso_6502[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(dso_6502[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(dso_LCD[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(dso_LCD[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(dso_LCD[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(dso_LCD[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(dso_LCD[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(dso_LCD[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(dso_LCD[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(dso_LCD[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(dso_as1802[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(dso_as1802[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(dso_as1802[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(dso_as1802[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(dso_as1802[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(dso_as1802[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(dso_as1802[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(dso_as1802[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(dso_as1802[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(dso_as1802[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(dso_as1802[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(dso_as1802[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(dso_as1802[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(dso_as1802[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(dso_as1802[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(dso_as1802[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(dso_as1802[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(dso_as1802[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(dso_as1802[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(dso_as1802[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(dso_as1802[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(dso_as1802[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(dso_as1802[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(dso_as1802[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(dso_as1802[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(dso_as1802[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(dso_as1802[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(dso_as2650[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(dso_as2650[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(dso_as2650[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(dso_as2650[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(dso_as2650[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(dso_as2650[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(dso_as2650[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(dso_as2650[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(dso_as2650[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(dso_as2650[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(dso_as2650[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(dso_as2650[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(dso_as2650[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(dso_as2650[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(dso_as2650[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(dso_as2650[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(dso_as2650[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(dso_as2650[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(dso_as2650[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(dso_as2650[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(dso_as2650[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(dso_as2650[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(dso_as2650[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(dso_as2650[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(dso_as2650[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(dso_as2650[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(dso_as2650[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(dso_as5401[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(dso_as5401[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(dso_as5401[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(dso_as5401[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(dso_as5401[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(dso_as5401[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(dso_as5401[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(dso_as5401[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(dso_as5401[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(dso_as5401[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(dso_as5401[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(dso_as5401[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(dso_as5401[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(dso_as5401[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(dso_as5401[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(dso_as5401[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(dso_as5401[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(dso_as5401[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(dso_as5401[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(dso_as5401[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(dso_as5401[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(dso_as5401[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(dso_as5401[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(dso_as5401[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(dso_as5401[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(dso_as5401[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(dso_as5401[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(dso_counter[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(dso_counter[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(dso_counter[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(dso_counter[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(dso_counter[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(dso_counter[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(dso_counter[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(dso_counter[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(dso_counter[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(dso_counter[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(dso_counter[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(dso_counter[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(dso_diceroll[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(dso_diceroll[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(dso_diceroll[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(dso_diceroll[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(dso_diceroll[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(dso_diceroll[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(dso_diceroll[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(dso_diceroll[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(dso_mc14500[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(dso_mc14500[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(dso_mc14500[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(dso_mc14500[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(dso_mc14500[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(dso_mc14500[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(dso_mc14500[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(dso_mc14500[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(dso_mc14500[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(dso_multiplier[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(dso_multiplier[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(dso_multiplier[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(dso_multiplier[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(dso_multiplier[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(dso_multiplier[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(dso_multiplier[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(dso_multiplier[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(dso_tbb1143[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(dso_tbb1143[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(dso_tbb1143[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(dso_tbb1143[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(dso_tbb1143[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(dso_tbb1143[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(dso_tbb1143[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(dso_tbb1143[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(dso_tune));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(io_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(io_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(io_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(io_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(io_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(io_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(io_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(io_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(io_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(io_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(oeb_6502));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(oeb_as1802));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(oeb_as2650));
 sky130_fd_sc_hd__diode_2 ANTENNA_input199_A (.DIODE(oeb_as5401));
 sky130_fd_sc_hd__diode_2 ANTENNA_input200_A (.DIODE(oeb_mc14500));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A1 (.DIODE(\wb_io_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A2 (.DIODE(\wb_io_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input201_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input202_A (.DIODE(wbs_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input203_A (.DIODE(wbs_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input204_A (.DIODE(wbs_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input205_A (.DIODE(wbs_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input206_A (.DIODE(wbs_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input207_A (.DIODE(wbs_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input208_A (.DIODE(wbs_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input209_A (.DIODE(wbs_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input210_A (.DIODE(wbs_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input211_A (.DIODE(wbs_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input212_A (.DIODE(wbs_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input213_A (.DIODE(wbs_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input214_A (.DIODE(wbs_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input215_A (.DIODE(wbs_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input216_A (.DIODE(wbs_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input217_A (.DIODE(wbs_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input218_A (.DIODE(wbs_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input219_A (.DIODE(wbs_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input220_A (.DIODE(wbs_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input221_A (.DIODE(wbs_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input222_A (.DIODE(wbs_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input223_A (.DIODE(wbs_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input224_A (.DIODE(wbs_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input225_A (.DIODE(wbs_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input226_A (.DIODE(wbs_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input227_A (.DIODE(wbs_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input228_A (.DIODE(wbs_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input229_A (.DIODE(wbs_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input230_A (.DIODE(wbs_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input231_A (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input232_A (.DIODE(wbs_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input233_A (.DIODE(wbs_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input234_A (.DIODE(wbs_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__B2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__B2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__A_N (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__B_N (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__A0 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__A0 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__A0 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__A0 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__A0 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__A0 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__A0 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__A0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__A0 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__A0 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__A0 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__A1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A0 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__A0 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__A0 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__A0 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A0 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A0 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__A0 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__A0 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__A0 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__A0 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__A0 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__A3 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A3 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_output267_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__A3 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__A3 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__A3 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__A3 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__B1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_output272_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__A3 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A3 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_output274_A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__A3 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__A3 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__0644__B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__A3 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__A3 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_output278_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__A3 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A3 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A3 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__D (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A3 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__B1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A1_N (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__B1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__B1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_output300_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__A3 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_output301_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A3 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__A2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output306_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_output309_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_output310_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_output311_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_output313_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_output314_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__B2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_output315_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__B2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_output316_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__B2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_output317_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_output319_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_output320_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_output322_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_output323_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_output324_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_output326_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_output331_A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__B2 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_output339_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_output341_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__A1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_output342_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__A1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_output343_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__A1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_output344_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_output345_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_output346_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A3 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1229__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__CLK (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__CLK (.DIODE(clknet_1_0__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1274__CLK (.DIODE(clknet_1_1__leaf_net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_output235_A (.DIODE(clknet_1_1__leaf_net235));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_580 ();
 assign io_oeb[0] = net373;
 assign io_oeb[10] = net383;
 assign io_oeb[1] = net374;
 assign io_oeb[2] = net375;
 assign io_oeb[3] = net376;
 assign io_oeb[4] = net377;
 assign io_oeb[5] = net378;
 assign io_oeb[6] = net379;
 assign io_oeb[7] = net380;
 assign io_oeb[8] = net381;
 assign io_oeb[9] = net382;
 assign io_out[0] = net357;
 assign io_out[10] = net367;
 assign io_out[1] = net358;
 assign io_out[2] = net359;
 assign io_out[3] = net360;
 assign io_out[4] = net361;
 assign io_out[5] = net362;
 assign io_out[6] = net363;
 assign io_out[7] = net364;
 assign io_out[8] = net365;
 assign io_out[9] = net366;
 assign wbs_dat_o[27] = net368;
 assign wbs_dat_o[28] = net369;
 assign wbs_dat_o[29] = net370;
 assign wbs_dat_o[30] = net371;
 assign wbs_dat_o[31] = net372;
endmodule

