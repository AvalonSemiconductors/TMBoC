// This is the unpowered netlist.
module tt2_tholin_namebadge (clk,
    rst,
    io_in,
    io_oeb,
    io_out);
 input clk;
 input rst;
 input [2:0] io_in;
 output [26:0] io_oeb;
 output [7:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire net49;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net50;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire clknet_0_clk;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire \lcd.num_state[0] ;
 wire \lcd.num_state[1] ;
 wire \lcd.rom_addr[0] ;
 wire \lcd.rom_addr[1] ;
 wire \lcd.rom_addr[3] ;
 wire \lcd.rom_addr[4] ;
 wire \lcd.rom_addr[5] ;
 wire \lcd.rom_addr[6] ;
 wire \lcd.round[0] ;
 wire \lcd.round[1] ;
 wire \lcd.s_ROM[0] ;
 wire \lcd.s_ROM[1] ;
 wire \lcd.s_ROM[2] ;
 wire \lcd.s_ROM[3] ;
 wire \lcd.s_ROM[4] ;
 wire \lcd.s_ROM[5] ;
 wire \lcd.s_ROM[6] ;
 wire \lcd.seq[0] ;
 wire \lcd.seq[1] ;
 wire \lcd.seq[2] ;
 wire \lcd.seq[3] ;
 wire \lcd.seq[4] ;
 wire \lcd.seq[5] ;
 wire \lcd.seq[6] ;
 wire \lcd.seq[7] ;
 wire \lcd.toggle ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_6 _369_ (.A(\lcd.toggle ),
    .Y(_340_));
 sky130_fd_sc_hd__inv_2 _370_ (.A(net36),
    .Y(_341_));
 sky130_fd_sc_hd__inv_2 _371_ (.A(net33),
    .Y(_342_));
 sky130_fd_sc_hd__inv_2 _372_ (.A(net45),
    .Y(_343_));
 sky130_fd_sc_hd__inv_2 _373_ (.A(\lcd.rom_addr[0] ),
    .Y(_344_));
 sky130_fd_sc_hd__inv_2 _374_ (.A(\lcd.rom_addr[1] ),
    .Y(_345_));
 sky130_fd_sc_hd__clkinv_2 _375_ (.A(net11),
    .Y(_346_));
 sky130_fd_sc_hd__nor2_8 _376_ (.A(\lcd.toggle ),
    .B(net4),
    .Y(_007_));
 sky130_fd_sc_hd__or2_4 _377_ (.A(net38),
    .B(net40),
    .X(_347_));
 sky130_fd_sc_hd__nor2_2 _378_ (.A(net31),
    .B(net34),
    .Y(_348_));
 sky130_fd_sc_hd__or2_4 _379_ (.A(net30),
    .B(net33),
    .X(_349_));
 sky130_fd_sc_hd__a211o_1 _380_ (.A1(net41),
    .A2(net43),
    .B1(net38),
    .C1(net40),
    .X(_350_));
 sky130_fd_sc_hd__and3b_4 _381_ (.A_N(_350_),
    .B(_341_),
    .C(_348_),
    .X(_351_));
 sky130_fd_sc_hd__or3_4 _382_ (.A(net35),
    .B(_349_),
    .C(_350_),
    .X(_352_));
 sky130_fd_sc_hd__or2_1 _383_ (.A(net40),
    .B(net41),
    .X(_353_));
 sky130_fd_sc_hd__nor3_1 _384_ (.A(net37),
    .B(net42),
    .C(_347_),
    .Y(_354_));
 sky130_fd_sc_hd__or4_1 _385_ (.A(net37),
    .B(net39),
    .C(\lcd.seq[3] ),
    .D(net42),
    .X(_355_));
 sky130_fd_sc_hd__and2_4 _386_ (.A(net31),
    .B(net34),
    .X(_356_));
 sky130_fd_sc_hd__and2b_4 _387_ (.A_N(\lcd.round[0] ),
    .B(\lcd.round[1] ),
    .X(_357_));
 sky130_fd_sc_hd__nand2b_4 _388_ (.A_N(\lcd.round[0] ),
    .B(\lcd.round[1] ),
    .Y(_358_));
 sky130_fd_sc_hd__nor2_2 _389_ (.A(net44),
    .B(net46),
    .Y(_359_));
 sky130_fd_sc_hd__nand4b_4 _390_ (.A_N(_355_),
    .B(_356_),
    .C(_357_),
    .D(_359_),
    .Y(_360_));
 sky130_fd_sc_hd__nor3_4 _391_ (.A(_340_),
    .B(_351_),
    .C(_360_),
    .Y(_361_));
 sky130_fd_sc_hd__nor2_4 _392_ (.A(_007_),
    .B(_361_),
    .Y(_362_));
 sky130_fd_sc_hd__or2_2 _393_ (.A(_007_),
    .B(_361_),
    .X(_363_));
 sky130_fd_sc_hd__nand2b_2 _394_ (.A_N(net43),
    .B(net38),
    .Y(_364_));
 sky130_fd_sc_hd__nand2_2 _395_ (.A(net40),
    .B(net41),
    .Y(_365_));
 sky130_fd_sc_hd__nand2b_1 _396_ (.A_N(net38),
    .B(net43),
    .Y(_366_));
 sky130_fd_sc_hd__or3b_1 _397_ (.A(net31),
    .B(net34),
    .C_N(net35),
    .X(_367_));
 sky130_fd_sc_hd__a221o_4 _398_ (.A1(_364_),
    .A2(_365_),
    .B1(_366_),
    .B2(_353_),
    .C1(_367_),
    .X(_368_));
 sky130_fd_sc_hd__and2_1 _399_ (.A(_357_),
    .B(_368_),
    .X(_033_));
 sky130_fd_sc_hd__and3_4 _400_ (.A(net39),
    .B(net40),
    .C(net41),
    .X(_034_));
 sky130_fd_sc_hd__nand3b_1 _401_ (.A_N(net33),
    .B(net35),
    .C(net30),
    .Y(_035_));
 sky130_fd_sc_hd__o21a_1 _402_ (.A1(net35),
    .A2(net33),
    .B1(net30),
    .X(_036_));
 sky130_fd_sc_hd__or3b_4 _403_ (.A(net36),
    .B(net34),
    .C_N(net32),
    .X(_037_));
 sky130_fd_sc_hd__and4_4 _404_ (.A(net30),
    .B(_341_),
    .C(_342_),
    .D(_034_),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _405_ (.A(_034_),
    .B(_037_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_2 _406_ (.A0(_368_),
    .A1(_039_),
    .S(_358_),
    .X(_040_));
 sky130_fd_sc_hd__and2_4 _407_ (.A(net35),
    .B(net33),
    .X(_041_));
 sky130_fd_sc_hd__o21ai_1 _408_ (.A1(net36),
    .A2(_034_),
    .B1(net34),
    .Y(_042_));
 sky130_fd_sc_hd__a211oi_4 _409_ (.A1(net33),
    .A2(_034_),
    .B1(_041_),
    .C1(net31),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _410_ (.A(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__and2b_4 _411_ (.A_N(\lcd.round[1] ),
    .B(\lcd.round[0] ),
    .X(_045_));
 sky130_fd_sc_hd__nand2b_4 _412_ (.A_N(\lcd.round[1] ),
    .B(\lcd.round[0] ),
    .Y(_046_));
 sky130_fd_sc_hd__xor2_4 _413_ (.A(\lcd.round[0] ),
    .B(\lcd.round[1] ),
    .X(_047_));
 sky130_fd_sc_hd__nor2_1 _414_ (.A(net41),
    .B(net43),
    .Y(_048_));
 sky130_fd_sc_hd__or3_2 _415_ (.A(net38),
    .B(net41),
    .C(net43),
    .X(_049_));
 sky130_fd_sc_hd__o21ai_1 _416_ (.A1(net39),
    .A2(net40),
    .B1(net36),
    .Y(_050_));
 sky130_fd_sc_hd__and3_4 _417_ (.A(net36),
    .B(_347_),
    .C(_049_),
    .X(_051_));
 sky130_fd_sc_hd__or4b_1 _418_ (.A(_349_),
    .B(_047_),
    .C(_050_),
    .D_N(_049_),
    .X(_052_));
 sky130_fd_sc_hd__o211a_4 _419_ (.A1(_043_),
    .A2(_047_),
    .B1(_052_),
    .C1(_352_),
    .X(_053_));
 sky130_fd_sc_hd__a211o_4 _420_ (.A1(net36),
    .A2(net38),
    .B1(net33),
    .C1(net30),
    .X(_054_));
 sky130_fd_sc_hd__a31o_4 _421_ (.A1(net35),
    .A2(net40),
    .A3(net41),
    .B1(_054_),
    .X(_055_));
 sky130_fd_sc_hd__o221a_4 _422_ (.A1(_356_),
    .A2(_034_),
    .B1(_035_),
    .B2(_364_),
    .C1(_036_),
    .X(_056_));
 sky130_fd_sc_hd__a21oi_4 _423_ (.A1(_347_),
    .A2(_041_),
    .B1(net32),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_1 _424_ (.A(_038_),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__o311a_1 _425_ (.A1(net38),
    .A2(net40),
    .A3(net41),
    .B1(net33),
    .C1(net35),
    .X(_059_));
 sky130_fd_sc_hd__and4bb_2 _426_ (.A_N(_347_),
    .B_N(net30),
    .C(net41),
    .D(_041_),
    .X(_060_));
 sky130_fd_sc_hd__o311ai_4 _427_ (.A1(_038_),
    .A2(_056_),
    .A3(_060_),
    .B1(_045_),
    .C1(_055_),
    .Y(_061_));
 sky130_fd_sc_hd__nor3_4 _428_ (.A(net35),
    .B(net38),
    .C(_349_),
    .Y(_062_));
 sky130_fd_sc_hd__or4_2 _429_ (.A(net30),
    .B(net35),
    .C(net33),
    .D(net38),
    .X(_063_));
 sky130_fd_sc_hd__nand2_1 _430_ (.A(_045_),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__nor2_1 _431_ (.A(net30),
    .B(_059_),
    .Y(_065_));
 sky130_fd_sc_hd__o31a_2 _432_ (.A1(net35),
    .A2(net38),
    .A3(net40),
    .B1(net33),
    .X(_066_));
 sky130_fd_sc_hd__nor2_1 _433_ (.A(net32),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__or3b_4 _434_ (.A(net30),
    .B(_059_),
    .C_N(_066_),
    .X(_068_));
 sky130_fd_sc_hd__or2_1 _435_ (.A(_357_),
    .B(_054_),
    .X(_069_));
 sky130_fd_sc_hd__a21o_2 _436_ (.A1(_068_),
    .A2(_069_),
    .B1(_064_),
    .X(_070_));
 sky130_fd_sc_hd__a41oi_4 _437_ (.A1(_040_),
    .A2(_053_),
    .A3(_061_),
    .A4(_070_),
    .B1(_340_),
    .Y(_071_));
 sky130_fd_sc_hd__a41o_4 _438_ (.A1(_040_),
    .A2(_053_),
    .A3(_061_),
    .A4(_070_),
    .B1(_340_),
    .X(_072_));
 sky130_fd_sc_hd__nor2_1 _439_ (.A(_038_),
    .B(_056_),
    .Y(_073_));
 sky130_fd_sc_hd__nor2_1 _440_ (.A(_343_),
    .B(\lcd.rom_addr[0] ),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_2 _441_ (.A(net45),
    .B(_344_),
    .Y(_075_));
 sky130_fd_sc_hd__and3_1 _442_ (.A(_362_),
    .B(_072_),
    .C(_074_),
    .X(_076_));
 sky130_fd_sc_hd__or3_1 _443_ (.A(net29),
    .B(_071_),
    .C(_075_),
    .X(_077_));
 sky130_fd_sc_hd__nor2_2 _444_ (.A(\lcd.rom_addr[1] ),
    .B(_075_),
    .Y(_078_));
 sky130_fd_sc_hd__and3_1 _445_ (.A(_362_),
    .B(_072_),
    .C(_078_),
    .X(_079_));
 sky130_fd_sc_hd__or4b_4 _446_ (.A(net11),
    .B(net29),
    .C(_071_),
    .D_N(_078_),
    .X(_080_));
 sky130_fd_sc_hd__nor3_2 _447_ (.A(\lcd.rom_addr[3] ),
    .B(\lcd.rom_addr[4] ),
    .C(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__a31o_2 _448_ (.A1(_347_),
    .A2(_041_),
    .A3(_049_),
    .B1(net31),
    .X(_082_));
 sky130_fd_sc_hd__a21oi_2 _449_ (.A1(net34),
    .A2(_051_),
    .B1(net32),
    .Y(_083_));
 sky130_fd_sc_hd__a21oi_1 _450_ (.A1(_357_),
    .A2(_082_),
    .B1(_340_),
    .Y(_084_));
 sky130_fd_sc_hd__a21o_2 _451_ (.A1(_357_),
    .A2(_082_),
    .B1(_340_),
    .X(_085_));
 sky130_fd_sc_hd__and3_4 _452_ (.A(_362_),
    .B(_072_),
    .C(_085_),
    .X(_086_));
 sky130_fd_sc_hd__or3_4 _453_ (.A(net29),
    .B(_071_),
    .C(_084_),
    .X(_087_));
 sky130_fd_sc_hd__o21a_1 _454_ (.A1(\lcd.rom_addr[3] ),
    .A2(_080_),
    .B1(\lcd.rom_addr[4] ),
    .X(_088_));
 sky130_fd_sc_hd__nor3_4 _455_ (.A(_081_),
    .B(net28),
    .C(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__clkinv_2 _456_ (.A(_089_),
    .Y(_020_));
 sky130_fd_sc_hd__o31a_4 _457_ (.A1(_343_),
    .A2(net29),
    .A3(_071_),
    .B1(\lcd.rom_addr[0] ),
    .X(_090_));
 sky130_fd_sc_hd__a31o_2 _458_ (.A1(net45),
    .A2(_362_),
    .A3(_072_),
    .B1(_344_),
    .X(_091_));
 sky130_fd_sc_hd__a211o_1 _459_ (.A1(_075_),
    .A2(_084_),
    .B1(net29),
    .C1(_071_),
    .X(_092_));
 sky130_fd_sc_hd__o211a_4 _460_ (.A1(_074_),
    .A2(_085_),
    .B1(_362_),
    .C1(_072_),
    .X(_093_));
 sky130_fd_sc_hd__nor2_4 _461_ (.A(_090_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__clkinv_4 _462_ (.A(_094_),
    .Y(_016_));
 sky130_fd_sc_hd__o31a_4 _463_ (.A1(_363_),
    .A2(_071_),
    .A3(_075_),
    .B1(\lcd.rom_addr[1] ),
    .X(_095_));
 sky130_fd_sc_hd__o211a_4 _464_ (.A1(_078_),
    .A2(_085_),
    .B1(_362_),
    .C1(_072_),
    .X(_096_));
 sky130_fd_sc_hd__nor2_8 _465_ (.A(_095_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _466_ (.A(_097_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_2 _467_ (.A(_345_),
    .B(_016_),
    .Y(_098_));
 sky130_fd_sc_hd__or3_4 _468_ (.A(_345_),
    .B(_090_),
    .C(_093_),
    .X(_099_));
 sky130_fd_sc_hd__a2111o_4 _469_ (.A1(_077_),
    .A2(_091_),
    .B1(_095_),
    .C1(_079_),
    .D1(_086_),
    .X(_100_));
 sky130_fd_sc_hd__and3_2 _470_ (.A(_345_),
    .B(_091_),
    .C(_092_),
    .X(_101_));
 sky130_fd_sc_hd__or3_4 _471_ (.A(\lcd.rom_addr[1] ),
    .B(_090_),
    .C(_093_),
    .X(_102_));
 sky130_fd_sc_hd__o22a_4 _472_ (.A1(_090_),
    .A2(_093_),
    .B1(_095_),
    .B2(_096_),
    .X(_103_));
 sky130_fd_sc_hd__a2bb2o_4 _473_ (.A1_N(_096_),
    .A2_N(_095_),
    .B1(_092_),
    .B2(_091_),
    .X(_104_));
 sky130_fd_sc_hd__nor2_2 _474_ (.A(_101_),
    .B(_103_),
    .Y(_105_));
 sky130_fd_sc_hd__a31o_2 _475_ (.A1(_362_),
    .A2(_072_),
    .A3(_078_),
    .B1(_346_),
    .X(_106_));
 sky130_fd_sc_hd__a21o_4 _476_ (.A1(_080_),
    .A2(_106_),
    .B1(net28),
    .X(_107_));
 sky130_fd_sc_hd__inv_2 _477_ (.A(_107_),
    .Y(_018_));
 sky130_fd_sc_hd__xor2_4 _478_ (.A(\lcd.rom_addr[3] ),
    .B(_080_),
    .X(_108_));
 sky130_fd_sc_hd__xnor2_4 _479_ (.A(\lcd.rom_addr[3] ),
    .B(_080_),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _480_ (.A(net28),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _481_ (.A(net23),
    .Y(_019_));
 sky130_fd_sc_hd__a31o_4 _482_ (.A1(\lcd.rom_addr[3] ),
    .A2(_080_),
    .A3(_106_),
    .B1(net28),
    .X(_111_));
 sky130_fd_sc_hd__a21oi_1 _483_ (.A1(_105_),
    .A2(_111_),
    .B1(net26),
    .Y(_112_));
 sky130_fd_sc_hd__nor2_1 _484_ (.A(_016_),
    .B(_107_),
    .Y(_113_));
 sky130_fd_sc_hd__or4_4 _485_ (.A(_346_),
    .B(_076_),
    .C(_086_),
    .D(_090_),
    .X(_114_));
 sky130_fd_sc_hd__or2_4 _486_ (.A(\lcd.rom_addr[1] ),
    .B(_114_),
    .X(_115_));
 sky130_fd_sc_hd__nand2_2 _487_ (.A(_102_),
    .B(_107_),
    .Y(_116_));
 sky130_fd_sc_hd__o211ai_1 _488_ (.A1(net17),
    .A2(_116_),
    .B1(_115_),
    .C1(_112_),
    .Y(_117_));
 sky130_fd_sc_hd__or4_2 _489_ (.A(\lcd.rom_addr[3] ),
    .B(\lcd.rom_addr[4] ),
    .C(\lcd.rom_addr[5] ),
    .D(_080_),
    .X(_118_));
 sky130_fd_sc_hd__nand2b_1 _490_ (.A_N(_081_),
    .B(\lcd.rom_addr[5] ),
    .Y(_119_));
 sky130_fd_sc_hd__and3_2 _491_ (.A(_087_),
    .B(_118_),
    .C(_119_),
    .X(_120_));
 sky130_fd_sc_hd__inv_2 _492_ (.A(net15),
    .Y(_021_));
 sky130_fd_sc_hd__or4_4 _493_ (.A(net11),
    .B(_076_),
    .C(_086_),
    .D(_090_),
    .X(_121_));
 sky130_fd_sc_hd__or2_4 _494_ (.A(net11),
    .B(_099_),
    .X(_122_));
 sky130_fd_sc_hd__or3_4 _495_ (.A(_346_),
    .B(_095_),
    .C(_096_),
    .X(_123_));
 sky130_fd_sc_hd__a31o_1 _496_ (.A1(net23),
    .A2(_122_),
    .A3(_123_),
    .B1(net20),
    .X(_124_));
 sky130_fd_sc_hd__o22a_4 _497_ (.A1(_097_),
    .A2(net25),
    .B1(_109_),
    .B2(net28),
    .X(_125_));
 sky130_fd_sc_hd__nand2_2 _498_ (.A(_099_),
    .B(net25),
    .Y(_126_));
 sky130_fd_sc_hd__a21o_1 _499_ (.A1(_102_),
    .A2(_104_),
    .B1(_107_),
    .X(_127_));
 sky130_fd_sc_hd__a21o_1 _500_ (.A1(_105_),
    .A2(_125_),
    .B1(_124_),
    .X(_128_));
 sky130_fd_sc_hd__nor2_1 _501_ (.A(\lcd.rom_addr[6] ),
    .B(_118_),
    .Y(_129_));
 sky130_fd_sc_hd__a211o_4 _502_ (.A1(\lcd.rom_addr[6] ),
    .A2(_118_),
    .B1(_129_),
    .C1(net28),
    .X(_022_));
 sky130_fd_sc_hd__inv_2 _503_ (.A(_022_),
    .Y(_130_));
 sky130_fd_sc_hd__o311a_2 _504_ (.A1(_101_),
    .A2(_103_),
    .A3(net24),
    .B1(_108_),
    .C1(_087_),
    .X(_131_));
 sky130_fd_sc_hd__a21o_1 _505_ (.A1(_126_),
    .A2(_131_),
    .B1(net20),
    .X(_132_));
 sky130_fd_sc_hd__o211a_1 _506_ (.A1(net28),
    .A2(_109_),
    .B1(_114_),
    .C1(_102_),
    .X(_133_));
 sky130_fd_sc_hd__a211o_1 _507_ (.A1(_126_),
    .A2(_131_),
    .B1(_133_),
    .C1(net20),
    .X(_134_));
 sky130_fd_sc_hd__nor2_1 _508_ (.A(net23),
    .B(_122_),
    .Y(_135_));
 sky130_fd_sc_hd__nor2_1 _509_ (.A(_103_),
    .B(net17),
    .Y(_136_));
 sky130_fd_sc_hd__and4_1 _510_ (.A(_104_),
    .B(net22),
    .C(_121_),
    .D(_123_),
    .X(_137_));
 sky130_fd_sc_hd__o311a_1 _511_ (.A1(net27),
    .A2(_135_),
    .A3(_137_),
    .B1(net14),
    .C1(_134_),
    .X(_138_));
 sky130_fd_sc_hd__a31o_1 _512_ (.A1(_117_),
    .A2(_021_),
    .A3(_128_),
    .B1(_138_),
    .X(_139_));
 sky130_fd_sc_hd__a221o_1 _513_ (.A1(_121_),
    .A2(_125_),
    .B1(_136_),
    .B2(_116_),
    .C1(net26),
    .X(_140_));
 sky130_fd_sc_hd__and4_2 _514_ (.A(_087_),
    .B(_016_),
    .C(_108_),
    .D(_123_),
    .X(_141_));
 sky130_fd_sc_hd__o21a_4 _515_ (.A1(net28),
    .A2(_109_),
    .B1(_123_),
    .X(_142_));
 sky130_fd_sc_hd__a211o_1 _516_ (.A1(_104_),
    .A2(_142_),
    .B1(_141_),
    .C1(net19),
    .X(_143_));
 sky130_fd_sc_hd__and2_1 _517_ (.A(net13),
    .B(_143_),
    .X(_144_));
 sky130_fd_sc_hd__nor2_2 _518_ (.A(_100_),
    .B(net24),
    .Y(_145_));
 sky130_fd_sc_hd__and2_2 _519_ (.A(_100_),
    .B(net24),
    .X(_146_));
 sky130_fd_sc_hd__nand2_2 _520_ (.A(_100_),
    .B(net24),
    .Y(_147_));
 sky130_fd_sc_hd__o211a_1 _521_ (.A1(_145_),
    .A2(_146_),
    .B1(_099_),
    .C1(_109_),
    .X(_148_));
 sky130_fd_sc_hd__a21o_1 _522_ (.A1(_127_),
    .A2(_131_),
    .B1(net20),
    .X(_149_));
 sky130_fd_sc_hd__and2_1 _523_ (.A(_099_),
    .B(_107_),
    .X(_150_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_099_),
    .B(_107_),
    .Y(_151_));
 sky130_fd_sc_hd__o211a_1 _525_ (.A1(_104_),
    .A2(net24),
    .B1(net22),
    .C1(_102_),
    .X(_152_));
 sky130_fd_sc_hd__a31o_1 _526_ (.A1(net16),
    .A2(_121_),
    .A3(_147_),
    .B1(net27),
    .X(_153_));
 sky130_fd_sc_hd__o22a_1 _527_ (.A1(_148_),
    .A2(_149_),
    .B1(_152_),
    .B2(_153_),
    .X(_154_));
 sky130_fd_sc_hd__a22o_1 _528_ (.A1(_140_),
    .A2(_144_),
    .B1(_154_),
    .B2(net14),
    .X(_155_));
 sky130_fd_sc_hd__mux2_1 _529_ (.A0(_139_),
    .A1(_155_),
    .S(_022_),
    .X(_000_));
 sky130_fd_sc_hd__and3_1 _530_ (.A(net22),
    .B(_116_),
    .C(_147_),
    .X(_156_));
 sky130_fd_sc_hd__a21o_1 _531_ (.A1(net17),
    .A2(_150_),
    .B1(net26),
    .X(_157_));
 sky130_fd_sc_hd__o21ai_1 _532_ (.A1(_156_),
    .A2(_157_),
    .B1(_132_),
    .Y(_158_));
 sky130_fd_sc_hd__or3_1 _533_ (.A(net21),
    .B(_108_),
    .C(_122_),
    .X(_159_));
 sky130_fd_sc_hd__a311o_1 _534_ (.A1(net17),
    .A2(_122_),
    .A3(_127_),
    .B1(_141_),
    .C1(net26),
    .X(_160_));
 sky130_fd_sc_hd__o32a_1 _535_ (.A1(_105_),
    .A2(net24),
    .A3(net22),
    .B1(_114_),
    .B2(_109_),
    .X(_161_));
 sky130_fd_sc_hd__nor2_1 _536_ (.A(net21),
    .B(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__o211a_1 _537_ (.A1(net21),
    .A2(_161_),
    .B1(_160_),
    .C1(_022_),
    .X(_163_));
 sky130_fd_sc_hd__a31o_1 _538_ (.A1(_130_),
    .A2(_158_),
    .A3(_159_),
    .B1(_163_),
    .X(_164_));
 sky130_fd_sc_hd__a31o_1 _539_ (.A1(net18),
    .A2(_114_),
    .A3(_116_),
    .B1(net19),
    .X(_165_));
 sky130_fd_sc_hd__a31o_1 _540_ (.A1(_017_),
    .A2(net23),
    .A3(_121_),
    .B1(_165_),
    .X(_166_));
 sky130_fd_sc_hd__nand2_1 _541_ (.A(net19),
    .B(_121_),
    .Y(_167_));
 sky130_fd_sc_hd__o211ai_4 _542_ (.A1(_125_),
    .A2(_167_),
    .B1(_166_),
    .C1(_130_),
    .Y(_168_));
 sky130_fd_sc_hd__a221o_1 _543_ (.A1(_123_),
    .A2(_131_),
    .B1(_147_),
    .B2(net17),
    .C1(net20),
    .X(_169_));
 sky130_fd_sc_hd__nor2_2 _544_ (.A(_107_),
    .B(_108_),
    .Y(_170_));
 sky130_fd_sc_hd__or2_2 _545_ (.A(_089_),
    .B(_170_),
    .X(_171_));
 sky130_fd_sc_hd__o211a_1 _546_ (.A1(_156_),
    .A2(_171_),
    .B1(_169_),
    .C1(_022_),
    .X(_172_));
 sky130_fd_sc_hd__nor2_2 _547_ (.A(net14),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a22oi_4 _548_ (.A1(net15),
    .A2(_164_),
    .B1(_168_),
    .B2(_173_),
    .Y(_001_));
 sky130_fd_sc_hd__o21a_1 _549_ (.A1(_105_),
    .A2(net24),
    .B1(_142_),
    .X(_174_));
 sky130_fd_sc_hd__o21a_1 _550_ (.A1(_145_),
    .A2(_146_),
    .B1(net22),
    .X(_175_));
 sky130_fd_sc_hd__nand2_2 _551_ (.A(_102_),
    .B(net24),
    .Y(_176_));
 sky130_fd_sc_hd__nor4_1 _552_ (.A(_098_),
    .B(net22),
    .C(_145_),
    .D(_146_),
    .Y(_177_));
 sky130_fd_sc_hd__a31o_1 _553_ (.A1(net22),
    .A2(_121_),
    .A3(_176_),
    .B1(net20),
    .X(_178_));
 sky130_fd_sc_hd__o32a_1 _554_ (.A1(net27),
    .A2(_174_),
    .A3(_175_),
    .B1(_177_),
    .B2(_178_),
    .X(_179_));
 sky130_fd_sc_hd__o211a_1 _555_ (.A1(_145_),
    .A2(_146_),
    .B1(_099_),
    .C1(net22),
    .X(_180_));
 sky130_fd_sc_hd__a21o_1 _556_ (.A1(net16),
    .A2(_126_),
    .B1(net20),
    .X(_181_));
 sky130_fd_sc_hd__a211oi_2 _557_ (.A1(_121_),
    .A2(_123_),
    .B1(net28),
    .C1(_109_),
    .Y(_182_));
 sky130_fd_sc_hd__or3_1 _558_ (.A(net27),
    .B(_142_),
    .C(_182_),
    .X(_183_));
 sky130_fd_sc_hd__o211a_1 _559_ (.A1(_180_),
    .A2(_181_),
    .B1(_183_),
    .C1(net14),
    .X(_184_));
 sky130_fd_sc_hd__a211o_1 _560_ (.A1(net13),
    .A2(_179_),
    .B1(_184_),
    .C1(_022_),
    .X(_185_));
 sky130_fd_sc_hd__o211a_4 _561_ (.A1(_100_),
    .A2(net24),
    .B1(_108_),
    .C1(_087_),
    .X(_186_));
 sky130_fd_sc_hd__a221o_1 _562_ (.A1(_114_),
    .A2(_125_),
    .B1(_186_),
    .B2(_115_),
    .C1(net20),
    .X(_187_));
 sky130_fd_sc_hd__a211o_1 _563_ (.A1(net16),
    .A2(_116_),
    .B1(_182_),
    .C1(net27),
    .X(_188_));
 sky130_fd_sc_hd__nand2_2 _564_ (.A(_346_),
    .B(_097_),
    .Y(_189_));
 sky130_fd_sc_hd__and3_1 _565_ (.A(_099_),
    .B(net16),
    .C(_189_),
    .X(_190_));
 sky130_fd_sc_hd__xnor2_2 _566_ (.A(_097_),
    .B(net24),
    .Y(_191_));
 sky130_fd_sc_hd__o22a_1 _567_ (.A1(_094_),
    .A2(net25),
    .B1(_109_),
    .B2(net28),
    .X(_192_));
 sky130_fd_sc_hd__a22o_1 _568_ (.A1(_016_),
    .A2(_107_),
    .B1(_108_),
    .B2(_087_),
    .X(_193_));
 sky130_fd_sc_hd__a211o_1 _569_ (.A1(net22),
    .A2(_191_),
    .B1(_192_),
    .C1(net27),
    .X(_194_));
 sky130_fd_sc_hd__o211a_1 _570_ (.A1(_124_),
    .A2(_190_),
    .B1(_194_),
    .C1(net14),
    .X(_195_));
 sky130_fd_sc_hd__a31o_1 _571_ (.A1(_021_),
    .A2(_187_),
    .A3(_188_),
    .B1(_195_),
    .X(_196_));
 sky130_fd_sc_hd__o21a_1 _572_ (.A1(_130_),
    .A2(_196_),
    .B1(_185_),
    .X(_002_));
 sky130_fd_sc_hd__and3_4 _573_ (.A(_016_),
    .B(net25),
    .C(_108_),
    .X(_197_));
 sky130_fd_sc_hd__a31o_1 _574_ (.A1(_099_),
    .A2(_123_),
    .A3(_192_),
    .B1(_197_),
    .X(_198_));
 sky130_fd_sc_hd__a21boi_1 _575_ (.A1(net21),
    .A2(_198_),
    .B1_N(_159_),
    .Y(_199_));
 sky130_fd_sc_hd__a31o_1 _576_ (.A1(_104_),
    .A2(net16),
    .A3(_176_),
    .B1(_197_),
    .X(_200_));
 sky130_fd_sc_hd__and4_1 _577_ (.A(net19),
    .B(_114_),
    .C(_189_),
    .D(_193_),
    .X(_201_));
 sky130_fd_sc_hd__a211o_1 _578_ (.A1(net27),
    .A2(_200_),
    .B1(_201_),
    .C1(net14),
    .X(_202_));
 sky130_fd_sc_hd__o21ai_1 _579_ (.A1(net13),
    .A2(_199_),
    .B1(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__a21oi_1 _580_ (.A1(_122_),
    .A2(_127_),
    .B1(net16),
    .Y(_204_));
 sky130_fd_sc_hd__a211o_1 _581_ (.A1(net16),
    .A2(_145_),
    .B1(_204_),
    .C1(net27),
    .X(_205_));
 sky130_fd_sc_hd__a211o_1 _582_ (.A1(_094_),
    .A2(_142_),
    .B1(_141_),
    .C1(net19),
    .X(_206_));
 sky130_fd_sc_hd__and3_1 _583_ (.A(net13),
    .B(_205_),
    .C(_206_),
    .X(_207_));
 sky130_fd_sc_hd__nand2_1 _584_ (.A(_097_),
    .B(_197_),
    .Y(_208_));
 sky130_fd_sc_hd__nand3_1 _585_ (.A(net21),
    .B(_189_),
    .C(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__a2111o_1 _586_ (.A1(_103_),
    .A2(_170_),
    .B1(_180_),
    .C1(_135_),
    .D1(net20),
    .X(_210_));
 sky130_fd_sc_hd__a31o_1 _587_ (.A1(net14),
    .A2(_209_),
    .A3(_210_),
    .B1(_022_),
    .X(_211_));
 sky130_fd_sc_hd__o22a_1 _588_ (.A1(_130_),
    .A2(_203_),
    .B1(_207_),
    .B2(_211_),
    .X(_003_));
 sky130_fd_sc_hd__nor2_2 _589_ (.A(net18),
    .B(_122_),
    .Y(_212_));
 sky130_fd_sc_hd__a221o_1 _590_ (.A1(_094_),
    .A2(_107_),
    .B1(_108_),
    .B2(_087_),
    .C1(_097_),
    .X(_213_));
 sky130_fd_sc_hd__o211a_1 _591_ (.A1(net18),
    .A2(_122_),
    .B1(_213_),
    .C1(net19),
    .X(_214_));
 sky130_fd_sc_hd__o2111a_1 _592_ (.A1(_104_),
    .A2(_111_),
    .B1(_114_),
    .C1(_189_),
    .D1(net27),
    .X(_215_));
 sky130_fd_sc_hd__nor3_1 _593_ (.A(net13),
    .B(_214_),
    .C(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__o21ai_1 _594_ (.A1(_101_),
    .A2(_192_),
    .B1(_115_),
    .Y(_217_));
 sky130_fd_sc_hd__nand2_1 _595_ (.A(net19),
    .B(_217_),
    .Y(_218_));
 sky130_fd_sc_hd__and2_2 _596_ (.A(_103_),
    .B(_111_),
    .X(_219_));
 sky130_fd_sc_hd__inv_2 _597_ (.A(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__a211o_1 _598_ (.A1(_108_),
    .A2(_113_),
    .B1(_219_),
    .C1(_020_),
    .X(_221_));
 sky130_fd_sc_hd__a31o_1 _599_ (.A1(net13),
    .A2(_218_),
    .A3(_221_),
    .B1(_216_),
    .X(_222_));
 sky130_fd_sc_hd__a32o_1 _600_ (.A1(net16),
    .A2(_151_),
    .A3(_176_),
    .B1(_186_),
    .B2(_126_),
    .X(_223_));
 sky130_fd_sc_hd__a211o_1 _601_ (.A1(net21),
    .A2(_223_),
    .B1(_162_),
    .C1(net13),
    .X(_224_));
 sky130_fd_sc_hd__o32a_1 _602_ (.A1(net19),
    .A2(_111_),
    .A3(_197_),
    .B1(_212_),
    .B2(_171_),
    .X(_225_));
 sky130_fd_sc_hd__o21a_1 _603_ (.A1(net15),
    .A2(_225_),
    .B1(_022_),
    .X(_226_));
 sky130_fd_sc_hd__a22o_1 _604_ (.A1(_130_),
    .A2(_222_),
    .B1(_224_),
    .B2(_226_),
    .X(_004_));
 sky130_fd_sc_hd__a21o_1 _605_ (.A1(_017_),
    .A2(_113_),
    .B1(net18),
    .X(_227_));
 sky130_fd_sc_hd__a31o_1 _606_ (.A1(_017_),
    .A2(net23),
    .A3(_113_),
    .B1(_219_),
    .X(_228_));
 sky130_fd_sc_hd__a211o_1 _607_ (.A1(net16),
    .A2(_150_),
    .B1(_146_),
    .C1(net20),
    .X(_229_));
 sky130_fd_sc_hd__a2bb2o_1 _608_ (.A1_N(_186_),
    .A2_N(_229_),
    .B1(_228_),
    .B2(net19),
    .X(_230_));
 sky130_fd_sc_hd__nand2_1 _609_ (.A(net15),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__or3_1 _610_ (.A(_099_),
    .B(net15),
    .C(_171_),
    .X(_232_));
 sky130_fd_sc_hd__a2111o_1 _611_ (.A1(_104_),
    .A2(net17),
    .B1(_111_),
    .C1(_186_),
    .D1(net21),
    .X(_233_));
 sky130_fd_sc_hd__a221o_1 _612_ (.A1(net23),
    .A2(_115_),
    .B1(_142_),
    .B2(_099_),
    .C1(net26),
    .X(_234_));
 sky130_fd_sc_hd__a21o_1 _613_ (.A1(_233_),
    .A2(_234_),
    .B1(net14),
    .X(_235_));
 sky130_fd_sc_hd__a21o_1 _614_ (.A1(_098_),
    .A2(_170_),
    .B1(net21),
    .X(_236_));
 sky130_fd_sc_hd__o311a_1 _615_ (.A1(net26),
    .A2(_212_),
    .A3(_219_),
    .B1(_236_),
    .C1(net15),
    .X(_237_));
 sky130_fd_sc_hd__and3b_1 _616_ (.A_N(_237_),
    .B(_130_),
    .C(_235_),
    .X(_238_));
 sky130_fd_sc_hd__a31o_1 _617_ (.A1(_022_),
    .A2(_231_),
    .A3(_232_),
    .B1(_238_),
    .X(_005_));
 sky130_fd_sc_hd__or3_1 _618_ (.A(net16),
    .B(_146_),
    .C(_150_),
    .X(_239_));
 sky130_fd_sc_hd__o21a_1 _619_ (.A1(net22),
    .A2(_115_),
    .B1(net26),
    .X(_240_));
 sky130_fd_sc_hd__a32o_1 _620_ (.A1(net21),
    .A2(_208_),
    .A3(_220_),
    .B1(_239_),
    .B2(_240_),
    .X(_241_));
 sky130_fd_sc_hd__o21a_1 _621_ (.A1(_136_),
    .A2(_142_),
    .B1(net21),
    .X(_242_));
 sky130_fd_sc_hd__a21o_1 _622_ (.A1(net26),
    .A2(_109_),
    .B1(net13),
    .X(_243_));
 sky130_fd_sc_hd__o22a_1 _623_ (.A1(net14),
    .A2(_241_),
    .B1(_242_),
    .B2(_243_),
    .X(_244_));
 sky130_fd_sc_hd__a21o_1 _624_ (.A1(_016_),
    .A2(_189_),
    .B1(net18),
    .X(_245_));
 sky130_fd_sc_hd__nand2_1 _625_ (.A(_115_),
    .B(_125_),
    .Y(_246_));
 sky130_fd_sc_hd__a32o_1 _626_ (.A1(net26),
    .A2(_227_),
    .A3(_246_),
    .B1(_245_),
    .B2(_112_),
    .X(_247_));
 sky130_fd_sc_hd__a21o_1 _627_ (.A1(_103_),
    .A2(_170_),
    .B1(net26),
    .X(_248_));
 sky130_fd_sc_hd__o211a_1 _628_ (.A1(_212_),
    .A2(_236_),
    .B1(_248_),
    .C1(net14),
    .X(_249_));
 sky130_fd_sc_hd__a21oi_1 _629_ (.A1(net13),
    .A2(_247_),
    .B1(_249_),
    .Y(_250_));
 sky130_fd_sc_hd__mux2_1 _630_ (.A0(_244_),
    .A1(_250_),
    .S(_022_),
    .X(_006_));
 sky130_fd_sc_hd__or2_1 _631_ (.A(net1),
    .B(net3),
    .X(_251_));
 sky130_fd_sc_hd__nand2_1 _632_ (.A(net1),
    .B(net3),
    .Y(_252_));
 sky130_fd_sc_hd__nand2_1 _633_ (.A(_251_),
    .B(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__xnor2_1 _634_ (.A(net2),
    .B(_253_),
    .Y(_009_));
 sky130_fd_sc_hd__a21bo_1 _635_ (.A1(net2),
    .A2(_251_),
    .B1_N(_252_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_4 _636_ (.A0(\lcd.s_ROM[4] ),
    .A1(\lcd.s_ROM[0] ),
    .S(net45),
    .X(_254_));
 sky130_fd_sc_hd__nand2_1 _637_ (.A(_037_),
    .B(_073_),
    .Y(_255_));
 sky130_fd_sc_hd__nand2_2 _638_ (.A(_057_),
    .B(_066_),
    .Y(_256_));
 sky130_fd_sc_hd__a22o_1 _639_ (.A1(_343_),
    .A2(_038_),
    .B1(_054_),
    .B2(_037_),
    .X(_257_));
 sky130_fd_sc_hd__o21a_1 _640_ (.A1(_254_),
    .A2(_255_),
    .B1(_256_),
    .X(_258_));
 sky130_fd_sc_hd__a2bb2o_1 _641_ (.A1_N(net45),
    .A2_N(_054_),
    .B1(_257_),
    .B2(_258_),
    .X(_259_));
 sky130_fd_sc_hd__a221o_1 _642_ (.A1(_062_),
    .A2(_254_),
    .B1(_259_),
    .B2(_055_),
    .C1(_046_),
    .X(_260_));
 sky130_fd_sc_hd__o22a_1 _643_ (.A1(net44),
    .A2(\lcd.num_state[1] ),
    .B1(\lcd.num_state[0] ),
    .B2(net42),
    .X(_261_));
 sky130_fd_sc_hd__o221a_1 _644_ (.A1(net42),
    .A2(net43),
    .B1(_343_),
    .B2(_261_),
    .C1(_041_),
    .X(_262_));
 sky130_fd_sc_hd__a21bo_1 _645_ (.A1(_042_),
    .A2(_254_),
    .B1_N(_057_),
    .X(_263_));
 sky130_fd_sc_hd__o21a_1 _646_ (.A1(_262_),
    .A2(_263_),
    .B1(_349_),
    .X(_264_));
 sky130_fd_sc_hd__a31o_1 _647_ (.A1(_343_),
    .A2(_348_),
    .A3(_051_),
    .B1(_045_),
    .X(_265_));
 sky130_fd_sc_hd__nor2_1 _648_ (.A(_349_),
    .B(_051_),
    .Y(_266_));
 sky130_fd_sc_hd__a211o_1 _649_ (.A1(_254_),
    .A2(_266_),
    .B1(_265_),
    .C1(_264_),
    .X(_267_));
 sky130_fd_sc_hd__o21a_1 _650_ (.A1(_082_),
    .A2(_254_),
    .B1(_033_),
    .X(_268_));
 sky130_fd_sc_hd__a31o_1 _651_ (.A1(_358_),
    .A2(_260_),
    .A3(_267_),
    .B1(_268_),
    .X(_269_));
 sky130_fd_sc_hd__or2_1 _652_ (.A(_351_),
    .B(_269_),
    .X(_270_));
 sky130_fd_sc_hd__and3_1 _653_ (.A(net46),
    .B(_348_),
    .C(_354_),
    .X(_271_));
 sky130_fd_sc_hd__a21o_1 _654_ (.A1(net41),
    .A2(net43),
    .B1(net46),
    .X(_272_));
 sky130_fd_sc_hd__or4_2 _655_ (.A(net40),
    .B(_048_),
    .C(_063_),
    .D(_272_),
    .X(_273_));
 sky130_fd_sc_hd__or4b_1 _656_ (.A(net36),
    .B(net43),
    .C(_347_),
    .D_N(net42),
    .X(_274_));
 sky130_fd_sc_hd__or3_1 _657_ (.A(_343_),
    .B(_349_),
    .C(_274_),
    .X(_275_));
 sky130_fd_sc_hd__nand3b_1 _658_ (.A_N(_271_),
    .B(_273_),
    .C(_275_),
    .Y(_276_));
 sky130_fd_sc_hd__mux2_1 _659_ (.A0(_273_),
    .A1(net44),
    .S(_271_),
    .X(_277_));
 sky130_fd_sc_hd__nor2_2 _660_ (.A(_340_),
    .B(_361_),
    .Y(_278_));
 sky130_fd_sc_hd__a32o_1 _661_ (.A1(_270_),
    .A2(_277_),
    .A3(_278_),
    .B1(net29),
    .B2(net12),
    .X(_010_));
 sky130_fd_sc_hd__mux2_4 _662_ (.A0(\lcd.s_ROM[5] ),
    .A1(\lcd.s_ROM[1] ),
    .S(net45),
    .X(_279_));
 sky130_fd_sc_hd__a21o_2 _663_ (.A1(_350_),
    .A2(_041_),
    .B1(net30),
    .X(_280_));
 sky130_fd_sc_hd__or3_1 _664_ (.A(_343_),
    .B(_043_),
    .C(_280_),
    .X(_281_));
 sky130_fd_sc_hd__a22o_1 _665_ (.A1(_266_),
    .A2(_279_),
    .B1(_281_),
    .B2(_349_),
    .X(_282_));
 sky130_fd_sc_hd__o2111a_1 _666_ (.A1(_044_),
    .A2(_279_),
    .B1(_282_),
    .C1(_046_),
    .D1(_358_),
    .X(_283_));
 sky130_fd_sc_hd__a21o_1 _667_ (.A1(net45),
    .A2(_034_),
    .B1(_037_),
    .X(_284_));
 sky130_fd_sc_hd__a32o_1 _668_ (.A1(_054_),
    .A2(_256_),
    .A3(_284_),
    .B1(_279_),
    .B2(_062_),
    .X(_285_));
 sky130_fd_sc_hd__o211a_1 _669_ (.A1(_255_),
    .A2(_279_),
    .B1(_285_),
    .C1(_045_),
    .X(_286_));
 sky130_fd_sc_hd__o21a_1 _670_ (.A1(_082_),
    .A2(_279_),
    .B1(_033_),
    .X(_287_));
 sky130_fd_sc_hd__or4_1 _671_ (.A(_351_),
    .B(_283_),
    .C(_286_),
    .D(_287_),
    .X(_288_));
 sky130_fd_sc_hd__o211a_1 _672_ (.A1(_045_),
    .A2(_275_),
    .B1(_278_),
    .C1(_273_),
    .X(_289_));
 sky130_fd_sc_hd__a22o_1 _673_ (.A1(net8),
    .A2(net29),
    .B1(_288_),
    .B2(_289_),
    .X(_011_));
 sky130_fd_sc_hd__a21boi_1 _674_ (.A1(net45),
    .A2(_038_),
    .B1_N(_256_),
    .Y(_290_));
 sky130_fd_sc_hd__mux2_2 _675_ (.A0(\lcd.s_ROM[6] ),
    .A1(\lcd.s_ROM[2] ),
    .S(net45),
    .X(_291_));
 sky130_fd_sc_hd__a41o_1 _676_ (.A1(_037_),
    .A2(_054_),
    .A3(_068_),
    .A4(_073_),
    .B1(_062_),
    .X(_292_));
 sky130_fd_sc_hd__a2bb2o_1 _677_ (.A1_N(_065_),
    .A2_N(_290_),
    .B1(_291_),
    .B2(_292_),
    .X(_293_));
 sky130_fd_sc_hd__nor2_1 _678_ (.A(net45),
    .B(_368_),
    .Y(_294_));
 sky130_fd_sc_hd__a31o_1 _679_ (.A1(_368_),
    .A2(_083_),
    .A3(_291_),
    .B1(_294_),
    .X(_295_));
 sky130_fd_sc_hd__and2_1 _680_ (.A(_357_),
    .B(_295_),
    .X(_296_));
 sky130_fd_sc_hd__a221o_1 _681_ (.A1(_348_),
    .A2(_051_),
    .B1(_291_),
    .B2(_043_),
    .C1(_045_),
    .X(_297_));
 sky130_fd_sc_hd__o211a_1 _682_ (.A1(_046_),
    .A2(_293_),
    .B1(_297_),
    .C1(_358_),
    .X(_298_));
 sky130_fd_sc_hd__or3_1 _683_ (.A(_351_),
    .B(_296_),
    .C(_298_),
    .X(_299_));
 sky130_fd_sc_hd__nand2_2 _684_ (.A(net44),
    .B(net46),
    .Y(_300_));
 sky130_fd_sc_hd__xnor2_1 _685_ (.A(net42),
    .B(_300_),
    .Y(_301_));
 sky130_fd_sc_hd__a31o_1 _686_ (.A1(net43),
    .A2(_046_),
    .A3(_271_),
    .B1(_352_),
    .X(_302_));
 sky130_fd_sc_hd__a31o_1 _687_ (.A1(_045_),
    .A2(_276_),
    .A3(_301_),
    .B1(_302_),
    .X(_303_));
 sky130_fd_sc_hd__a32o_1 _688_ (.A1(_278_),
    .A2(_299_),
    .A3(_303_),
    .B1(net29),
    .B2(net9),
    .X(_012_));
 sky130_fd_sc_hd__o21bai_1 _689_ (.A1(_057_),
    .A2(_255_),
    .B1_N(_067_),
    .Y(_304_));
 sky130_fd_sc_hd__nand2_1 _690_ (.A(\lcd.seq[0] ),
    .B(\lcd.s_ROM[3] ),
    .Y(_305_));
 sky130_fd_sc_hd__inv_2 _691_ (.A(_305_),
    .Y(_306_));
 sky130_fd_sc_hd__and2_1 _692_ (.A(_068_),
    .B(_306_),
    .X(_307_));
 sky130_fd_sc_hd__o41a_1 _693_ (.A1(net46),
    .A2(_058_),
    .A3(_065_),
    .A4(_067_),
    .B1(_054_),
    .X(_308_));
 sky130_fd_sc_hd__a21bo_1 _694_ (.A1(_304_),
    .A2(_307_),
    .B1_N(_308_),
    .X(_309_));
 sky130_fd_sc_hd__a22o_1 _695_ (.A1(_062_),
    .A2(_306_),
    .B1(_309_),
    .B2(_055_),
    .X(_310_));
 sky130_fd_sc_hd__a21o_1 _696_ (.A1(net34),
    .A2(_043_),
    .B1(_266_),
    .X(_311_));
 sky130_fd_sc_hd__a21o_1 _697_ (.A1(_306_),
    .A2(_311_),
    .B1(_265_),
    .X(_312_));
 sky130_fd_sc_hd__o211a_1 _698_ (.A1(_046_),
    .A2(_310_),
    .B1(_312_),
    .C1(_358_),
    .X(_313_));
 sky130_fd_sc_hd__a31o_1 _699_ (.A1(_368_),
    .A2(_083_),
    .A3(_306_),
    .B1(_294_),
    .X(_314_));
 sky130_fd_sc_hd__a211o_1 _700_ (.A1(_357_),
    .A2(_314_),
    .B1(_313_),
    .C1(_351_),
    .X(_315_));
 sky130_fd_sc_hd__nand2b_1 _701_ (.A_N(_359_),
    .B(_300_),
    .Y(_316_));
 sky130_fd_sc_hd__a31o_1 _702_ (.A1(_045_),
    .A2(_276_),
    .A3(_316_),
    .B1(_302_),
    .X(_317_));
 sky130_fd_sc_hd__a32o_1 _703_ (.A1(_278_),
    .A2(_315_),
    .A3(_317_),
    .B1(net29),
    .B2(net10),
    .X(_013_));
 sky130_fd_sc_hd__nor2_2 _704_ (.A(_365_),
    .B(_300_),
    .Y(_318_));
 sky130_fd_sc_hd__and3_2 _705_ (.A(net37),
    .B(net39),
    .C(_318_),
    .X(_319_));
 sky130_fd_sc_hd__and3_1 _706_ (.A(net47),
    .B(_356_),
    .C(_319_),
    .X(_320_));
 sky130_fd_sc_hd__a21oi_1 _707_ (.A1(\lcd.round[0] ),
    .A2(\lcd.round[1] ),
    .B1(_340_),
    .Y(_321_));
 sky130_fd_sc_hd__a211o_1 _708_ (.A1(net47),
    .A2(_352_),
    .B1(_321_),
    .C1(_007_),
    .X(_322_));
 sky130_fd_sc_hd__and2b_1 _709_ (.A_N(_320_),
    .B(_322_),
    .X(_323_));
 sky130_fd_sc_hd__mux2_1 _710_ (.A0(_320_),
    .A1(_323_),
    .S(\lcd.round[0] ),
    .X(_014_));
 sky130_fd_sc_hd__a22o_1 _711_ (.A1(_047_),
    .A2(_320_),
    .B1(_323_),
    .B2(\lcd.round[1] ),
    .X(_015_));
 sky130_fd_sc_hd__nor2_1 _712_ (.A(_340_),
    .B(net46),
    .Y(_324_));
 sky130_fd_sc_hd__a22o_1 _713_ (.A1(net46),
    .A2(_007_),
    .B1(_360_),
    .B2(_324_),
    .X(_024_));
 sky130_fd_sc_hd__nand2_1 _714_ (.A(_360_),
    .B(_316_),
    .Y(_325_));
 sky130_fd_sc_hd__a22o_1 _715_ (.A1(net44),
    .A2(_007_),
    .B1(_325_),
    .B2(net47),
    .X(_025_));
 sky130_fd_sc_hd__a41o_1 _716_ (.A1(_354_),
    .A2(_356_),
    .A3(_357_),
    .A4(_359_),
    .B1(_301_),
    .X(_326_));
 sky130_fd_sc_hd__a22o_1 _717_ (.A1(net42),
    .A2(_007_),
    .B1(_326_),
    .B2(net47),
    .X(_026_));
 sky130_fd_sc_hd__a31oi_1 _718_ (.A1(net42),
    .A2(net44),
    .A3(net46),
    .B1(\lcd.seq[3] ),
    .Y(_327_));
 sky130_fd_sc_hd__o21ai_1 _719_ (.A1(_318_),
    .A2(_327_),
    .B1(_360_),
    .Y(_328_));
 sky130_fd_sc_hd__a22o_1 _720_ (.A1(\lcd.seq[3] ),
    .A2(_007_),
    .B1(_328_),
    .B2(net47),
    .X(_027_));
 sky130_fd_sc_hd__nor2_1 _721_ (.A(net39),
    .B(_318_),
    .Y(_329_));
 sky130_fd_sc_hd__a31o_1 _722_ (.A1(net43),
    .A2(net46),
    .A3(_034_),
    .B1(_329_),
    .X(_330_));
 sky130_fd_sc_hd__nand2_1 _723_ (.A(_360_),
    .B(_330_),
    .Y(_331_));
 sky130_fd_sc_hd__a22o_1 _724_ (.A1(net39),
    .A2(_007_),
    .B1(_331_),
    .B2(net47),
    .X(_028_));
 sky130_fd_sc_hd__a21oi_1 _725_ (.A1(net39),
    .A2(_318_),
    .B1(net37),
    .Y(_332_));
 sky130_fd_sc_hd__o21ai_1 _726_ (.A1(_319_),
    .A2(_332_),
    .B1(_360_),
    .Y(_333_));
 sky130_fd_sc_hd__a22o_1 _727_ (.A1(net37),
    .A2(_007_),
    .B1(_333_),
    .B2(net47),
    .X(_029_));
 sky130_fd_sc_hd__and3_1 _728_ (.A(net47),
    .B(\lcd.seq[6] ),
    .C(_319_),
    .X(_334_));
 sky130_fd_sc_hd__a21oi_1 _729_ (.A1(_340_),
    .A2(net4),
    .B1(_334_),
    .Y(_335_));
 sky130_fd_sc_hd__a21o_1 _730_ (.A1(net47),
    .A2(_319_),
    .B1(\lcd.seq[6] ),
    .X(_336_));
 sky130_fd_sc_hd__and2_1 _731_ (.A(_335_),
    .B(_336_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _732_ (.A0(_334_),
    .A1(_335_),
    .S(\lcd.seq[7] ),
    .X(_031_));
 sky130_fd_sc_hd__a21o_1 _733_ (.A1(_054_),
    .A2(_304_),
    .B1(_064_),
    .X(_337_));
 sky130_fd_sc_hd__o221ai_4 _734_ (.A1(_349_),
    .A2(_051_),
    .B1(_280_),
    .B2(_342_),
    .C1(_046_),
    .Y(_338_));
 sky130_fd_sc_hd__a32o_1 _735_ (.A1(_358_),
    .A2(_337_),
    .A3(_338_),
    .B1(_033_),
    .B2(_083_),
    .X(_339_));
 sky130_fd_sc_hd__a32o_1 _736_ (.A1(_352_),
    .A2(_278_),
    .A3(_339_),
    .B1(net29),
    .B2(net5),
    .X(_032_));
 sky130_fd_sc_hd__nor2_1 _737_ (.A(net47),
    .B(net4),
    .Y(_023_));
 sky130_fd_sc_hd__dfxtp_2 _738_ (.CLK(clknet_2_2__leaf_clk),
    .D(_010_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_2 _739_ (.CLK(clknet_2_2__leaf_clk),
    .D(_011_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _740_ (.CLK(clknet_2_0__leaf_clk),
    .D(_012_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _741_ (.CLK(clknet_2_2__leaf_clk),
    .D(_013_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _742_ (.CLK(clknet_2_3__leaf_clk),
    .D(_009_),
    .Q(\lcd.num_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _743_ (.CLK(clknet_2_3__leaf_clk),
    .D(_008_),
    .Q(\lcd.num_state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _744_ (.CLK(clknet_2_0__leaf_clk),
    .D(_014_),
    .Q(\lcd.round[0] ));
 sky130_fd_sc_hd__dfxtp_4 _745_ (.CLK(clknet_2_0__leaf_clk),
    .D(_015_),
    .Q(\lcd.round[1] ));
 sky130_fd_sc_hd__dfxtp_2 _746_ (.CLK(clknet_2_2__leaf_clk),
    .D(_016_),
    .Q(\lcd.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _747_ (.CLK(clknet_2_2__leaf_clk),
    .D(_017_),
    .Q(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_4 _748_ (.CLK(clknet_2_2__leaf_clk),
    .D(net25),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_4 _749_ (.CLK(clknet_2_2__leaf_clk),
    .D(net18),
    .Q(\lcd.rom_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _750_ (.CLK(clknet_2_3__leaf_clk),
    .D(net19),
    .Q(\lcd.rom_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _751_ (.CLK(clknet_2_3__leaf_clk),
    .D(net13),
    .Q(\lcd.rom_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _752_ (.CLK(clknet_2_3__leaf_clk),
    .D(_022_),
    .Q(\lcd.rom_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _753_ (.CLK(clknet_2_1__leaf_clk),
    .D(_023_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_4 _754_ (.CLK(clknet_2_0__leaf_clk),
    .D(_007_),
    .Q(\lcd.toggle ));
 sky130_fd_sc_hd__dfxtp_1 _755_ (.CLK(clknet_2_2__leaf_clk),
    .D(_000_),
    .Q(\lcd.s_ROM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _756_ (.CLK(clknet_2_1__leaf_clk),
    .D(_001_),
    .Q(\lcd.s_ROM[1] ));
 sky130_fd_sc_hd__dfxtp_1 _757_ (.CLK(clknet_2_2__leaf_clk),
    .D(_002_),
    .Q(\lcd.s_ROM[2] ));
 sky130_fd_sc_hd__dfxtp_1 _758_ (.CLK(clknet_2_3__leaf_clk),
    .D(_003_),
    .Q(\lcd.s_ROM[3] ));
 sky130_fd_sc_hd__dfxtp_1 _759_ (.CLK(clknet_2_1__leaf_clk),
    .D(_004_),
    .Q(\lcd.s_ROM[4] ));
 sky130_fd_sc_hd__dfxtp_1 _760_ (.CLK(clknet_2_3__leaf_clk),
    .D(_005_),
    .Q(\lcd.s_ROM[5] ));
 sky130_fd_sc_hd__dfxtp_1 _761_ (.CLK(clknet_2_3__leaf_clk),
    .D(_006_),
    .Q(\lcd.s_ROM[6] ));
 sky130_fd_sc_hd__dfxtp_1 _762_ (.CLK(clknet_2_0__leaf_clk),
    .D(_024_),
    .Q(\lcd.seq[0] ));
 sky130_fd_sc_hd__dfxtp_1 _763_ (.CLK(clknet_2_0__leaf_clk),
    .D(_025_),
    .Q(\lcd.seq[1] ));
 sky130_fd_sc_hd__dfxtp_1 _764_ (.CLK(clknet_2_0__leaf_clk),
    .D(_026_),
    .Q(\lcd.seq[2] ));
 sky130_fd_sc_hd__dfxtp_2 _765_ (.CLK(clknet_2_1__leaf_clk),
    .D(_027_),
    .Q(\lcd.seq[3] ));
 sky130_fd_sc_hd__dfxtp_1 _766_ (.CLK(clknet_2_0__leaf_clk),
    .D(_028_),
    .Q(\lcd.seq[4] ));
 sky130_fd_sc_hd__dfxtp_1 _767_ (.CLK(clknet_2_3__leaf_clk),
    .D(_029_),
    .Q(\lcd.seq[5] ));
 sky130_fd_sc_hd__dfxtp_1 _768_ (.CLK(clknet_2_1__leaf_clk),
    .D(_030_),
    .Q(\lcd.seq[6] ));
 sky130_fd_sc_hd__dfxtp_1 _769_ (.CLK(clknet_2_1__leaf_clk),
    .D(_031_),
    .Q(\lcd.seq[7] ));
 sky130_fd_sc_hd__dfxtp_1 _770_ (.CLK(clknet_2_0__leaf_clk),
    .D(_032_),
    .Q(net5));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_74 (.LO(net74));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_2 _798_ (.A(net12),
    .X(net7));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(rst),
    .X(net4));
 sky130_fd_sc_hd__buf_4 output5 (.A(net5),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output6 (.A(net6),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output7 (.A(net7),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output8 (.A(net8),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output9 (.A(net9),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output10 (.A(net10),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output11 (.A(net11),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_4 fanout13 (.A(_021_),
    .X(net13));
 sky130_fd_sc_hd__buf_4 fanout14 (.A(_120_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(_120_),
    .X(net15));
 sky130_fd_sc_hd__buf_4 fanout16 (.A(net18),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net18),
    .X(net17));
 sky130_fd_sc_hd__buf_4 fanout18 (.A(_019_),
    .X(net18));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(_020_),
    .X(net19));
 sky130_fd_sc_hd__buf_4 fanout20 (.A(_020_),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout21 (.A(_020_),
    .X(net21));
 sky130_fd_sc_hd__buf_4 fanout22 (.A(_110_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(_110_),
    .X(net23));
 sky130_fd_sc_hd__buf_6 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_4 fanout25 (.A(_018_),
    .X(net25));
 sky130_fd_sc_hd__buf_4 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout27 (.A(_089_),
    .X(net27));
 sky130_fd_sc_hd__buf_8 fanout28 (.A(_086_),
    .X(net28));
 sky130_fd_sc_hd__buf_4 fanout29 (.A(_363_),
    .X(net29));
 sky130_fd_sc_hd__buf_4 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(\lcd.seq[7] ),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_8 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__buf_4 fanout34 (.A(\lcd.seq[6] ),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_4 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(\lcd.seq[5] ),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(\lcd.seq[4] ),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(\lcd.seq[3] ),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(\lcd.seq[2] ),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(\lcd.seq[1] ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(\lcd.seq[1] ),
    .X(net44));
 sky130_fd_sc_hd__buf_6 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_6 fanout46 (.A(\lcd.seq[0] ),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(\lcd.toggle ),
    .X(net47));
 sky130_fd_sc_hd__conb_1 tt2_tholin_namebadge_48 (.LO(net48));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__746__D (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__A1 (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__573__A (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__568__A1 (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__514__B (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__A (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__467__B (.DIODE(_016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__752__D (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__630__S (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__617__A1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__603__B1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__587__B1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__560__C1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__546__C1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__537__C1 (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__529__S (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__503__A (.DIODE(_022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__722__A3 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__667__A2 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__422__A2 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__409__A2 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__408__A2 (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__405__A (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__404__D (.DIODE(_034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__438__A2 (.DIODE(_053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__437__A2 (.DIODE(_053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__590__C1 (.DIODE(_097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__584__A (.DIODE(_097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__566__A (.DIODE(_097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__564__B (.DIODE(_097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__A1 (.DIODE(_097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__A (.DIODE(_097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__612__B2 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__610__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__574__A1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__565__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__555__B1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__524__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__523__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__521__B1 (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__A (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__B (.DIODE(_099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__611__A1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__592__A1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__576__A1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__525__A1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__516__A1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__A (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__499__A2 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__590__A2 (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__568__A2 (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__544__A (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__524__B (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__523__B (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__499__B1 (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__487__B (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__B (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__477__A (.DIODE(_107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__622__A2 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__567__B1 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__557__C1 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__535__B2 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__521__C1 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__515__A2 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__506__A2 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__B1 (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__B (.DIODE(_109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__557__A1 (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__553__A2 (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__541__B (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__540__A3 (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__526__A2 (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__513__A1 (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__C (.DIODE(_121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__591__A2 (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__589__B (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__580__A1 (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__534__A2 (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__533__C (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__508__B (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__A2 (.DIODE(_122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__650__A2 (.DIODE(_254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__649__A1 (.DIODE(_254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__645__A2 (.DIODE(_254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__642__A2 (.DIODE(_254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__640__A1 (.DIODE(_254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__670__A2 (.DIODE(_279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__669__A2 (.DIODE(_279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__668__B1 (.DIODE(_279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__666__A2 (.DIODE(_279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__665__A2 (.DIODE(_279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__729__A1 (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__712__A (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__707__B1 (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__660__A (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__451__B1 (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__450__B1 (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__438__B1 (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__437__B1 (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__391__A (.DIODE(_340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__716__A3 (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__700__A1 (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__680__A (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__451__A1 (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__450__A1 (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__435__A (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__399__A (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__C (.DIODE(_357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__699__A1 (.DIODE(_368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__679__A1 (.DIODE(_368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__678__B (.DIODE(_368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__406__A0 (.DIODE(_368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__399__B (.DIODE(_368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA__486__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__471__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__463__B1 (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__444__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__374__A (.DIODE(\lcd.rom_addr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_output5_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__736__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output8_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__673__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__703__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output11_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__493__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__446__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__375__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_output12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__798__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__661__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__560__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__517__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__583__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__622__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__601__C1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__579__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__593__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__599__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__751__D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__629__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__749__D (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__605__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__539__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__589__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__591__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__567__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__748__D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__573__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__515__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__557__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__506__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__567__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__455__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__476__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__502__C1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__482__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__636__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__675__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__662__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__458__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__372__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__678__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__667__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__641__A1_N (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__441__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__674__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__693__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__722__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__718__A3 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__389__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__684__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__713__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__712__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__654__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__653__A (.DIODE(net46));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_236 ();
 assign io_oeb[0] = net48;
 assign io_oeb[10] = net58;
 assign io_oeb[11] = net59;
 assign io_oeb[12] = net60;
 assign io_oeb[13] = net61;
 assign io_oeb[14] = net62;
 assign io_oeb[15] = net63;
 assign io_oeb[16] = net64;
 assign io_oeb[17] = net65;
 assign io_oeb[18] = net66;
 assign io_oeb[19] = net67;
 assign io_oeb[1] = net49;
 assign io_oeb[20] = net68;
 assign io_oeb[21] = net69;
 assign io_oeb[22] = net70;
 assign io_oeb[23] = net71;
 assign io_oeb[24] = net72;
 assign io_oeb[25] = net73;
 assign io_oeb[26] = net74;
 assign io_oeb[2] = net50;
 assign io_oeb[3] = net51;
 assign io_oeb[4] = net52;
 assign io_oeb[5] = net53;
 assign io_oeb[6] = net54;
 assign io_oeb[7] = net55;
 assign io_oeb[8] = net56;
 assign io_oeb[9] = net57;
endmodule

