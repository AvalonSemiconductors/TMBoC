magic
tech sky130B
magscale 1 2
timestamp 1682095494
<< viali >>
rect 13369 19465 13403 19499
rect 17969 19465 18003 19499
rect 10977 19397 11011 19431
rect 12256 19397 12290 19431
rect 14381 19397 14415 19431
rect 15301 19397 15335 19431
rect 18797 19397 18831 19431
rect 2329 19329 2363 19363
rect 2513 19329 2547 19363
rect 14565 19329 14599 19363
rect 17141 19329 17175 19363
rect 18153 19329 18187 19363
rect 18613 19329 18647 19363
rect 11989 19261 12023 19295
rect 17417 19261 17451 19295
rect 2145 19125 2179 19159
rect 11069 19125 11103 19159
rect 14749 19125 14783 19159
rect 15393 19125 15427 19159
rect 17233 19125 17267 19159
rect 17325 19125 17359 19159
rect 7021 18921 7055 18955
rect 10701 18853 10735 18887
rect 13093 18853 13127 18887
rect 15117 18853 15151 18887
rect 17049 18785 17083 18819
rect 5365 18717 5399 18751
rect 8401 18717 8435 18751
rect 9321 18717 9355 18751
rect 11713 18717 11747 18751
rect 11980 18717 12014 18751
rect 14933 18717 14967 18751
rect 16405 18717 16439 18751
rect 16497 18717 16531 18751
rect 17325 18717 17359 18751
rect 17417 18717 17451 18751
rect 17509 18717 17543 18751
rect 17693 18717 17727 18751
rect 2329 18649 2363 18683
rect 3065 18649 3099 18683
rect 5098 18649 5132 18683
rect 8156 18649 8190 18683
rect 9588 18649 9622 18683
rect 14749 18649 14783 18683
rect 15577 18649 15611 18683
rect 15761 18649 15795 18683
rect 3985 18581 4019 18615
rect 15945 18581 15979 18615
rect 8953 18377 8987 18411
rect 4914 18309 4948 18343
rect 7840 18309 7874 18343
rect 9680 18309 9714 18343
rect 17141 18309 17175 18343
rect 2053 18241 2087 18275
rect 2145 18241 2179 18275
rect 2789 18241 2823 18275
rect 2973 18241 3007 18275
rect 7573 18241 7607 18275
rect 12072 18241 12106 18275
rect 14749 18241 14783 18275
rect 14933 18241 14967 18275
rect 15025 18241 15059 18275
rect 15577 18241 15611 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 17785 18241 17819 18275
rect 17969 18241 18003 18275
rect 5181 18173 5215 18207
rect 9413 18173 9447 18207
rect 11805 18173 11839 18207
rect 15945 18173 15979 18207
rect 17049 18173 17083 18207
rect 3801 18105 3835 18139
rect 15577 18105 15611 18139
rect 15761 18105 15795 18139
rect 16865 18105 16899 18139
rect 2329 18037 2363 18071
rect 3157 18037 3191 18071
rect 10793 18037 10827 18071
rect 13185 18037 13219 18071
rect 15853 18037 15887 18071
rect 17877 18037 17911 18071
rect 14657 17833 14691 17867
rect 18705 17833 18739 17867
rect 19625 17833 19659 17867
rect 7297 17765 7331 17799
rect 16865 17765 16899 17799
rect 15025 17697 15059 17731
rect 16313 17697 16347 17731
rect 1869 17629 1903 17663
rect 2053 17629 2087 17663
rect 2145 17629 2179 17663
rect 5190 17629 5224 17663
rect 5457 17629 5491 17663
rect 5917 17629 5951 17663
rect 14841 17629 14875 17663
rect 16497 17629 16531 17663
rect 18337 17629 18371 17663
rect 6184 17561 6218 17595
rect 15577 17561 15611 17595
rect 15761 17561 15795 17595
rect 16681 17561 16715 17595
rect 18521 17561 18555 17595
rect 19593 17561 19627 17595
rect 19809 17561 19843 17595
rect 1967 17493 2001 17527
rect 4077 17493 4111 17527
rect 16589 17493 16623 17527
rect 19441 17493 19475 17527
rect 2145 17153 2179 17187
rect 4822 17153 4856 17187
rect 5089 17153 5123 17187
rect 9956 17153 9990 17187
rect 11980 17153 12014 17187
rect 16957 17153 16991 17187
rect 19441 17153 19475 17187
rect 19625 17153 19659 17187
rect 1869 17085 1903 17119
rect 9689 17085 9723 17119
rect 11713 17085 11747 17119
rect 17509 17085 17543 17119
rect 1961 17017 1995 17051
rect 3709 17017 3743 17051
rect 2329 16949 2363 16983
rect 11069 16949 11103 16983
rect 13093 16949 13127 16983
rect 19533 16949 19567 16983
rect 10609 16745 10643 16779
rect 16681 16745 16715 16779
rect 13461 16677 13495 16711
rect 15393 16677 15427 16711
rect 2329 16609 2363 16643
rect 9229 16609 9263 16643
rect 12081 16609 12115 16643
rect 2053 16541 2087 16575
rect 2145 16541 2179 16575
rect 6653 16541 6687 16575
rect 7113 16541 7147 16575
rect 15025 16541 15059 16575
rect 15209 16541 15243 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 17969 16541 18003 16575
rect 19441 16541 19475 16575
rect 19625 16541 19659 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 6386 16473 6420 16507
rect 7380 16473 7414 16507
rect 9474 16473 9508 16507
rect 12348 16473 12382 16507
rect 16589 16473 16623 16507
rect 17417 16473 17451 16507
rect 17785 16473 17819 16507
rect 20085 16473 20119 16507
rect 5273 16405 5307 16439
rect 8493 16405 8527 16439
rect 17601 16405 17635 16439
rect 17693 16405 17727 16439
rect 2237 16201 2271 16235
rect 2789 16201 2823 16235
rect 14473 16201 14507 16235
rect 15301 16201 15335 16235
rect 17601 16201 17635 16235
rect 19809 16201 19843 16235
rect 3902 16133 3936 16167
rect 12440 16133 12474 16167
rect 1961 16065 1995 16099
rect 2053 16065 2087 16099
rect 4169 16065 4203 16099
rect 5742 16065 5776 16099
rect 6009 16065 6043 16099
rect 8033 16065 8067 16099
rect 8300 16065 8334 16099
rect 12173 16065 12207 16099
rect 14289 16065 14323 16099
rect 14473 16065 14507 16099
rect 16129 16065 16163 16099
rect 16313 16065 16347 16099
rect 16865 16065 16899 16099
rect 16957 16065 16991 16099
rect 17141 16065 17175 16099
rect 17601 16065 17635 16099
rect 18337 16065 18371 16099
rect 18521 16065 18555 16099
rect 18613 16065 18647 16099
rect 19625 16065 19659 16099
rect 15025 15997 15059 16031
rect 15209 15997 15243 16031
rect 17877 15997 17911 16031
rect 19441 15997 19475 16031
rect 15669 15929 15703 15963
rect 17141 15929 17175 15963
rect 17693 15929 17727 15963
rect 18337 15929 18371 15963
rect 4629 15861 4663 15895
rect 9413 15861 9447 15895
rect 13553 15861 13587 15895
rect 16129 15861 16163 15895
rect 5733 15657 5767 15691
rect 11713 15657 11747 15691
rect 15393 15657 15427 15691
rect 17417 15657 17451 15691
rect 17601 15657 17635 15691
rect 1961 15589 1995 15623
rect 15025 15521 15059 15555
rect 2237 15453 2271 15487
rect 15209 15453 15243 15487
rect 1961 15385 1995 15419
rect 7021 15385 7055 15419
rect 10425 15385 10459 15419
rect 17233 15385 17267 15419
rect 17449 15385 17483 15419
rect 2145 15317 2179 15351
rect 2513 15113 2547 15147
rect 9597 15113 9631 15147
rect 8309 15045 8343 15079
rect 2329 14977 2363 15011
rect 11713 14977 11747 15011
rect 11980 14977 12014 15011
rect 19533 14977 19567 15011
rect 2053 14909 2087 14943
rect 2145 14909 2179 14943
rect 14933 14909 14967 14943
rect 13093 14841 13127 14875
rect 15301 14841 15335 14875
rect 15393 14773 15427 14807
rect 19625 14773 19659 14807
rect 11161 14569 11195 14603
rect 16865 14569 16899 14603
rect 16957 14569 16991 14603
rect 19993 14569 20027 14603
rect 15117 14501 15151 14535
rect 15209 14501 15243 14535
rect 19441 14501 19475 14535
rect 3985 14433 4019 14467
rect 5641 14433 5675 14467
rect 9597 14433 9631 14467
rect 2145 14365 2179 14399
rect 2237 14365 2271 14399
rect 5365 14365 5399 14399
rect 7205 14365 7239 14399
rect 9873 14365 9907 14399
rect 12173 14365 12207 14399
rect 15025 14365 15059 14399
rect 15301 14365 15335 14399
rect 16589 14365 16623 14399
rect 16773 14365 16807 14399
rect 17049 14365 17083 14399
rect 17785 14365 17819 14399
rect 17969 14365 18003 14399
rect 19809 14365 19843 14399
rect 7472 14297 7506 14331
rect 12440 14297 12474 14331
rect 19717 14297 19751 14331
rect 2421 14229 2455 14263
rect 8585 14229 8619 14263
rect 13553 14229 13587 14263
rect 14841 14229 14875 14263
rect 17325 14229 17359 14263
rect 18153 14229 18187 14263
rect 19625 14229 19659 14263
rect 9045 14025 9079 14059
rect 13553 14025 13587 14059
rect 16957 14025 16991 14059
rect 18797 14025 18831 14059
rect 2881 13957 2915 13991
rect 7674 13957 7708 13991
rect 12440 13957 12474 13991
rect 17141 13957 17175 13991
rect 18429 13957 18463 13991
rect 18629 13957 18663 13991
rect 2237 13889 2271 13923
rect 3065 13889 3099 13923
rect 3249 13889 3283 13923
rect 5089 13889 5123 13923
rect 7941 13889 7975 13923
rect 10158 13889 10192 13923
rect 14933 13889 14967 13923
rect 15393 13889 15427 13923
rect 19533 13889 19567 13923
rect 19625 13889 19659 13923
rect 19717 13889 19751 13923
rect 19901 13889 19935 13923
rect 1961 13821 1995 13855
rect 2053 13821 2087 13855
rect 5365 13821 5399 13855
rect 10425 13821 10459 13855
rect 12173 13821 12207 13855
rect 15669 13821 15703 13855
rect 17509 13821 17543 13855
rect 19257 13821 19291 13855
rect 2421 13753 2455 13787
rect 3985 13753 4019 13787
rect 15117 13753 15151 13787
rect 15301 13753 15335 13787
rect 6561 13685 6595 13719
rect 15209 13685 15243 13719
rect 17141 13685 17175 13719
rect 18613 13685 18647 13719
rect 2329 13481 2363 13515
rect 17325 13481 17359 13515
rect 19441 13481 19475 13515
rect 19625 13481 19659 13515
rect 19993 13413 20027 13447
rect 2053 13277 2087 13311
rect 2145 13277 2179 13311
rect 6009 13277 6043 13311
rect 16865 13277 16899 13311
rect 17141 13277 17175 13311
rect 6276 13209 6310 13243
rect 7389 13141 7423 13175
rect 16957 13141 16991 13175
rect 19625 13141 19659 13175
rect 19625 12937 19659 12971
rect 1869 12869 1903 12903
rect 2053 12869 2087 12903
rect 17233 12869 17267 12903
rect 18705 12869 18739 12903
rect 2145 12801 2179 12835
rect 4169 12801 4203 12835
rect 4436 12801 4470 12835
rect 8217 12801 8251 12835
rect 11713 12801 11747 12835
rect 11980 12801 12014 12835
rect 18521 12801 18555 12835
rect 19165 12801 19199 12835
rect 19257 12801 19291 12835
rect 19441 12801 19475 12835
rect 8493 12733 8527 12767
rect 18337 12733 18371 12767
rect 1869 12665 1903 12699
rect 17601 12665 17635 12699
rect 5549 12597 5583 12631
rect 9781 12597 9815 12631
rect 13093 12597 13127 12631
rect 17049 12597 17083 12631
rect 17233 12597 17267 12631
rect 15209 12393 15243 12427
rect 15669 12393 15703 12427
rect 17969 12393 18003 12427
rect 18705 12393 18739 12427
rect 19809 12393 19843 12427
rect 19993 12393 20027 12427
rect 13093 12325 13127 12359
rect 15761 12325 15795 12359
rect 19441 12325 19475 12359
rect 1685 12257 1719 12291
rect 3985 12257 4019 12291
rect 14749 12257 14783 12291
rect 17141 12257 17175 12291
rect 1777 12189 1811 12223
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 5365 12189 5399 12223
rect 5641 12189 5675 12223
rect 7205 12189 7239 12223
rect 9597 12189 9631 12223
rect 11713 12189 11747 12223
rect 14841 12189 14875 12223
rect 16129 12189 16163 12223
rect 17417 12189 17451 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 18613 12189 18647 12223
rect 18797 12189 18831 12223
rect 7450 12121 7484 12155
rect 9864 12121 9898 12155
rect 11980 12121 12014 12155
rect 17233 12121 17267 12155
rect 8585 12053 8619 12087
rect 10977 12053 11011 12087
rect 19809 12053 19843 12087
rect 1777 11849 1811 11883
rect 13737 11849 13771 11883
rect 18797 11849 18831 11883
rect 19809 11849 19843 11883
rect 3525 11781 3559 11815
rect 19441 11781 19475 11815
rect 19533 11781 19567 11815
rect 1685 11713 1719 11747
rect 1961 11713 1995 11747
rect 5181 11713 5215 11747
rect 6561 11713 6595 11747
rect 6828 11713 6862 11747
rect 12357 11713 12391 11747
rect 12624 11713 12658 11747
rect 18429 11713 18463 11747
rect 18613 11713 18647 11747
rect 19257 11713 19291 11747
rect 19625 11713 19659 11747
rect 4905 11645 4939 11679
rect 15025 11645 15059 11679
rect 17417 11645 17451 11679
rect 1961 11577 1995 11611
rect 15301 11577 15335 11611
rect 16865 11577 16899 11611
rect 17325 11577 17359 11611
rect 7941 11509 7975 11543
rect 15485 11509 15519 11543
rect 17233 11509 17267 11543
rect 17693 11509 17727 11543
rect 2237 11305 2271 11339
rect 16681 11305 16715 11339
rect 19717 11305 19751 11339
rect 6837 11237 6871 11271
rect 17325 11169 17359 11203
rect 18613 11169 18647 11203
rect 2053 11101 2087 11135
rect 2237 11101 2271 11135
rect 5457 11101 5491 11135
rect 15393 11101 15427 11135
rect 17141 11101 17175 11135
rect 18797 11101 18831 11135
rect 18889 11101 18923 11135
rect 19625 11101 19659 11135
rect 5724 11033 5758 11067
rect 15025 11033 15059 11067
rect 17049 10965 17083 10999
rect 18613 10965 18647 10999
rect 16957 10761 16991 10795
rect 18521 10761 18555 10795
rect 12532 10693 12566 10727
rect 17125 10693 17159 10727
rect 17325 10693 17359 10727
rect 18705 10693 18739 10727
rect 2237 10625 2271 10659
rect 2329 10625 2363 10659
rect 4730 10625 4764 10659
rect 4997 10625 5031 10659
rect 8033 10625 8067 10659
rect 12265 10625 12299 10659
rect 15761 10625 15795 10659
rect 18429 10625 18463 10659
rect 19441 10625 19475 10659
rect 19533 10625 19567 10659
rect 19625 10625 19659 10659
rect 2053 10557 2087 10591
rect 2145 10557 2179 10591
rect 8309 10557 8343 10591
rect 15485 10557 15519 10591
rect 3617 10489 3651 10523
rect 18705 10489 18739 10523
rect 2513 10421 2547 10455
rect 9597 10421 9631 10455
rect 13645 10421 13679 10455
rect 15209 10421 15243 10455
rect 15393 10421 15427 10455
rect 17141 10421 17175 10455
rect 19257 10421 19291 10455
rect 2789 10217 2823 10251
rect 5549 10217 5583 10251
rect 15255 10217 15289 10251
rect 16221 10217 16255 10251
rect 17601 10217 17635 10251
rect 2145 10149 2179 10183
rect 17049 10149 17083 10183
rect 12173 10081 12207 10115
rect 1869 10013 1903 10047
rect 2605 10013 2639 10047
rect 2789 10013 2823 10047
rect 7757 10013 7791 10047
rect 14933 10013 14967 10047
rect 15117 10013 15151 10047
rect 15393 10013 15427 10047
rect 16313 10013 16347 10047
rect 16589 10013 16623 10047
rect 17325 10013 17359 10047
rect 18613 10013 18647 10047
rect 19625 10013 19659 10047
rect 19901 10013 19935 10047
rect 20085 10013 20119 10047
rect 2145 9945 2179 9979
rect 7021 9945 7055 9979
rect 10425 9945 10459 9979
rect 1961 9877 1995 9911
rect 7849 9877 7883 9911
rect 15025 9877 15059 9911
rect 16037 9877 16071 9911
rect 17233 9877 17267 9911
rect 17417 9877 17451 9911
rect 18797 9877 18831 9911
rect 19441 9877 19475 9911
rect 17325 9673 17359 9707
rect 12532 9605 12566 9639
rect 17969 9605 18003 9639
rect 19533 9605 19567 9639
rect 4638 9537 4672 9571
rect 4905 9537 4939 9571
rect 7757 9537 7791 9571
rect 8024 9537 8058 9571
rect 9781 9537 9815 9571
rect 10048 9537 10082 9571
rect 12265 9537 12299 9571
rect 14933 9537 14967 9571
rect 17417 9537 17451 9571
rect 17877 9537 17911 9571
rect 18061 9537 18095 9571
rect 19349 9537 19383 9571
rect 19625 9537 19659 9571
rect 19717 9537 19751 9571
rect 15209 9469 15243 9503
rect 13645 9401 13679 9435
rect 19901 9401 19935 9435
rect 3525 9333 3559 9367
rect 9137 9333 9171 9367
rect 11161 9333 11195 9367
rect 15025 9333 15059 9367
rect 15117 9333 15151 9367
rect 4261 9129 4295 9163
rect 6561 9129 6595 9163
rect 13553 9129 13587 9163
rect 15071 9129 15105 9163
rect 17233 9129 17267 9163
rect 17417 9129 17451 9163
rect 19901 9129 19935 9163
rect 8493 9061 8527 9095
rect 15209 9061 15243 9095
rect 2605 8993 2639 9027
rect 9781 8993 9815 9027
rect 15301 8993 15335 9027
rect 2697 8925 2731 8959
rect 4169 8925 4203 8959
rect 4353 8925 4387 8959
rect 5181 8925 5215 8959
rect 7113 8925 7147 8959
rect 9137 8925 9171 8959
rect 12173 8925 12207 8959
rect 14933 8925 14967 8959
rect 19533 8925 19567 8959
rect 19625 8925 19659 8959
rect 19717 8925 19751 8959
rect 5426 8857 5460 8891
rect 7380 8857 7414 8891
rect 10048 8857 10082 8891
rect 12440 8857 12474 8891
rect 17049 8857 17083 8891
rect 1869 8789 1903 8823
rect 9229 8789 9263 8823
rect 11161 8789 11195 8823
rect 15577 8789 15611 8823
rect 17249 8789 17283 8823
rect 4629 8585 4663 8619
rect 5733 8585 5767 8619
rect 6745 8585 6779 8619
rect 7941 8585 7975 8619
rect 10793 8585 10827 8619
rect 12909 8585 12943 8619
rect 14749 8585 14783 8619
rect 17509 8585 17543 8619
rect 19533 8585 19567 8619
rect 8861 8517 8895 8551
rect 9781 8517 9815 8551
rect 10149 8517 10183 8551
rect 11865 8517 11899 8551
rect 12081 8517 12115 8551
rect 14013 8517 14047 8551
rect 15301 8517 15335 8551
rect 15393 8517 15427 8551
rect 16957 8517 16991 8551
rect 2053 8449 2087 8483
rect 2237 8449 2271 8483
rect 5641 8449 5675 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 7757 8449 7791 8483
rect 9229 8449 9263 8483
rect 9321 8449 9355 8483
rect 10241 8449 10275 8483
rect 11161 8449 11195 8483
rect 12850 8449 12884 8483
rect 13369 8449 13403 8483
rect 13921 8449 13955 8483
rect 15025 8449 15059 8483
rect 16129 8449 16163 8483
rect 16313 8449 16347 8483
rect 16865 8449 16899 8483
rect 17233 8449 17267 8483
rect 19165 8449 19199 8483
rect 3985 8381 4019 8415
rect 4353 8381 4387 8415
rect 4445 8381 4479 8415
rect 8953 8381 8987 8415
rect 9873 8381 9907 8415
rect 11069 8381 11103 8415
rect 14933 8381 14967 8415
rect 17325 8381 17359 8415
rect 19257 8381 19291 8415
rect 13277 8313 13311 8347
rect 16221 8313 16255 8347
rect 9045 8245 9079 8279
rect 9965 8245 9999 8279
rect 11161 8245 11195 8279
rect 11713 8245 11747 8279
rect 11897 8245 11931 8279
rect 12725 8245 12759 8279
rect 19165 8245 19199 8279
rect 6653 8041 6687 8075
rect 7665 8041 7699 8075
rect 9321 8041 9355 8075
rect 11345 8041 11379 8075
rect 12081 8041 12115 8075
rect 12909 8041 12943 8075
rect 17233 8041 17267 8075
rect 18797 8041 18831 8075
rect 19625 8041 19659 8075
rect 4537 7973 4571 8007
rect 12173 7973 12207 8007
rect 2053 7905 2087 7939
rect 7573 7905 7607 7939
rect 7757 7905 7791 7939
rect 12265 7905 12299 7939
rect 17325 7905 17359 7939
rect 2237 7837 2271 7871
rect 4353 7837 4387 7871
rect 4629 7837 4663 7871
rect 4997 7837 5031 7871
rect 6009 7837 6043 7871
rect 6193 7837 6227 7871
rect 6837 7837 6871 7871
rect 7849 7837 7883 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 11069 7837 11103 7871
rect 11989 7837 12023 7871
rect 12725 7837 12759 7871
rect 14381 7837 14415 7871
rect 14841 7837 14875 7871
rect 17049 7837 17083 7871
rect 17969 7837 18003 7871
rect 18245 7837 18279 7871
rect 18705 7837 18739 7871
rect 18889 7837 18923 7871
rect 7021 7769 7055 7803
rect 11161 7769 11195 7803
rect 11345 7769 11379 7803
rect 14565 7769 14599 7803
rect 19809 7769 19843 7803
rect 2421 7701 2455 7735
rect 6193 7701 6227 7735
rect 9505 7701 9539 7735
rect 16865 7701 16899 7735
rect 19441 7701 19475 7735
rect 19609 7701 19643 7735
rect 4077 7497 4111 7531
rect 4445 7497 4479 7531
rect 5181 7497 5215 7531
rect 19441 7497 19475 7531
rect 10057 7429 10091 7463
rect 10241 7429 10275 7463
rect 13553 7429 13587 7463
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 4261 7361 4295 7395
rect 4537 7361 4571 7395
rect 5089 7361 5123 7395
rect 5273 7361 5307 7395
rect 5917 7361 5951 7395
rect 10333 7361 10367 7395
rect 13829 7361 13863 7395
rect 14841 7361 14875 7395
rect 15025 7361 15059 7395
rect 15761 7361 15795 7395
rect 16129 7361 16163 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 17141 7361 17175 7395
rect 17233 7361 17267 7395
rect 19073 7361 19107 7395
rect 19257 7361 19291 7395
rect 2329 7293 2363 7327
rect 2513 7293 2547 7327
rect 5825 7293 5859 7327
rect 13737 7293 13771 7327
rect 14473 7293 14507 7327
rect 14657 7293 14691 7327
rect 17969 7293 18003 7327
rect 18429 7293 18463 7327
rect 10057 7225 10091 7259
rect 14013 7225 14047 7259
rect 15577 7225 15611 7259
rect 18061 7225 18095 7259
rect 2145 7157 2179 7191
rect 13645 7157 13679 7191
rect 16037 7157 16071 7191
rect 17509 7157 17543 7191
rect 5181 6953 5215 6987
rect 10333 6953 10367 6987
rect 6469 6885 6503 6919
rect 11713 6885 11747 6919
rect 12265 6885 12299 6919
rect 17417 6885 17451 6919
rect 5365 6817 5399 6851
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 12909 6817 12943 6851
rect 1869 6749 1903 6783
rect 2145 6749 2179 6783
rect 5457 6749 5491 6783
rect 6285 6749 6319 6783
rect 7665 6749 7699 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 7941 6749 7975 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 13185 6749 13219 6783
rect 14289 6749 14323 6783
rect 14381 6749 14415 6783
rect 14565 6749 14599 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 17417 6749 17451 6783
rect 17877 6749 17911 6783
rect 18061 6749 18095 6783
rect 18153 6749 18187 6783
rect 10517 6681 10551 6715
rect 13001 6681 13035 6715
rect 15025 6681 15059 6715
rect 2881 6613 2915 6647
rect 7481 6613 7515 6647
rect 10149 6613 10183 6647
rect 10317 6613 10351 6647
rect 11897 6613 11931 6647
rect 18153 6613 18187 6647
rect 1961 6409 1995 6443
rect 9597 6409 9631 6443
rect 11897 6409 11931 6443
rect 12081 6409 12115 6443
rect 17893 6409 17927 6443
rect 18061 6409 18095 6443
rect 19349 6409 19383 6443
rect 3065 6341 3099 6375
rect 3801 6341 3835 6375
rect 4813 6341 4847 6375
rect 7389 6341 7423 6375
rect 17693 6341 17727 6375
rect 2053 6273 2087 6307
rect 2973 6273 3007 6307
rect 3157 6273 3191 6307
rect 3985 6273 4019 6307
rect 4997 6273 5031 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6837 6273 6871 6307
rect 7021 6273 7055 6307
rect 7757 6273 7791 6307
rect 7941 6273 7975 6307
rect 8677 6273 8711 6307
rect 8953 6273 8987 6307
rect 9137 6273 9171 6307
rect 9781 6273 9815 6307
rect 9873 6273 9907 6307
rect 10057 6273 10091 6307
rect 10149 6273 10183 6307
rect 10885 6273 10919 6307
rect 11161 6273 11195 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 17079 6273 17113 6307
rect 17233 6273 17267 6307
rect 19257 6273 19291 6307
rect 3709 6205 3743 6239
rect 5733 6205 5767 6239
rect 6561 6205 6595 6239
rect 8861 6205 8895 6239
rect 11069 6205 11103 6239
rect 12265 6205 12299 6239
rect 13921 6205 13955 6239
rect 8769 6137 8803 6171
rect 13645 6137 13679 6171
rect 16865 6137 16899 6171
rect 4261 6069 4295 6103
rect 5181 6069 5215 6103
rect 8493 6069 8527 6103
rect 10701 6069 10735 6103
rect 13461 6069 13495 6103
rect 17877 6069 17911 6103
rect 2973 5865 3007 5899
rect 10701 5865 10735 5899
rect 12909 5865 12943 5899
rect 13277 5865 13311 5899
rect 6009 5797 6043 5831
rect 8309 5797 8343 5831
rect 10793 5797 10827 5831
rect 14933 5729 14967 5763
rect 15025 5729 15059 5763
rect 15485 5729 15519 5763
rect 16405 5729 16439 5763
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 2513 5661 2547 5695
rect 3157 5661 3191 5695
rect 3341 5661 3375 5695
rect 6193 5661 6227 5695
rect 7573 5661 7607 5695
rect 7849 5661 7883 5695
rect 8401 5661 8435 5695
rect 9413 5661 9447 5695
rect 9919 5661 9953 5695
rect 10149 5661 10183 5695
rect 10701 5661 10735 5695
rect 13185 5661 13219 5695
rect 13277 5661 13311 5695
rect 15945 5661 15979 5695
rect 16497 5661 16531 5695
rect 17325 5661 17359 5695
rect 17601 5661 17635 5695
rect 6561 5593 6595 5627
rect 10977 5593 11011 5627
rect 6285 5525 6319 5559
rect 6377 5525 6411 5559
rect 10241 5525 10275 5559
rect 15301 5525 15335 5559
rect 16129 5525 16163 5559
rect 17785 5525 17819 5559
rect 6009 5321 6043 5355
rect 7297 5321 7331 5355
rect 11805 5321 11839 5355
rect 13553 5321 13587 5355
rect 13921 5321 13955 5355
rect 2973 5253 3007 5287
rect 16313 5253 16347 5287
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 7757 5185 7791 5219
rect 11713 5185 11747 5219
rect 14013 5185 14047 5219
rect 14105 5185 14139 5219
rect 15025 5185 15059 5219
rect 15301 5185 15335 5219
rect 15853 5185 15887 5219
rect 16037 5185 16071 5219
rect 2145 5117 2179 5151
rect 7665 5117 7699 5151
rect 13369 5117 13403 5151
rect 10885 4777 10919 4811
rect 12817 4777 12851 4811
rect 13185 4777 13219 4811
rect 15209 4777 15243 4811
rect 15577 4709 15611 4743
rect 5089 4641 5123 4675
rect 7389 4641 7423 4675
rect 11529 4641 11563 4675
rect 11805 4641 11839 4675
rect 13277 4641 13311 4675
rect 15485 4641 15519 4675
rect 15706 4641 15740 4675
rect 4077 4573 4111 4607
rect 6285 4573 6319 4607
rect 6377 4573 6411 4607
rect 6561 4573 6595 4607
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 7941 4573 7975 4607
rect 10609 4573 10643 4607
rect 10885 4573 10919 4607
rect 11713 4573 11747 4607
rect 11897 4573 11931 4607
rect 11989 4573 12023 4607
rect 13001 4573 13035 4607
rect 15853 4573 15887 4607
rect 10701 4505 10735 4539
rect 12909 4233 12943 4267
rect 11805 4097 11839 4131
rect 11989 4097 12023 4131
rect 12817 4097 12851 4131
rect 13001 4097 13035 4131
rect 11897 4029 11931 4063
rect 2145 2397 2179 2431
rect 4813 2397 4847 2431
rect 7481 2397 7515 2431
rect 9689 2397 9723 2431
rect 12357 2397 12391 2431
rect 15025 2397 15059 2431
rect 17693 2397 17727 2431
rect 19901 2397 19935 2431
rect 1869 2329 1903 2363
rect 4537 2329 4571 2363
rect 7205 2329 7239 2363
rect 9965 2329 9999 2363
rect 12633 2329 12667 2363
rect 15301 2329 15335 2363
rect 17969 2329 18003 2363
rect 20177 2329 20211 2363
<< metal1 >>
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 14366 19700 14372 19712
rect 11296 19672 14372 19700
rect 11296 19660 11302 19672
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 1104 19610 21043 19632
rect 1104 19558 5894 19610
rect 5946 19558 5958 19610
rect 6010 19558 6022 19610
rect 6074 19558 6086 19610
rect 6138 19558 6150 19610
rect 6202 19558 10839 19610
rect 10891 19558 10903 19610
rect 10955 19558 10967 19610
rect 11019 19558 11031 19610
rect 11083 19558 11095 19610
rect 11147 19558 15784 19610
rect 15836 19558 15848 19610
rect 15900 19558 15912 19610
rect 15964 19558 15976 19610
rect 16028 19558 16040 19610
rect 16092 19558 20729 19610
rect 20781 19558 20793 19610
rect 20845 19558 20857 19610
rect 20909 19558 20921 19610
rect 20973 19558 20985 19610
rect 21037 19558 21043 19610
rect 1104 19536 21043 19558
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 13722 19496 13728 19508
rect 13403 19468 13728 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 17957 19499 18015 19505
rect 17957 19496 17969 19499
rect 17144 19468 17969 19496
rect 10686 19388 10692 19440
rect 10744 19428 10750 19440
rect 10965 19431 11023 19437
rect 10965 19428 10977 19431
rect 10744 19400 10977 19428
rect 10744 19388 10750 19400
rect 10965 19397 10977 19400
rect 11011 19397 11023 19431
rect 10965 19391 11023 19397
rect 12244 19431 12302 19437
rect 12244 19397 12256 19431
rect 12290 19428 12302 19431
rect 14182 19428 14188 19440
rect 12290 19400 14188 19428
rect 12290 19397 12302 19400
rect 12244 19391 12302 19397
rect 14182 19388 14188 19400
rect 14240 19388 14246 19440
rect 14366 19428 14372 19440
rect 14327 19400 14372 19428
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 15289 19431 15347 19437
rect 15289 19428 15301 19431
rect 14476 19400 15301 19428
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 2406 19360 2412 19372
rect 2363 19332 2412 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 2406 19320 2412 19332
rect 2464 19320 2470 19372
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 6822 19360 6828 19372
rect 2547 19332 6828 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 6822 19320 6828 19332
rect 6880 19320 6886 19372
rect 14476 19360 14504 19400
rect 15289 19397 15301 19400
rect 15335 19397 15347 19431
rect 15289 19391 15347 19397
rect 13740 19332 14504 19360
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11756 19264 11989 19292
rect 11756 19252 11762 19264
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 2133 19159 2191 19165
rect 2133 19125 2145 19159
rect 2179 19156 2191 19159
rect 4890 19156 4896 19168
rect 2179 19128 4896 19156
rect 2179 19125 2191 19128
rect 2133 19119 2191 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 11057 19159 11115 19165
rect 11057 19125 11069 19159
rect 11103 19156 11115 19159
rect 13740 19156 13768 19332
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 14608 19332 14653 19360
rect 14608 19320 14614 19332
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 17144 19369 17172 19468
rect 17957 19465 17969 19468
rect 18003 19465 18015 19499
rect 17957 19459 18015 19465
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 18785 19431 18843 19437
rect 18785 19428 18797 19431
rect 18288 19400 18797 19428
rect 18288 19388 18294 19400
rect 18785 19397 18797 19400
rect 18831 19397 18843 19431
rect 18785 19391 18843 19397
rect 17129 19363 17187 19369
rect 17129 19360 17141 19363
rect 16264 19332 17141 19360
rect 16264 19320 16270 19332
rect 17129 19329 17141 19332
rect 17175 19329 17187 19363
rect 17129 19323 17187 19329
rect 18141 19363 18199 19369
rect 18141 19329 18153 19363
rect 18187 19360 18199 19363
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 18187 19332 18613 19360
rect 18187 19329 18199 19332
rect 18141 19323 18199 19329
rect 18601 19329 18613 19332
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19292 17463 19295
rect 19334 19292 19340 19304
rect 17451 19264 19340 19292
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 14090 19184 14096 19236
rect 14148 19224 14154 19236
rect 16574 19224 16580 19236
rect 14148 19196 16580 19224
rect 14148 19184 14154 19196
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 14734 19156 14740 19168
rect 11103 19128 13768 19156
rect 14695 19128 14740 19156
rect 11103 19125 11115 19128
rect 11057 19119 11115 19125
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15378 19156 15384 19168
rect 15339 19128 15384 19156
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 17218 19156 17224 19168
rect 17179 19128 17224 19156
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17494 19156 17500 19168
rect 17359 19128 17500 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 1104 19066 20884 19088
rect 1104 19014 3422 19066
rect 3474 19014 3486 19066
rect 3538 19014 3550 19066
rect 3602 19014 3614 19066
rect 3666 19014 3678 19066
rect 3730 19014 8367 19066
rect 8419 19014 8431 19066
rect 8483 19014 8495 19066
rect 8547 19014 8559 19066
rect 8611 19014 8623 19066
rect 8675 19014 13312 19066
rect 13364 19014 13376 19066
rect 13428 19014 13440 19066
rect 13492 19014 13504 19066
rect 13556 19014 13568 19066
rect 13620 19014 18257 19066
rect 18309 19014 18321 19066
rect 18373 19014 18385 19066
rect 18437 19014 18449 19066
rect 18501 19014 18513 19066
rect 18565 19014 20884 19066
rect 1104 18992 20884 19014
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 7009 18955 7067 18961
rect 7009 18952 7021 18955
rect 6880 18924 7021 18952
rect 6880 18912 6886 18924
rect 7009 18921 7021 18924
rect 7055 18921 7067 18955
rect 14734 18952 14740 18964
rect 7009 18915 7067 18921
rect 9140 18924 14740 18952
rect 5350 18748 5356 18760
rect 5311 18720 5356 18748
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 7616 18720 8401 18748
rect 7616 18708 7622 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 2314 18680 2320 18692
rect 2275 18652 2320 18680
rect 2314 18640 2320 18652
rect 2372 18640 2378 18692
rect 2406 18640 2412 18692
rect 2464 18680 2470 18692
rect 3053 18683 3111 18689
rect 3053 18680 3065 18683
rect 2464 18652 3065 18680
rect 2464 18640 2470 18652
rect 3053 18649 3065 18652
rect 3099 18649 3111 18683
rect 3053 18643 3111 18649
rect 4154 18640 4160 18692
rect 4212 18680 4218 18692
rect 5086 18683 5144 18689
rect 5086 18680 5098 18683
rect 4212 18652 5098 18680
rect 4212 18640 4218 18652
rect 5086 18649 5098 18652
rect 5132 18649 5144 18683
rect 5086 18643 5144 18649
rect 8144 18683 8202 18689
rect 8144 18649 8156 18683
rect 8190 18680 8202 18683
rect 9140 18680 9168 18924
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15010 18912 15016 18964
rect 15068 18952 15074 18964
rect 15068 18924 17632 18952
rect 15068 18912 15074 18924
rect 10689 18887 10747 18893
rect 10689 18853 10701 18887
rect 10735 18884 10747 18887
rect 11238 18884 11244 18896
rect 10735 18856 11244 18884
rect 10735 18853 10747 18856
rect 10689 18847 10747 18853
rect 11238 18844 11244 18856
rect 11296 18844 11302 18896
rect 13081 18887 13139 18893
rect 13081 18853 13093 18887
rect 13127 18884 13139 18887
rect 14090 18884 14096 18896
rect 13127 18856 14096 18884
rect 13127 18853 13139 18856
rect 13081 18847 13139 18853
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 15105 18887 15163 18893
rect 15105 18884 15117 18887
rect 14240 18856 15117 18884
rect 14240 18844 14246 18856
rect 15105 18853 15117 18856
rect 15151 18853 15163 18887
rect 15105 18847 15163 18853
rect 17037 18819 17095 18825
rect 17037 18816 17049 18819
rect 14016 18788 17049 18816
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 9272 18720 9321 18748
rect 9272 18708 9278 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 11698 18748 11704 18760
rect 11659 18720 11704 18748
rect 9309 18711 9367 18717
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 11968 18751 12026 18757
rect 11968 18717 11980 18751
rect 12014 18748 12026 18751
rect 14016 18748 14044 18788
rect 17037 18785 17049 18788
rect 17083 18785 17095 18819
rect 17604 18816 17632 18924
rect 17604 18788 17724 18816
rect 17037 18779 17095 18785
rect 12014 18720 14044 18748
rect 12014 18717 12026 18720
rect 11968 18711 12026 18717
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14921 18751 14979 18757
rect 14921 18748 14933 18751
rect 14608 18720 14933 18748
rect 14608 18708 14614 18720
rect 14921 18717 14933 18720
rect 14967 18748 14979 18751
rect 16393 18751 16451 18757
rect 14967 18720 15700 18748
rect 14967 18717 14979 18720
rect 14921 18711 14979 18717
rect 15672 18692 15700 18720
rect 16393 18717 16405 18751
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18748 16543 18751
rect 17218 18748 17224 18760
rect 16531 18720 17224 18748
rect 16531 18717 16543 18720
rect 16485 18711 16543 18717
rect 8190 18652 9168 18680
rect 9576 18683 9634 18689
rect 8190 18649 8202 18652
rect 8144 18643 8202 18649
rect 9576 18649 9588 18683
rect 9622 18680 9634 18683
rect 13630 18680 13636 18692
rect 9622 18652 11836 18680
rect 9622 18649 9634 18652
rect 9576 18643 9634 18649
rect 2958 18572 2964 18624
rect 3016 18612 3022 18624
rect 3973 18615 4031 18621
rect 3973 18612 3985 18615
rect 3016 18584 3985 18612
rect 3016 18572 3022 18584
rect 3973 18581 3985 18584
rect 4019 18581 4031 18615
rect 11808 18612 11836 18652
rect 12406 18652 13636 18680
rect 12406 18612 12434 18652
rect 13630 18640 13636 18652
rect 13688 18640 13694 18692
rect 14734 18680 14740 18692
rect 14695 18652 14740 18680
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 15565 18683 15623 18689
rect 15565 18680 15577 18683
rect 15028 18652 15577 18680
rect 11808 18584 12434 18612
rect 3973 18575 4031 18581
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 15028 18612 15056 18652
rect 15565 18649 15577 18652
rect 15611 18649 15623 18683
rect 15565 18643 15623 18649
rect 15654 18640 15660 18692
rect 15712 18680 15718 18692
rect 15749 18683 15807 18689
rect 15749 18680 15761 18683
rect 15712 18652 15761 18680
rect 15712 18640 15718 18652
rect 15749 18649 15761 18652
rect 15795 18649 15807 18683
rect 16408 18680 16436 18711
rect 17218 18708 17224 18720
rect 17276 18748 17282 18760
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 17276 18720 17325 18748
rect 17276 18708 17282 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 16574 18680 16580 18692
rect 16408 18652 16580 18680
rect 15749 18643 15807 18649
rect 16574 18640 16580 18652
rect 16632 18680 16638 18692
rect 17034 18680 17040 18692
rect 16632 18652 17040 18680
rect 16632 18640 16638 18652
rect 17034 18640 17040 18652
rect 17092 18640 17098 18692
rect 17420 18680 17448 18711
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 17696 18757 17724 18788
rect 17681 18751 17739 18757
rect 17552 18720 17597 18748
rect 17552 18708 17558 18720
rect 17681 18717 17693 18751
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 19334 18680 19340 18692
rect 17420 18652 19340 18680
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 13964 18584 15056 18612
rect 13964 18572 13970 18584
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 15252 18584 15945 18612
rect 15252 18572 15258 18584
rect 15933 18581 15945 18584
rect 15979 18581 15991 18615
rect 15933 18575 15991 18581
rect 1104 18522 21043 18544
rect 1104 18470 5894 18522
rect 5946 18470 5958 18522
rect 6010 18470 6022 18522
rect 6074 18470 6086 18522
rect 6138 18470 6150 18522
rect 6202 18470 10839 18522
rect 10891 18470 10903 18522
rect 10955 18470 10967 18522
rect 11019 18470 11031 18522
rect 11083 18470 11095 18522
rect 11147 18470 15784 18522
rect 15836 18470 15848 18522
rect 15900 18470 15912 18522
rect 15964 18470 15976 18522
rect 16028 18470 16040 18522
rect 16092 18470 20729 18522
rect 20781 18470 20793 18522
rect 20845 18470 20857 18522
rect 20909 18470 20921 18522
rect 20973 18470 20985 18522
rect 21037 18470 21043 18522
rect 1104 18448 21043 18470
rect 8941 18411 8999 18417
rect 8941 18377 8953 18411
rect 8987 18408 8999 18411
rect 14734 18408 14740 18420
rect 8987 18380 14740 18408
rect 8987 18377 8999 18380
rect 8941 18371 8999 18377
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 2056 18312 2820 18340
rect 2056 18284 2084 18312
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2792 18281 2820 18312
rect 4890 18300 4896 18352
rect 4948 18349 4954 18352
rect 4948 18340 4960 18349
rect 7828 18343 7886 18349
rect 4948 18312 4993 18340
rect 4948 18303 4960 18312
rect 7828 18309 7840 18343
rect 7874 18340 7886 18343
rect 8202 18340 8208 18352
rect 7874 18312 8208 18340
rect 7874 18309 7886 18312
rect 7828 18303 7886 18309
rect 4948 18300 4954 18303
rect 8202 18300 8208 18312
rect 8260 18300 8266 18352
rect 9668 18343 9726 18349
rect 9668 18309 9680 18343
rect 9714 18340 9726 18343
rect 9714 18312 14780 18340
rect 9714 18309 9726 18312
rect 9668 18303 9726 18309
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18241 2835 18275
rect 2958 18272 2964 18284
rect 2919 18244 2964 18272
rect 2777 18235 2835 18241
rect 2148 18136 2176 18235
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 7558 18272 7564 18284
rect 7519 18244 7564 18272
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 14752 18281 14780 18312
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 16632 18312 17141 18340
rect 16632 18300 16638 18312
rect 17129 18309 17141 18312
rect 17175 18340 17187 18343
rect 17862 18340 17868 18352
rect 17175 18312 17868 18340
rect 17175 18309 17187 18312
rect 17129 18303 17187 18309
rect 17862 18300 17868 18312
rect 17920 18340 17926 18352
rect 17920 18312 18000 18340
rect 17920 18300 17926 18312
rect 12060 18275 12118 18281
rect 12060 18241 12072 18275
rect 12106 18272 12118 18275
rect 14737 18275 14795 18281
rect 12106 18244 14044 18272
rect 12106 18241 12118 18244
rect 12060 18235 12118 18241
rect 5169 18207 5227 18213
rect 5169 18173 5181 18207
rect 5215 18204 5227 18207
rect 5350 18204 5356 18216
rect 5215 18176 5356 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 9272 18176 9413 18204
rect 9272 18164 9278 18176
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 9401 18167 9459 18173
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 11756 18176 11805 18204
rect 11756 18164 11762 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 3789 18139 3847 18145
rect 3789 18136 3801 18139
rect 2148 18108 3801 18136
rect 3789 18105 3801 18108
rect 3835 18105 3847 18139
rect 13906 18136 13912 18148
rect 3789 18099 3847 18105
rect 13096 18108 13912 18136
rect 2317 18071 2375 18077
rect 2317 18037 2329 18071
rect 2363 18068 2375 18071
rect 3050 18068 3056 18080
rect 2363 18040 3056 18068
rect 2363 18037 2375 18040
rect 2317 18031 2375 18037
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 6178 18068 6184 18080
rect 3191 18040 6184 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18068 10839 18071
rect 13096 18068 13124 18108
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 14016 18136 14044 18244
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14918 18272 14924 18284
rect 14879 18244 14924 18272
rect 14737 18235 14795 18241
rect 14918 18232 14924 18244
rect 14976 18232 14982 18284
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15562 18272 15568 18284
rect 15068 18244 15113 18272
rect 15523 18244 15568 18272
rect 15068 18232 15074 18244
rect 15562 18232 15568 18244
rect 15620 18232 15626 18284
rect 16666 18272 16672 18284
rect 15672 18244 16672 18272
rect 15565 18139 15623 18145
rect 15565 18136 15577 18139
rect 14016 18108 15577 18136
rect 15565 18105 15577 18108
rect 15611 18105 15623 18139
rect 15565 18099 15623 18105
rect 10827 18040 13124 18068
rect 13173 18071 13231 18077
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 13173 18037 13185 18071
rect 13219 18068 13231 18071
rect 14826 18068 14832 18080
rect 13219 18040 14832 18068
rect 13219 18037 13231 18040
rect 13173 18031 13231 18037
rect 14826 18028 14832 18040
rect 14884 18068 14890 18080
rect 15672 18068 15700 18244
rect 16666 18232 16672 18244
rect 16724 18272 16730 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16724 18244 16865 18272
rect 16724 18232 16730 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17972 18281 18000 18312
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 17000 18244 17233 18272
rect 17000 18232 17006 18244
rect 17221 18241 17233 18244
rect 17267 18272 17279 18275
rect 17773 18275 17831 18281
rect 17773 18272 17785 18275
rect 17267 18244 17785 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17773 18241 17785 18244
rect 17819 18241 17831 18275
rect 17773 18235 17831 18241
rect 17957 18275 18015 18281
rect 17957 18241 17969 18275
rect 18003 18241 18015 18275
rect 17957 18235 18015 18241
rect 15933 18207 15991 18213
rect 15933 18173 15945 18207
rect 15979 18204 15991 18207
rect 16206 18204 16212 18216
rect 15979 18176 16212 18204
rect 15979 18173 15991 18176
rect 15933 18167 15991 18173
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 17034 18204 17040 18216
rect 16995 18176 17040 18204
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 15749 18139 15807 18145
rect 15749 18105 15761 18139
rect 15795 18136 15807 18139
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 15795 18108 16865 18136
rect 15795 18105 15807 18108
rect 15749 18099 15807 18105
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 16853 18099 16911 18105
rect 15838 18068 15844 18080
rect 14884 18040 15700 18068
rect 15799 18040 15844 18068
rect 14884 18028 14890 18040
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 19334 18068 19340 18080
rect 17911 18040 19340 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 1104 17978 20884 18000
rect 1104 17926 3422 17978
rect 3474 17926 3486 17978
rect 3538 17926 3550 17978
rect 3602 17926 3614 17978
rect 3666 17926 3678 17978
rect 3730 17926 8367 17978
rect 8419 17926 8431 17978
rect 8483 17926 8495 17978
rect 8547 17926 8559 17978
rect 8611 17926 8623 17978
rect 8675 17926 13312 17978
rect 13364 17926 13376 17978
rect 13428 17926 13440 17978
rect 13492 17926 13504 17978
rect 13556 17926 13568 17978
rect 13620 17926 18257 17978
rect 18309 17926 18321 17978
rect 18373 17926 18385 17978
rect 18437 17926 18449 17978
rect 18501 17926 18513 17978
rect 18565 17926 20884 17978
rect 1104 17904 20884 17926
rect 2314 17864 2320 17876
rect 1872 17836 2320 17864
rect 1762 17620 1768 17672
rect 1820 17660 1826 17672
rect 1872 17669 1900 17836
rect 2314 17824 2320 17836
rect 2372 17864 2378 17876
rect 2372 17836 7236 17864
rect 2372 17824 2378 17836
rect 7208 17728 7236 17836
rect 13630 17824 13636 17876
rect 13688 17864 13694 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 13688 17836 14657 17864
rect 13688 17824 13694 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 18693 17867 18751 17873
rect 18693 17833 18705 17867
rect 18739 17864 18751 17867
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 18739 17836 19625 17864
rect 18739 17833 18751 17836
rect 18693 17827 18751 17833
rect 19613 17833 19625 17836
rect 19659 17833 19671 17867
rect 19613 17827 19671 17833
rect 7285 17799 7343 17805
rect 7285 17765 7297 17799
rect 7331 17796 7343 17799
rect 14918 17796 14924 17808
rect 7331 17768 14924 17796
rect 7331 17765 7343 17768
rect 7285 17759 7343 17765
rect 14918 17756 14924 17768
rect 14976 17756 14982 17808
rect 16853 17799 16911 17805
rect 15028 17768 16804 17796
rect 15028 17740 15056 17768
rect 7208 17700 12434 17728
rect 1857 17663 1915 17669
rect 1857 17660 1869 17663
rect 1820 17632 1869 17660
rect 1820 17620 1826 17632
rect 1857 17629 1869 17632
rect 1903 17629 1915 17663
rect 1857 17623 1915 17629
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 2041 17663 2099 17669
rect 2041 17660 2053 17663
rect 2004 17632 2053 17660
rect 2004 17620 2010 17632
rect 2041 17629 2053 17632
rect 2087 17629 2099 17663
rect 2041 17623 2099 17629
rect 2130 17620 2136 17672
rect 2188 17660 2194 17672
rect 2188 17632 2233 17660
rect 2188 17620 2194 17632
rect 3050 17620 3056 17672
rect 3108 17660 3114 17672
rect 5178 17663 5236 17669
rect 5178 17660 5190 17663
rect 3108 17632 5190 17660
rect 3108 17620 3114 17632
rect 5178 17629 5190 17632
rect 5224 17629 5236 17663
rect 5178 17623 5236 17629
rect 5350 17620 5356 17672
rect 5408 17660 5414 17672
rect 5445 17663 5503 17669
rect 5445 17660 5457 17663
rect 5408 17632 5457 17660
rect 5408 17620 5414 17632
rect 5445 17629 5457 17632
rect 5491 17660 5503 17663
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 5491 17632 5917 17660
rect 5491 17629 5503 17632
rect 5445 17623 5503 17629
rect 5905 17629 5917 17632
rect 5951 17660 5963 17663
rect 7558 17660 7564 17672
rect 5951 17632 7564 17660
rect 5951 17629 5963 17632
rect 5905 17623 5963 17629
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 6178 17601 6184 17604
rect 6172 17592 6184 17601
rect 6139 17564 6184 17592
rect 6172 17555 6184 17564
rect 6178 17552 6184 17555
rect 6236 17552 6242 17604
rect 12406 17592 12434 17700
rect 14182 17688 14188 17740
rect 14240 17728 14246 17740
rect 15010 17728 15016 17740
rect 14240 17700 15016 17728
rect 14240 17688 14246 17700
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 15562 17688 15568 17740
rect 15620 17728 15626 17740
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 15620 17700 16313 17728
rect 15620 17688 15626 17700
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16776 17728 16804 17768
rect 16853 17765 16865 17799
rect 16899 17796 16911 17799
rect 17034 17796 17040 17808
rect 16899 17768 17040 17796
rect 16899 17765 16911 17768
rect 16853 17759 16911 17765
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 16776 17700 19840 17728
rect 16301 17691 16359 17697
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 13780 17632 14841 17660
rect 13780 17620 13786 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17660 16543 17663
rect 16942 17660 16948 17672
rect 16531 17632 16948 17660
rect 16531 17629 16543 17632
rect 16485 17623 16543 17629
rect 16942 17620 16948 17632
rect 17000 17660 17006 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 17000 17632 18337 17660
rect 17000 17620 17006 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 19812 17604 19840 17700
rect 15378 17592 15384 17604
rect 12406 17564 15384 17592
rect 15378 17552 15384 17564
rect 15436 17592 15442 17604
rect 15565 17595 15623 17601
rect 15565 17592 15577 17595
rect 15436 17564 15577 17592
rect 15436 17552 15442 17564
rect 15565 17561 15577 17564
rect 15611 17561 15623 17595
rect 15565 17555 15623 17561
rect 15749 17595 15807 17601
rect 15749 17561 15761 17595
rect 15795 17592 15807 17595
rect 15838 17592 15844 17604
rect 15795 17564 15844 17592
rect 15795 17561 15807 17564
rect 15749 17555 15807 17561
rect 15838 17552 15844 17564
rect 15896 17592 15902 17604
rect 16298 17592 16304 17604
rect 15896 17564 16304 17592
rect 15896 17552 15902 17564
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 16666 17592 16672 17604
rect 16627 17564 16672 17592
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 17862 17552 17868 17604
rect 17920 17592 17926 17604
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 17920 17564 18521 17592
rect 17920 17552 17926 17564
rect 18509 17561 18521 17564
rect 18555 17561 18567 17595
rect 18509 17555 18567 17561
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19581 17595 19639 17601
rect 19581 17592 19593 17595
rect 19392 17564 19593 17592
rect 19392 17552 19398 17564
rect 19581 17561 19593 17564
rect 19627 17561 19639 17595
rect 19794 17592 19800 17604
rect 19707 17564 19800 17592
rect 19581 17555 19639 17561
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 1946 17524 1952 17536
rect 2004 17533 2010 17536
rect 1913 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17487 2013 17533
rect 2004 17484 2010 17487
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 4065 17527 4123 17533
rect 4065 17524 4077 17527
rect 3200 17496 4077 17524
rect 3200 17484 3206 17496
rect 4065 17493 4077 17496
rect 4111 17493 4123 17527
rect 16574 17524 16580 17536
rect 16535 17496 16580 17524
rect 4065 17487 4123 17493
rect 16574 17484 16580 17496
rect 16632 17484 16638 17536
rect 19426 17524 19432 17536
rect 19387 17496 19432 17524
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 1104 17434 21043 17456
rect 1104 17382 5894 17434
rect 5946 17382 5958 17434
rect 6010 17382 6022 17434
rect 6074 17382 6086 17434
rect 6138 17382 6150 17434
rect 6202 17382 10839 17434
rect 10891 17382 10903 17434
rect 10955 17382 10967 17434
rect 11019 17382 11031 17434
rect 11083 17382 11095 17434
rect 11147 17382 15784 17434
rect 15836 17382 15848 17434
rect 15900 17382 15912 17434
rect 15964 17382 15976 17434
rect 16028 17382 16040 17434
rect 16092 17382 20729 17434
rect 20781 17382 20793 17434
rect 20845 17382 20857 17434
rect 20909 17382 20921 17434
rect 20973 17382 20985 17434
rect 21037 17382 21043 17434
rect 1104 17360 21043 17382
rect 1946 17144 1952 17196
rect 2004 17184 2010 17196
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 2004 17156 2145 17184
rect 2004 17144 2010 17156
rect 2133 17153 2145 17156
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 4246 17144 4252 17196
rect 4304 17184 4310 17196
rect 4810 17187 4868 17193
rect 4810 17184 4822 17187
rect 4304 17156 4822 17184
rect 4304 17144 4310 17156
rect 4810 17153 4822 17156
rect 4856 17153 4868 17187
rect 4810 17147 4868 17153
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5350 17184 5356 17196
rect 5123 17156 5356 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 9944 17187 10002 17193
rect 9944 17153 9956 17187
rect 9990 17184 10002 17187
rect 11146 17184 11152 17196
rect 9990 17156 11152 17184
rect 9990 17153 10002 17156
rect 9944 17147 10002 17153
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 11968 17187 12026 17193
rect 11968 17153 11980 17187
rect 12014 17184 12026 17187
rect 13722 17184 13728 17196
rect 12014 17156 13728 17184
rect 12014 17153 12026 17156
rect 11968 17147 12026 17153
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16945 17187 17003 17193
rect 16945 17184 16957 17187
rect 15436 17156 16957 17184
rect 15436 17144 15442 17156
rect 16945 17153 16957 17156
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 19518 17184 19524 17196
rect 19475 17156 19524 17184
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17184 19671 17187
rect 19702 17184 19708 17196
rect 19659 17156 19708 17184
rect 19659 17153 19671 17156
rect 19613 17147 19671 17153
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 1854 17116 1860 17128
rect 1815 17088 1860 17116
rect 1854 17076 1860 17088
rect 1912 17076 1918 17128
rect 9214 17076 9220 17128
rect 9272 17116 9278 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9272 17088 9689 17116
rect 9272 17076 9278 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 11698 17116 11704 17128
rect 11659 17088 11704 17116
rect 9677 17079 9735 17085
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 17494 17116 17500 17128
rect 17455 17088 17500 17116
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 1949 17051 2007 17057
rect 1949 17017 1961 17051
rect 1995 17048 2007 17051
rect 2130 17048 2136 17060
rect 1995 17020 2136 17048
rect 1995 17017 2007 17020
rect 1949 17011 2007 17017
rect 2130 17008 2136 17020
rect 2188 17048 2194 17060
rect 3697 17051 3755 17057
rect 3697 17048 3709 17051
rect 2188 17020 3709 17048
rect 2188 17008 2194 17020
rect 3697 17017 3709 17020
rect 3743 17017 3755 17051
rect 16850 17048 16856 17060
rect 3697 17011 3755 17017
rect 13004 17020 16856 17048
rect 2317 16983 2375 16989
rect 2317 16949 2329 16983
rect 2363 16980 2375 16983
rect 3878 16980 3884 16992
rect 2363 16952 3884 16980
rect 2363 16949 2375 16952
rect 2317 16943 2375 16949
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 11057 16983 11115 16989
rect 11057 16949 11069 16983
rect 11103 16980 11115 16983
rect 13004 16980 13032 17020
rect 16850 17008 16856 17020
rect 16908 17008 16914 17060
rect 11103 16952 13032 16980
rect 13081 16983 13139 16989
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 13081 16949 13093 16983
rect 13127 16980 13139 16983
rect 14274 16980 14280 16992
rect 13127 16952 14280 16980
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 14274 16940 14280 16952
rect 14332 16980 14338 16992
rect 15102 16980 15108 16992
rect 14332 16952 15108 16980
rect 14332 16940 14338 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 19521 16983 19579 16989
rect 19521 16949 19533 16983
rect 19567 16980 19579 16983
rect 19610 16980 19616 16992
rect 19567 16952 19616 16980
rect 19567 16949 19579 16952
rect 19521 16943 19579 16949
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 1104 16890 20884 16912
rect 1104 16838 3422 16890
rect 3474 16838 3486 16890
rect 3538 16838 3550 16890
rect 3602 16838 3614 16890
rect 3666 16838 3678 16890
rect 3730 16838 8367 16890
rect 8419 16838 8431 16890
rect 8483 16838 8495 16890
rect 8547 16838 8559 16890
rect 8611 16838 8623 16890
rect 8675 16838 13312 16890
rect 13364 16838 13376 16890
rect 13428 16838 13440 16890
rect 13492 16838 13504 16890
rect 13556 16838 13568 16890
rect 13620 16838 18257 16890
rect 18309 16838 18321 16890
rect 18373 16838 18385 16890
rect 18437 16838 18449 16890
rect 18501 16838 18513 16890
rect 18565 16838 20884 16890
rect 1104 16816 20884 16838
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 8294 16776 8300 16788
rect 4028 16748 8300 16776
rect 4028 16736 4034 16748
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 10594 16776 10600 16788
rect 10555 16748 10600 16776
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 11204 16748 16681 16776
rect 11204 16736 11210 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 2774 16708 2780 16720
rect 2148 16680 2780 16708
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2148 16581 2176 16680
rect 2774 16668 2780 16680
rect 2832 16668 2838 16720
rect 13449 16711 13507 16717
rect 13449 16677 13461 16711
rect 13495 16708 13507 16711
rect 13630 16708 13636 16720
rect 13495 16680 13636 16708
rect 13495 16677 13507 16680
rect 13449 16671 13507 16677
rect 13630 16668 13636 16680
rect 13688 16668 13694 16720
rect 15381 16711 15439 16717
rect 15381 16677 15393 16711
rect 15427 16708 15439 16711
rect 16574 16708 16580 16720
rect 15427 16680 16580 16708
rect 15427 16677 15439 16680
rect 15381 16671 15439 16677
rect 16574 16668 16580 16680
rect 16632 16668 16638 16720
rect 19794 16708 19800 16720
rect 19444 16680 19800 16708
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 5442 16640 5448 16652
rect 2363 16612 5448 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 9214 16640 9220 16652
rect 9175 16612 9220 16640
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12069 16643 12127 16649
rect 12069 16640 12081 16643
rect 11756 16612 12081 16640
rect 11756 16600 11762 16612
rect 12069 16609 12081 16612
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 14936 16612 15240 16640
rect 14936 16584 14964 16612
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 6641 16575 6699 16581
rect 6641 16541 6653 16575
rect 6687 16572 6699 16575
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6687 16544 7113 16572
rect 6687 16541 6699 16544
rect 6641 16535 6699 16541
rect 7101 16541 7113 16544
rect 7147 16572 7159 16575
rect 10502 16572 10508 16584
rect 7147 16544 7604 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 7576 16516 7604 16544
rect 8404 16544 10508 16572
rect 2222 16464 2228 16516
rect 2280 16504 2286 16516
rect 6374 16507 6432 16513
rect 6374 16504 6386 16507
rect 2280 16476 6386 16504
rect 2280 16464 2286 16476
rect 6374 16473 6386 16476
rect 6420 16473 6432 16507
rect 6374 16467 6432 16473
rect 7368 16507 7426 16513
rect 7368 16473 7380 16507
rect 7414 16504 7426 16507
rect 7414 16476 7512 16504
rect 7414 16473 7426 16476
rect 7368 16467 7426 16473
rect 5258 16436 5264 16448
rect 5219 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 7484 16436 7512 16476
rect 7558 16464 7564 16516
rect 7616 16464 7622 16516
rect 8404 16436 8432 16544
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 14918 16572 14924 16584
rect 10612 16544 14924 16572
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9462 16507 9520 16513
rect 9462 16504 9474 16507
rect 9364 16476 9474 16504
rect 9364 16464 9370 16476
rect 9462 16473 9474 16476
rect 9508 16473 9520 16507
rect 10612 16504 10640 16544
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 15010 16532 15016 16584
rect 15068 16572 15074 16584
rect 15212 16581 15240 16612
rect 15197 16575 15255 16581
rect 15068 16544 15113 16572
rect 15068 16532 15074 16544
rect 15197 16541 15209 16575
rect 15243 16541 15255 16575
rect 16758 16572 16764 16584
rect 16719 16544 16764 16572
rect 15197 16535 15255 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 16942 16572 16948 16584
rect 16899 16544 16948 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 16942 16532 16948 16544
rect 17000 16572 17006 16584
rect 17957 16575 18015 16581
rect 17957 16572 17969 16575
rect 17000 16544 17969 16572
rect 17000 16532 17006 16544
rect 17957 16541 17969 16544
rect 18003 16541 18015 16575
rect 17957 16535 18015 16541
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 19334 16572 19340 16584
rect 18196 16544 19340 16572
rect 18196 16532 18202 16544
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 19444 16581 19472 16680
rect 19794 16668 19800 16680
rect 19852 16668 19858 16720
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 19576 16612 19748 16640
rect 19576 16600 19582 16612
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19610 16572 19616 16584
rect 19571 16544 19616 16572
rect 19429 16535 19487 16541
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 19720 16581 19748 16612
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 19852 16544 19897 16572
rect 19852 16532 19858 16544
rect 9462 16467 9520 16473
rect 10520 16476 10640 16504
rect 12336 16507 12394 16513
rect 7484 16408 8432 16436
rect 8481 16439 8539 16445
rect 8481 16405 8493 16439
rect 8527 16436 8539 16439
rect 10520 16436 10548 16476
rect 12336 16473 12348 16507
rect 12382 16504 12394 16507
rect 14734 16504 14740 16516
rect 12382 16476 14740 16504
rect 12382 16473 12394 16476
rect 12336 16467 12394 16473
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 16574 16504 16580 16516
rect 16535 16476 16580 16504
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 17402 16504 17408 16516
rect 17363 16476 17408 16504
rect 17402 16464 17408 16476
rect 17460 16464 17466 16516
rect 17773 16507 17831 16513
rect 17773 16473 17785 16507
rect 17819 16504 17831 16507
rect 17819 16476 17908 16504
rect 17819 16473 17831 16476
rect 17773 16467 17831 16473
rect 8527 16408 10548 16436
rect 8527 16405 8539 16408
rect 8481 16399 8539 16405
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 17589 16439 17647 16445
rect 17589 16436 17601 16439
rect 16908 16408 17601 16436
rect 16908 16396 16914 16408
rect 17589 16405 17601 16408
rect 17635 16405 17647 16439
rect 17589 16399 17647 16405
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 17880 16436 17908 16476
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 20073 16507 20131 16513
rect 20073 16504 20085 16507
rect 18104 16476 20085 16504
rect 18104 16464 18110 16476
rect 20073 16473 20085 16476
rect 20119 16473 20131 16507
rect 20073 16467 20131 16473
rect 19518 16436 19524 16448
rect 17736 16408 17781 16436
rect 17880 16408 19524 16436
rect 17736 16396 17742 16408
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 1104 16346 21043 16368
rect 1104 16294 5894 16346
rect 5946 16294 5958 16346
rect 6010 16294 6022 16346
rect 6074 16294 6086 16346
rect 6138 16294 6150 16346
rect 6202 16294 10839 16346
rect 10891 16294 10903 16346
rect 10955 16294 10967 16346
rect 11019 16294 11031 16346
rect 11083 16294 11095 16346
rect 11147 16294 15784 16346
rect 15836 16294 15848 16346
rect 15900 16294 15912 16346
rect 15964 16294 15976 16346
rect 16028 16294 16040 16346
rect 16092 16294 20729 16346
rect 20781 16294 20793 16346
rect 20845 16294 20857 16346
rect 20909 16294 20921 16346
rect 20973 16294 20985 16346
rect 21037 16294 21043 16346
rect 1104 16272 21043 16294
rect 2222 16232 2228 16244
rect 2183 16204 2228 16232
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 2832 16204 2877 16232
rect 2832 16192 2838 16204
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 11882 16232 11888 16244
rect 10652 16204 11888 16232
rect 10652 16192 10658 16204
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 14507 16204 15301 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 17589 16235 17647 16241
rect 17589 16201 17601 16235
rect 17635 16201 17647 16235
rect 19794 16232 19800 16244
rect 19755 16204 19800 16232
rect 17589 16195 17647 16201
rect 3878 16124 3884 16176
rect 3936 16173 3942 16176
rect 3936 16164 3948 16173
rect 12428 16167 12486 16173
rect 3936 16136 3981 16164
rect 4172 16136 6040 16164
rect 3936 16127 3948 16136
rect 3936 16124 3942 16127
rect 1946 16096 1952 16108
rect 1907 16068 1952 16096
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 4172 16105 4200 16136
rect 6012 16108 6040 16136
rect 12428 16133 12440 16167
rect 12474 16164 12486 16167
rect 17604 16164 17632 16195
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 19702 16164 19708 16176
rect 12474 16136 17632 16164
rect 18524 16136 19708 16164
rect 12474 16133 12486 16136
rect 12428 16127 12486 16133
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4157 16059 4215 16065
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 5730 16099 5788 16105
rect 5730 16096 5742 16099
rect 5500 16068 5742 16096
rect 5500 16056 5506 16068
rect 5730 16065 5742 16068
rect 5776 16065 5788 16099
rect 5994 16096 6000 16108
rect 5907 16068 6000 16096
rect 5730 16059 5788 16065
rect 5994 16056 6000 16068
rect 6052 16096 6058 16108
rect 7558 16096 7564 16108
rect 6052 16068 7564 16096
rect 6052 16056 6058 16068
rect 7558 16056 7564 16068
rect 7616 16096 7622 16108
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 7616 16068 8033 16096
rect 7616 16056 7622 16068
rect 8021 16065 8033 16068
rect 8067 16065 8079 16099
rect 8021 16059 8079 16065
rect 8288 16099 8346 16105
rect 8288 16065 8300 16099
rect 8334 16096 8346 16099
rect 9122 16096 9128 16108
rect 8334 16068 9128 16096
rect 8334 16065 8346 16068
rect 8288 16059 8346 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11756 16068 12173 16096
rect 11756 16056 11762 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 14274 16096 14280 16108
rect 14235 16068 14280 16096
rect 12161 16059 12219 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14458 16096 14464 16108
rect 14419 16068 14464 16096
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 15028 16096 15148 16102
rect 15562 16096 15568 16108
rect 15028 16074 15568 16096
rect 15028 16037 15056 16074
rect 15120 16068 15568 16074
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 16117 16099 16175 16105
rect 16117 16096 16129 16099
rect 15672 16068 16129 16096
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 15997 15071 16031
rect 15013 15991 15071 15997
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15252 16000 15297 16028
rect 15252 15988 15258 16000
rect 2746 15932 2912 15960
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 2746 15892 2774 15932
rect 2464 15864 2774 15892
rect 2884 15892 2912 15932
rect 13722 15920 13728 15972
rect 13780 15960 13786 15972
rect 15672 15969 15700 16068
rect 16117 16065 16129 16068
rect 16163 16065 16175 16099
rect 16298 16096 16304 16108
rect 16259 16068 16304 16096
rect 16117 16059 16175 16065
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 16850 16096 16856 16108
rect 16811 16068 16856 16096
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 16942 16056 16948 16108
rect 17000 16096 17006 16108
rect 17129 16099 17187 16105
rect 17000 16068 17045 16096
rect 17000 16056 17006 16068
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 17586 16096 17592 16108
rect 17175 16068 17592 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18524 16105 18552 16136
rect 18325 16099 18383 16105
rect 18325 16096 18337 16099
rect 17736 16068 18337 16096
rect 17736 16056 17742 16068
rect 18325 16065 18337 16068
rect 18371 16065 18383 16099
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18325 16059 18383 16065
rect 18432 16068 18521 16096
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 17494 16028 17500 16040
rect 16632 16000 17500 16028
rect 16632 15988 16638 16000
rect 17494 15988 17500 16000
rect 17552 16028 17558 16040
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 17552 16000 17877 16028
rect 17552 15988 17558 16000
rect 17865 15997 17877 16000
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 15657 15963 15715 15969
rect 13780 15932 15240 15960
rect 13780 15920 13786 15932
rect 4617 15895 4675 15901
rect 4617 15892 4629 15895
rect 2884 15864 4629 15892
rect 2464 15852 2470 15864
rect 4617 15861 4629 15864
rect 4663 15861 4675 15895
rect 4617 15855 4675 15861
rect 9401 15895 9459 15901
rect 9401 15861 9413 15895
rect 9447 15892 9459 15895
rect 9490 15892 9496 15904
rect 9447 15864 9496 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 13541 15895 13599 15901
rect 13541 15861 13553 15895
rect 13587 15892 13599 15895
rect 15102 15892 15108 15904
rect 13587 15864 15108 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 15212 15892 15240 15932
rect 15657 15929 15669 15963
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 16758 15920 16764 15972
rect 16816 15960 16822 15972
rect 17129 15963 17187 15969
rect 17129 15960 17141 15963
rect 16816 15932 17141 15960
rect 16816 15920 16822 15932
rect 17129 15929 17141 15932
rect 17175 15929 17187 15963
rect 17129 15923 17187 15929
rect 17681 15963 17739 15969
rect 17681 15929 17693 15963
rect 17727 15960 17739 15963
rect 18325 15963 18383 15969
rect 18325 15960 18337 15963
rect 17727 15932 18337 15960
rect 17727 15929 17739 15932
rect 17681 15923 17739 15929
rect 18325 15929 18337 15932
rect 18371 15929 18383 15963
rect 18325 15923 18383 15929
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 15212 15864 16129 15892
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 18432 15892 18460 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18509 16059 18567 16065
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 19518 16096 19524 16108
rect 18647 16068 19524 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 19518 16056 19524 16068
rect 19576 16056 19582 16108
rect 19628 16105 19656 16136
rect 19702 16124 19708 16136
rect 19760 16124 19766 16176
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19426 16028 19432 16040
rect 19387 16000 19432 16028
rect 19426 15988 19432 16000
rect 19484 15988 19490 16040
rect 17368 15864 18460 15892
rect 17368 15852 17374 15864
rect 1104 15802 20884 15824
rect 1104 15750 3422 15802
rect 3474 15750 3486 15802
rect 3538 15750 3550 15802
rect 3602 15750 3614 15802
rect 3666 15750 3678 15802
rect 3730 15750 8367 15802
rect 8419 15750 8431 15802
rect 8483 15750 8495 15802
rect 8547 15750 8559 15802
rect 8611 15750 8623 15802
rect 8675 15750 13312 15802
rect 13364 15750 13376 15802
rect 13428 15750 13440 15802
rect 13492 15750 13504 15802
rect 13556 15750 13568 15802
rect 13620 15750 18257 15802
rect 18309 15750 18321 15802
rect 18373 15750 18385 15802
rect 18437 15750 18449 15802
rect 18501 15750 18513 15802
rect 18565 15750 20884 15802
rect 1104 15728 20884 15750
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5721 15691 5779 15697
rect 5721 15688 5733 15691
rect 5684 15660 5733 15688
rect 5684 15648 5690 15660
rect 5721 15657 5733 15660
rect 5767 15688 5779 15691
rect 5994 15688 6000 15700
rect 5767 15660 6000 15688
rect 5767 15657 5779 15660
rect 5721 15651 5779 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 15381 15691 15439 15697
rect 15381 15657 15393 15691
rect 15427 15688 15439 15691
rect 17405 15691 17463 15697
rect 17405 15688 17417 15691
rect 15427 15660 17417 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 17405 15657 17417 15660
rect 17451 15657 17463 15691
rect 17586 15688 17592 15700
rect 17547 15660 17592 15688
rect 17405 15651 17463 15657
rect 1949 15623 2007 15629
rect 1949 15589 1961 15623
rect 1995 15620 2007 15623
rect 2314 15620 2320 15632
rect 1995 15592 2320 15620
rect 1995 15589 2007 15592
rect 1949 15583 2007 15589
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 14458 15580 14464 15632
rect 14516 15620 14522 15632
rect 17034 15620 17040 15632
rect 14516 15592 17040 15620
rect 14516 15580 14522 15592
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 17420 15620 17448 15651
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 17862 15648 17868 15700
rect 17920 15688 17926 15700
rect 19426 15688 19432 15700
rect 17920 15660 19432 15688
rect 17920 15648 17926 15660
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 17678 15620 17684 15632
rect 17420 15592 17684 15620
rect 17678 15580 17684 15592
rect 17736 15580 17742 15632
rect 15010 15552 15016 15564
rect 14923 15524 15016 15552
rect 15010 15512 15016 15524
rect 15068 15552 15074 15564
rect 15286 15552 15292 15564
rect 15068 15524 15292 15552
rect 15068 15512 15074 15524
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 17862 15552 17868 15564
rect 17000 15524 17868 15552
rect 17000 15512 17006 15524
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15484 2283 15487
rect 2406 15484 2412 15496
rect 2271 15456 2412 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 15102 15444 15108 15496
rect 15160 15484 15166 15496
rect 15197 15487 15255 15493
rect 15197 15484 15209 15487
rect 15160 15456 15209 15484
rect 15160 15444 15166 15456
rect 15197 15453 15209 15456
rect 15243 15453 15255 15487
rect 15197 15447 15255 15453
rect 1949 15419 2007 15425
rect 1949 15385 1961 15419
rect 1995 15416 2007 15419
rect 2498 15416 2504 15428
rect 1995 15388 2504 15416
rect 1995 15385 2007 15388
rect 1949 15379 2007 15385
rect 2498 15376 2504 15388
rect 2556 15376 2562 15428
rect 7009 15419 7067 15425
rect 7009 15385 7021 15419
rect 7055 15416 7067 15419
rect 9582 15416 9588 15428
rect 7055 15388 9588 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 9582 15376 9588 15388
rect 9640 15416 9646 15428
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 9640 15388 10425 15416
rect 9640 15376 9646 15388
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 10413 15379 10471 15385
rect 13630 15376 13636 15428
rect 13688 15416 13694 15428
rect 16666 15416 16672 15428
rect 13688 15388 16672 15416
rect 13688 15376 13694 15388
rect 16666 15376 16672 15388
rect 16724 15416 16730 15428
rect 17221 15419 17279 15425
rect 17221 15416 17233 15419
rect 16724 15388 17233 15416
rect 16724 15376 16730 15388
rect 17221 15385 17233 15388
rect 17267 15416 17279 15419
rect 17310 15416 17316 15428
rect 17267 15388 17316 15416
rect 17267 15385 17279 15388
rect 17221 15379 17279 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17437 15419 17495 15425
rect 17437 15385 17449 15419
rect 17483 15416 17495 15419
rect 19518 15416 19524 15428
rect 17483 15388 19524 15416
rect 17483 15385 17495 15388
rect 17437 15379 17495 15385
rect 19518 15376 19524 15388
rect 19576 15376 19582 15428
rect 2038 15308 2044 15360
rect 2096 15348 2102 15360
rect 2133 15351 2191 15357
rect 2133 15348 2145 15351
rect 2096 15320 2145 15348
rect 2096 15308 2102 15320
rect 2133 15317 2145 15320
rect 2179 15317 2191 15351
rect 2133 15311 2191 15317
rect 1104 15258 21043 15280
rect 1104 15206 5894 15258
rect 5946 15206 5958 15258
rect 6010 15206 6022 15258
rect 6074 15206 6086 15258
rect 6138 15206 6150 15258
rect 6202 15206 10839 15258
rect 10891 15206 10903 15258
rect 10955 15206 10967 15258
rect 11019 15206 11031 15258
rect 11083 15206 11095 15258
rect 11147 15206 15784 15258
rect 15836 15206 15848 15258
rect 15900 15206 15912 15258
rect 15964 15206 15976 15258
rect 16028 15206 16040 15258
rect 16092 15206 20729 15258
rect 20781 15206 20793 15258
rect 20845 15206 20857 15258
rect 20909 15206 20921 15258
rect 20973 15206 20985 15258
rect 21037 15206 21043 15258
rect 1104 15184 21043 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 4154 15144 4160 15156
rect 2547 15116 4160 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 9582 15144 9588 15156
rect 9543 15116 9588 15144
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 8294 15076 8300 15088
rect 8255 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15036 8358 15088
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 11698 15008 11704 15020
rect 9272 14980 11704 15008
rect 9272 14968 9278 14980
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 11968 15011 12026 15017
rect 11968 14977 11980 15011
rect 12014 15008 12026 15011
rect 16942 15008 16948 15020
rect 12014 14980 16948 15008
rect 12014 14977 12026 14980
rect 11968 14971 12026 14977
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 19518 15008 19524 15020
rect 19479 14980 19524 15008
rect 19518 14968 19524 14980
rect 19576 14968 19582 15020
rect 1946 14900 1952 14952
rect 2004 14940 2010 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 2004 14912 2053 14940
rect 2004 14900 2010 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14940 2191 14943
rect 2406 14940 2412 14952
rect 2179 14912 2412 14940
rect 2179 14909 2191 14912
rect 2133 14903 2191 14909
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 16850 14940 16856 14952
rect 14967 14912 16856 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 13081 14875 13139 14881
rect 13081 14841 13093 14875
rect 13127 14872 13139 14875
rect 14936 14872 14964 14903
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 13127 14844 14964 14872
rect 15289 14875 15347 14881
rect 13127 14841 13139 14844
rect 13081 14835 13139 14841
rect 15289 14841 15301 14875
rect 15335 14872 15347 14875
rect 15470 14872 15476 14884
rect 15335 14844 15476 14872
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 15470 14832 15476 14844
rect 15528 14832 15534 14884
rect 15378 14804 15384 14816
rect 15339 14776 15384 14804
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 19613 14807 19671 14813
rect 19613 14773 19625 14807
rect 19659 14804 19671 14807
rect 19702 14804 19708 14816
rect 19659 14776 19708 14804
rect 19659 14773 19671 14776
rect 19613 14767 19671 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 1104 14714 20884 14736
rect 1104 14662 3422 14714
rect 3474 14662 3486 14714
rect 3538 14662 3550 14714
rect 3602 14662 3614 14714
rect 3666 14662 3678 14714
rect 3730 14662 8367 14714
rect 8419 14662 8431 14714
rect 8483 14662 8495 14714
rect 8547 14662 8559 14714
rect 8611 14662 8623 14714
rect 8675 14662 13312 14714
rect 13364 14662 13376 14714
rect 13428 14662 13440 14714
rect 13492 14662 13504 14714
rect 13556 14662 13568 14714
rect 13620 14662 18257 14714
rect 18309 14662 18321 14714
rect 18373 14662 18385 14714
rect 18437 14662 18449 14714
rect 18501 14662 18513 14714
rect 18565 14662 20884 14714
rect 1104 14640 20884 14662
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 15470 14600 15476 14612
rect 11195 14572 15476 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 16816 14572 16865 14600
rect 16816 14560 16822 14572
rect 16853 14569 16865 14572
rect 16899 14569 16911 14603
rect 16853 14563 16911 14569
rect 16945 14603 17003 14609
rect 16945 14569 16957 14603
rect 16991 14600 17003 14603
rect 17126 14600 17132 14612
rect 16991 14572 17132 14600
rect 16991 14569 17003 14572
rect 16945 14563 17003 14569
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 19981 14603 20039 14609
rect 19981 14600 19993 14603
rect 19576 14572 19993 14600
rect 19576 14560 19582 14572
rect 19981 14569 19993 14572
rect 20027 14569 20039 14603
rect 19981 14563 20039 14569
rect 14918 14492 14924 14544
rect 14976 14532 14982 14544
rect 15105 14535 15163 14541
rect 15105 14532 15117 14535
rect 14976 14504 15117 14532
rect 14976 14492 14982 14504
rect 15105 14501 15117 14504
rect 15151 14501 15163 14535
rect 15105 14495 15163 14501
rect 15197 14535 15255 14541
rect 15197 14501 15209 14535
rect 15243 14532 15255 14535
rect 15378 14532 15384 14544
rect 15243 14504 15384 14532
rect 15243 14501 15255 14504
rect 15197 14495 15255 14501
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 18414 14532 18420 14544
rect 16500 14504 18420 14532
rect 1946 14424 1952 14476
rect 2004 14464 2010 14476
rect 3973 14467 4031 14473
rect 3973 14464 3985 14467
rect 2004 14436 3985 14464
rect 2004 14424 2010 14436
rect 3973 14433 3985 14436
rect 4019 14433 4031 14467
rect 5626 14464 5632 14476
rect 5587 14436 5632 14464
rect 3973 14427 4031 14433
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9585 14467 9643 14473
rect 9585 14464 9597 14467
rect 9272 14436 9597 14464
rect 9272 14424 9278 14436
rect 9585 14433 9597 14436
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 16500 14464 16528 14504
rect 18414 14492 18420 14504
rect 18472 14532 18478 14544
rect 19150 14532 19156 14544
rect 18472 14504 19156 14532
rect 18472 14492 18478 14504
rect 19150 14492 19156 14504
rect 19208 14532 19214 14544
rect 19429 14535 19487 14541
rect 19429 14532 19441 14535
rect 19208 14504 19441 14532
rect 19208 14492 19214 14504
rect 19429 14501 19441 14504
rect 19475 14501 19487 14535
rect 19429 14495 19487 14501
rect 14700 14436 16528 14464
rect 16592 14436 18000 14464
rect 14700 14424 14706 14436
rect 16592 14408 16620 14436
rect 2130 14396 2136 14408
rect 2043 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 5258 14396 5264 14408
rect 2271 14368 5264 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 5258 14356 5264 14368
rect 5316 14356 5322 14408
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 7193 14399 7251 14405
rect 5408 14368 5453 14396
rect 5408 14356 5414 14368
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 7926 14396 7932 14408
rect 7239 14368 7932 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 15010 14396 15016 14408
rect 14971 14368 15016 14396
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 16574 14396 16580 14408
rect 16535 14368 16580 14396
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16666 14356 16672 14408
rect 16724 14396 16730 14408
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16724 14368 16773 14396
rect 16724 14356 16730 14368
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17770 14396 17776 14408
rect 17092 14368 17137 14396
rect 17731 14368 17776 14396
rect 17092 14356 17098 14368
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 17972 14405 18000 14436
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 18748 14436 19932 14464
rect 18748 14424 18754 14436
rect 17957 14399 18015 14405
rect 17957 14365 17969 14399
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 18598 14356 18604 14408
rect 18656 14396 18662 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 18656 14368 19809 14396
rect 18656 14356 18662 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 2148 14328 2176 14356
rect 2314 14328 2320 14340
rect 2148 14300 2320 14328
rect 2314 14288 2320 14300
rect 2372 14288 2378 14340
rect 7460 14331 7518 14337
rect 7460 14297 7472 14331
rect 7506 14328 7518 14331
rect 7558 14328 7564 14340
rect 7506 14300 7564 14328
rect 7506 14297 7518 14300
rect 7460 14291 7518 14297
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 12428 14331 12486 14337
rect 12428 14297 12440 14331
rect 12474 14328 12486 14331
rect 19334 14328 19340 14340
rect 12474 14300 19340 14328
rect 12474 14297 12486 14300
rect 12428 14291 12486 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 19705 14331 19763 14337
rect 19705 14297 19717 14331
rect 19751 14328 19763 14331
rect 19904 14328 19932 14436
rect 19751 14300 19932 14328
rect 19751 14297 19763 14300
rect 19705 14291 19763 14297
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 8573 14263 8631 14269
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 8754 14260 8760 14272
rect 8619 14232 8760 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 13541 14263 13599 14269
rect 13541 14229 13553 14263
rect 13587 14260 13599 14263
rect 14642 14260 14648 14272
rect 13587 14232 14648 14260
rect 13587 14229 13599 14232
rect 13541 14223 13599 14229
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 14826 14260 14832 14272
rect 14787 14232 14832 14260
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 16114 14260 16120 14272
rect 15252 14232 16120 14260
rect 15252 14220 15258 14232
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17310 14260 17316 14272
rect 17271 14232 17316 14260
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 19518 14260 19524 14272
rect 18187 14232 19524 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 19518 14220 19524 14232
rect 19576 14260 19582 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 19576 14232 19625 14260
rect 19576 14220 19582 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 1104 14170 21043 14192
rect 1104 14118 5894 14170
rect 5946 14118 5958 14170
rect 6010 14118 6022 14170
rect 6074 14118 6086 14170
rect 6138 14118 6150 14170
rect 6202 14118 10839 14170
rect 10891 14118 10903 14170
rect 10955 14118 10967 14170
rect 11019 14118 11031 14170
rect 11083 14118 11095 14170
rect 11147 14118 15784 14170
rect 15836 14118 15848 14170
rect 15900 14118 15912 14170
rect 15964 14118 15976 14170
rect 16028 14118 16040 14170
rect 16092 14118 20729 14170
rect 20781 14118 20793 14170
rect 20845 14118 20857 14170
rect 20909 14118 20921 14170
rect 20973 14118 20985 14170
rect 21037 14118 21043 14170
rect 1104 14096 21043 14118
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 9033 14059 9091 14065
rect 2464 14028 5304 14056
rect 2464 14016 2470 14028
rect 2869 13991 2927 13997
rect 2869 13988 2881 13991
rect 2746 13960 2881 13988
rect 1854 13880 1860 13932
rect 1912 13920 1918 13932
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 1912 13892 2237 13920
rect 1912 13880 1918 13892
rect 2225 13889 2237 13892
rect 2271 13889 2283 13923
rect 2225 13883 2283 13889
rect 2406 13880 2412 13932
rect 2464 13920 2470 13932
rect 2746 13920 2774 13960
rect 2869 13957 2881 13960
rect 2915 13957 2927 13991
rect 5276 13988 5304 14028
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 13541 14059 13599 14065
rect 9079 14028 12388 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 7662 13991 7720 13997
rect 7662 13988 7674 13991
rect 2869 13951 2927 13957
rect 2976 13960 3832 13988
rect 5276 13960 7674 13988
rect 2464 13892 2774 13920
rect 2464 13880 2470 13892
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13852 2099 13855
rect 2130 13852 2136 13864
rect 2087 13824 2136 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 2130 13812 2136 13824
rect 2188 13852 2194 13864
rect 2976 13852 3004 13960
rect 3053 13923 3111 13929
rect 3053 13889 3065 13923
rect 3099 13920 3111 13923
rect 3142 13920 3148 13932
rect 3099 13892 3148 13920
rect 3099 13889 3111 13892
rect 3053 13883 3111 13889
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13920 3295 13923
rect 3602 13920 3608 13932
rect 3283 13892 3608 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 2188 13824 3004 13852
rect 2188 13812 2194 13824
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13784 2467 13787
rect 2866 13784 2872 13796
rect 2455 13756 2872 13784
rect 2455 13753 2467 13756
rect 2409 13747 2467 13753
rect 2866 13744 2872 13756
rect 2924 13744 2930 13796
rect 3804 13716 3832 13960
rect 7662 13957 7674 13960
rect 7708 13957 7720 13991
rect 7662 13951 7720 13957
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4028 13892 5089 13920
rect 4028 13880 4034 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 7926 13920 7932 13932
rect 7887 13892 7932 13920
rect 5077 13883 5135 13889
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 10134 13920 10140 13932
rect 10192 13929 10198 13932
rect 10104 13892 10140 13920
rect 10134 13880 10140 13892
rect 10192 13883 10204 13929
rect 12360 13920 12388 14028
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 16574 14056 16580 14068
rect 13587 14028 16580 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 16942 14056 16948 14068
rect 16903 14028 16948 14056
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 18785 14059 18843 14065
rect 18785 14025 18797 14059
rect 18831 14025 18843 14059
rect 18785 14019 18843 14025
rect 12428 13991 12486 13997
rect 12428 13957 12440 13991
rect 12474 13988 12486 13991
rect 17126 13988 17132 14000
rect 12474 13960 15884 13988
rect 17087 13960 17132 13988
rect 12474 13957 12486 13960
rect 12428 13951 12486 13957
rect 14918 13920 14924 13932
rect 12360 13892 14320 13920
rect 14879 13892 14924 13920
rect 10192 13880 10198 13883
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 5534 13852 5540 13864
rect 5399 13824 5540 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 11698 13852 11704 13864
rect 10459 13824 11704 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 11698 13812 11704 13824
rect 11756 13852 11762 13864
rect 12158 13852 12164 13864
rect 11756 13824 12164 13852
rect 11756 13812 11762 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 14292 13852 14320 13892
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 15344 13892 15393 13920
rect 15344 13880 15350 13892
rect 15381 13889 15393 13892
rect 15427 13920 15439 13923
rect 15856 13920 15884 13960
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 18414 13988 18420 14000
rect 18375 13960 18420 13988
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 18598 13948 18604 14000
rect 18656 13997 18662 14000
rect 18656 13991 18675 13997
rect 18663 13957 18675 13991
rect 18800 13988 18828 14019
rect 19978 13988 19984 14000
rect 18800 13960 19984 13988
rect 18656 13951 18675 13957
rect 18656 13948 18662 13951
rect 19518 13920 19524 13932
rect 15427 13892 15792 13920
rect 15856 13892 19288 13920
rect 19479 13892 19524 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 15194 13852 15200 13864
rect 14292 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 15654 13852 15660 13864
rect 15615 13824 15660 13852
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15764 13852 15792 13892
rect 19260 13861 19288 13892
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 19628 13929 19656 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 19702 13880 19708 13932
rect 19760 13920 19766 13932
rect 19889 13923 19947 13929
rect 19760 13892 19805 13920
rect 19760 13880 19766 13892
rect 19889 13889 19901 13923
rect 19935 13889 19947 13923
rect 19889 13883 19947 13889
rect 17497 13855 17555 13861
rect 15764 13824 16620 13852
rect 3970 13784 3976 13796
rect 3931 13756 3976 13784
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 14274 13744 14280 13796
rect 14332 13784 14338 13796
rect 15105 13787 15163 13793
rect 15105 13784 15117 13787
rect 14332 13756 15117 13784
rect 14332 13744 14338 13756
rect 15105 13753 15117 13756
rect 15151 13753 15163 13787
rect 15286 13784 15292 13796
rect 15247 13756 15292 13784
rect 15105 13747 15163 13753
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 16592 13784 16620 13824
rect 17497 13821 17509 13855
rect 17543 13852 17555 13855
rect 19245 13855 19303 13861
rect 17543 13824 18644 13852
rect 17543 13821 17555 13824
rect 17497 13815 17555 13821
rect 17770 13784 17776 13796
rect 16592 13756 17776 13784
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 3804 13688 6561 13716
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6549 13679 6607 13685
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 17129 13719 17187 13725
rect 15252 13688 15297 13716
rect 15252 13676 15258 13688
rect 17129 13685 17141 13719
rect 17175 13716 17187 13719
rect 17218 13716 17224 13728
rect 17175 13688 17224 13716
rect 17175 13685 17187 13688
rect 17129 13679 17187 13685
rect 17218 13676 17224 13688
rect 17276 13676 17282 13728
rect 18616 13725 18644 13824
rect 19245 13821 19257 13855
rect 19291 13821 19303 13855
rect 19904 13852 19932 13883
rect 19245 13815 19303 13821
rect 19720 13824 19932 13852
rect 19720 13796 19748 13824
rect 19702 13744 19708 13796
rect 19760 13744 19766 13796
rect 18601 13719 18659 13725
rect 18601 13685 18613 13719
rect 18647 13716 18659 13719
rect 18690 13716 18696 13728
rect 18647 13688 18696 13716
rect 18647 13685 18659 13688
rect 18601 13679 18659 13685
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 1104 13626 20884 13648
rect 1104 13574 3422 13626
rect 3474 13574 3486 13626
rect 3538 13574 3550 13626
rect 3602 13574 3614 13626
rect 3666 13574 3678 13626
rect 3730 13574 8367 13626
rect 8419 13574 8431 13626
rect 8483 13574 8495 13626
rect 8547 13574 8559 13626
rect 8611 13574 8623 13626
rect 8675 13574 13312 13626
rect 13364 13574 13376 13626
rect 13428 13574 13440 13626
rect 13492 13574 13504 13626
rect 13556 13574 13568 13626
rect 13620 13574 18257 13626
rect 18309 13574 18321 13626
rect 18373 13574 18385 13626
rect 18437 13574 18449 13626
rect 18501 13574 18513 13626
rect 18565 13574 20884 13626
rect 1104 13552 20884 13574
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 5350 13512 5356 13524
rect 2363 13484 5356 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 17126 13472 17132 13524
rect 17184 13512 17190 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 17184 13484 17325 13512
rect 17184 13472 17190 13484
rect 17313 13481 17325 13484
rect 17359 13481 17371 13515
rect 17313 13475 17371 13481
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 19392 13484 19441 13512
rect 19392 13472 19398 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 19610 13512 19616 13524
rect 19571 13484 19616 13512
rect 19429 13475 19487 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 2866 13404 2872 13456
rect 2924 13444 2930 13456
rect 4246 13444 4252 13456
rect 2924 13416 4252 13444
rect 2924 13404 2930 13416
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 19978 13444 19984 13456
rect 19939 13416 19984 13444
rect 19978 13404 19984 13416
rect 20036 13404 20042 13456
rect 3970 13376 3976 13388
rect 2056 13348 3976 13376
rect 2056 13320 2084 13348
rect 3970 13336 3976 13348
rect 4028 13336 4034 13388
rect 2038 13308 2044 13320
rect 1999 13280 2044 13308
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2314 13308 2320 13320
rect 2179 13280 2320 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5592 13280 6009 13308
rect 5592 13268 5598 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 16850 13308 16856 13320
rect 16811 13280 16856 13308
rect 5997 13271 6055 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13308 17187 13311
rect 17954 13308 17960 13320
rect 17175 13280 17960 13308
rect 17175 13277 17187 13280
rect 17129 13271 17187 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 6264 13243 6322 13249
rect 6264 13209 6276 13243
rect 6310 13240 6322 13243
rect 6454 13240 6460 13252
rect 6310 13212 6460 13240
rect 6310 13209 6322 13212
rect 6264 13203 6322 13209
rect 6454 13200 6460 13212
rect 6512 13200 6518 13252
rect 7377 13175 7435 13181
rect 7377 13141 7389 13175
rect 7423 13172 7435 13175
rect 7466 13172 7472 13184
rect 7423 13144 7472 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 16945 13175 17003 13181
rect 16945 13141 16957 13175
rect 16991 13172 17003 13175
rect 17770 13172 17776 13184
rect 16991 13144 17776 13172
rect 16991 13141 17003 13144
rect 16945 13135 17003 13141
rect 17770 13132 17776 13144
rect 17828 13172 17834 13184
rect 19242 13172 19248 13184
rect 17828 13144 19248 13172
rect 17828 13132 17834 13144
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 19613 13175 19671 13181
rect 19613 13141 19625 13175
rect 19659 13172 19671 13175
rect 19702 13172 19708 13184
rect 19659 13144 19708 13172
rect 19659 13141 19671 13144
rect 19613 13135 19671 13141
rect 19702 13132 19708 13144
rect 19760 13132 19766 13184
rect 1104 13082 21043 13104
rect 1104 13030 5894 13082
rect 5946 13030 5958 13082
rect 6010 13030 6022 13082
rect 6074 13030 6086 13082
rect 6138 13030 6150 13082
rect 6202 13030 10839 13082
rect 10891 13030 10903 13082
rect 10955 13030 10967 13082
rect 11019 13030 11031 13082
rect 11083 13030 11095 13082
rect 11147 13030 15784 13082
rect 15836 13030 15848 13082
rect 15900 13030 15912 13082
rect 15964 13030 15976 13082
rect 16028 13030 16040 13082
rect 16092 13030 20729 13082
rect 20781 13030 20793 13082
rect 20845 13030 20857 13082
rect 20909 13030 20921 13082
rect 20973 13030 20985 13082
rect 21037 13030 21043 13082
rect 1104 13008 21043 13030
rect 19610 12968 19616 12980
rect 19571 12940 19616 12968
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 1762 12860 1768 12912
rect 1820 12900 1826 12912
rect 1857 12903 1915 12909
rect 1857 12900 1869 12903
rect 1820 12872 1869 12900
rect 1820 12860 1826 12872
rect 1857 12869 1869 12872
rect 1903 12869 1915 12903
rect 1857 12863 1915 12869
rect 1946 12860 1952 12912
rect 2004 12900 2010 12912
rect 2041 12903 2099 12909
rect 2041 12900 2053 12903
rect 2004 12872 2053 12900
rect 2004 12860 2010 12872
rect 2041 12869 2053 12872
rect 2087 12900 2099 12903
rect 2498 12900 2504 12912
rect 2087 12872 2504 12900
rect 2087 12869 2099 12872
rect 2041 12863 2099 12869
rect 2498 12860 2504 12872
rect 2556 12860 2562 12912
rect 5534 12900 5540 12912
rect 4172 12872 5540 12900
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 4172 12841 4200 12872
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 17218 12900 17224 12912
rect 17131 12872 17224 12900
rect 17218 12860 17224 12872
rect 17276 12900 17282 12912
rect 17770 12900 17776 12912
rect 17276 12872 17776 12900
rect 17276 12860 17282 12872
rect 17770 12860 17776 12872
rect 17828 12860 17834 12912
rect 18693 12903 18751 12909
rect 18693 12869 18705 12903
rect 18739 12900 18751 12903
rect 19334 12900 19340 12912
rect 18739 12872 19340 12900
rect 18739 12869 18751 12872
rect 18693 12863 18751 12869
rect 19334 12860 19340 12872
rect 19392 12900 19398 12912
rect 19392 12872 19472 12900
rect 19392 12860 19398 12872
rect 4430 12841 4436 12844
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 4424 12795 4436 12841
rect 4488 12832 4494 12844
rect 4488 12804 4524 12832
rect 4430 12792 4436 12795
rect 4488 12792 4494 12804
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7984 12804 8217 12832
rect 7984 12792 7990 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 8205 12795 8263 12801
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 11968 12835 12026 12841
rect 11968 12801 11980 12835
rect 12014 12832 12026 12835
rect 18509 12835 18567 12841
rect 12014 12804 18092 12832
rect 12014 12801 12026 12804
rect 11968 12795 12026 12801
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 8846 12764 8852 12776
rect 8527 12736 8852 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 17589 12699 17647 12705
rect 17589 12665 17601 12699
rect 17635 12696 17647 12699
rect 17954 12696 17960 12708
rect 17635 12668 17960 12696
rect 17635 12665 17647 12668
rect 17589 12659 17647 12665
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 18064 12696 18092 12804
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 18598 12832 18604 12844
rect 18555 12804 18604 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 19150 12832 19156 12844
rect 19111 12804 19156 12832
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19242 12792 19248 12844
rect 19300 12832 19306 12844
rect 19444 12841 19472 12872
rect 19429 12835 19487 12841
rect 19300 12804 19393 12832
rect 19300 12792 19306 12804
rect 19429 12801 19441 12835
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 18690 12764 18696 12776
rect 18371 12736 18696 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 19260 12764 19288 12792
rect 19610 12764 19616 12776
rect 19260 12736 19616 12764
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19978 12696 19984 12708
rect 18064 12668 19984 12696
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 5537 12631 5595 12637
rect 5537 12597 5549 12631
rect 5583 12628 5595 12631
rect 5626 12628 5632 12640
rect 5583 12600 5632 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 11238 12628 11244 12640
rect 9815 12600 11244 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 13081 12631 13139 12637
rect 13081 12597 13093 12631
rect 13127 12628 13139 12631
rect 14734 12628 14740 12640
rect 13127 12600 14740 12628
rect 13127 12597 13139 12600
rect 13081 12591 13139 12597
rect 14734 12588 14740 12600
rect 14792 12588 14798 12640
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 15436 12600 17049 12628
rect 15436 12588 15442 12600
rect 17037 12597 17049 12600
rect 17083 12597 17095 12631
rect 17037 12591 17095 12597
rect 17221 12631 17279 12637
rect 17221 12597 17233 12631
rect 17267 12628 17279 12631
rect 18690 12628 18696 12640
rect 17267 12600 18696 12628
rect 17267 12597 17279 12600
rect 17221 12591 17279 12597
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 1104 12538 20884 12560
rect 1104 12486 3422 12538
rect 3474 12486 3486 12538
rect 3538 12486 3550 12538
rect 3602 12486 3614 12538
rect 3666 12486 3678 12538
rect 3730 12486 8367 12538
rect 8419 12486 8431 12538
rect 8483 12486 8495 12538
rect 8547 12486 8559 12538
rect 8611 12486 8623 12538
rect 8675 12486 13312 12538
rect 13364 12486 13376 12538
rect 13428 12486 13440 12538
rect 13492 12486 13504 12538
rect 13556 12486 13568 12538
rect 13620 12486 18257 12538
rect 18309 12486 18321 12538
rect 18373 12486 18385 12538
rect 18437 12486 18449 12538
rect 18501 12486 18513 12538
rect 18565 12486 20884 12538
rect 1104 12464 20884 12486
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 15194 12424 15200 12436
rect 11940 12396 13032 12424
rect 15155 12396 15200 12424
rect 11940 12384 11946 12396
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 1854 12288 1860 12300
rect 1719 12260 1860 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 1854 12248 1860 12260
rect 1912 12288 1918 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 1912 12260 3985 12288
rect 1912 12248 1918 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1765 12183 1823 12189
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 1780 12152 1808 12183
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 2179 12192 5365 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5592 12192 5641 12220
rect 5592 12180 5598 12192
rect 5629 12189 5641 12192
rect 5675 12220 5687 12223
rect 6546 12220 6552 12232
rect 5675 12192 6552 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 6546 12180 6552 12192
rect 6604 12220 6610 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6604 12192 7205 12220
rect 6604 12180 6610 12192
rect 7193 12189 7205 12192
rect 7239 12220 7251 12223
rect 7926 12220 7932 12232
rect 7239 12192 7932 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 11698 12220 11704 12232
rect 9631 12192 11704 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 13004 12220 13032 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 15657 12427 15715 12433
rect 15657 12424 15669 12427
rect 15344 12396 15669 12424
rect 15344 12384 15350 12396
rect 15657 12393 15669 12396
rect 15703 12393 15715 12427
rect 17954 12424 17960 12436
rect 17915 12396 17960 12424
rect 15657 12387 15715 12393
rect 17954 12384 17960 12396
rect 18012 12384 18018 12436
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19702 12384 19708 12436
rect 19760 12424 19766 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19760 12396 19809 12424
rect 19760 12384 19766 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19797 12387 19855 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 13081 12359 13139 12365
rect 13081 12325 13093 12359
rect 13127 12356 13139 12359
rect 13127 12328 15424 12356
rect 13127 12325 13139 12328
rect 13081 12319 13139 12325
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 13872 12260 14749 12288
rect 13872 12248 13878 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 15396 12288 15424 12328
rect 15562 12316 15568 12368
rect 15620 12356 15626 12368
rect 15749 12359 15807 12365
rect 15749 12356 15761 12359
rect 15620 12328 15761 12356
rect 15620 12316 15626 12328
rect 15749 12325 15761 12328
rect 15795 12325 15807 12359
rect 15749 12319 15807 12325
rect 16206 12316 16212 12368
rect 16264 12356 16270 12368
rect 18046 12356 18052 12368
rect 16264 12328 18052 12356
rect 16264 12316 16270 12328
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 15396 12260 17141 12288
rect 14737 12251 14795 12257
rect 17129 12257 17141 12260
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 13004 12192 14841 12220
rect 14829 12189 14841 12192
rect 14875 12220 14887 12223
rect 16114 12220 16120 12232
rect 14875 12192 15976 12220
rect 16075 12192 16120 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 7438 12155 7496 12161
rect 7438 12152 7450 12155
rect 1728 12124 1808 12152
rect 5828 12124 7450 12152
rect 1728 12112 1734 12124
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 5828 12084 5856 12124
rect 7438 12121 7450 12124
rect 7484 12121 7496 12155
rect 7438 12115 7496 12121
rect 9852 12155 9910 12161
rect 9852 12121 9864 12155
rect 9898 12152 9910 12155
rect 10594 12152 10600 12164
rect 9898 12124 10600 12152
rect 9898 12121 9910 12124
rect 9852 12115 9910 12121
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 11968 12155 12026 12161
rect 11968 12121 11980 12155
rect 12014 12152 12026 12155
rect 12014 12124 12434 12152
rect 12014 12121 12026 12124
rect 11968 12115 12026 12121
rect 4304 12056 5856 12084
rect 8573 12087 8631 12093
rect 4304 12044 4310 12056
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 9674 12084 9680 12096
rect 8619 12056 9680 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 10965 12087 11023 12093
rect 10965 12053 10977 12087
rect 11011 12084 11023 12087
rect 11606 12084 11612 12096
rect 11011 12056 11612 12084
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12406 12084 12434 12124
rect 14734 12112 14740 12164
rect 14792 12152 14798 12164
rect 15102 12152 15108 12164
rect 14792 12124 15108 12152
rect 14792 12112 14798 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15948 12152 15976 12192
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 17420 12229 17448 12328
rect 18046 12316 18052 12328
rect 18104 12316 18110 12368
rect 19334 12316 19340 12368
rect 19392 12356 19398 12368
rect 19429 12359 19487 12365
rect 19429 12356 19441 12359
rect 19392 12328 19441 12356
rect 19392 12316 19398 12328
rect 19429 12325 19441 12328
rect 19475 12325 19487 12359
rect 19429 12319 19487 12325
rect 17972 12260 18828 12288
rect 17972 12232 18000 12260
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 17954 12220 17960 12232
rect 17867 12192 17960 12220
rect 17405 12183 17463 12189
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 18800 12229 18828 12260
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12220 18199 12223
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18187 12192 18613 12220
rect 18187 12189 18199 12192
rect 18141 12183 18199 12189
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 16574 12152 16580 12164
rect 15948 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 17218 12152 17224 12164
rect 17179 12124 17224 12152
rect 17218 12112 17224 12124
rect 17276 12152 17282 12164
rect 18156 12152 18184 12183
rect 19702 12152 19708 12164
rect 17276 12124 18184 12152
rect 19260 12124 19708 12152
rect 17276 12112 17282 12124
rect 15378 12084 15384 12096
rect 12406 12056 15384 12084
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 17770 12044 17776 12096
rect 17828 12084 17834 12096
rect 19260 12084 19288 12124
rect 19702 12112 19708 12124
rect 19760 12112 19766 12164
rect 19794 12084 19800 12096
rect 17828 12056 19288 12084
rect 19755 12056 19800 12084
rect 17828 12044 17834 12056
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 1104 11994 21043 12016
rect 1104 11942 5894 11994
rect 5946 11942 5958 11994
rect 6010 11942 6022 11994
rect 6074 11942 6086 11994
rect 6138 11942 6150 11994
rect 6202 11942 10839 11994
rect 10891 11942 10903 11994
rect 10955 11942 10967 11994
rect 11019 11942 11031 11994
rect 11083 11942 11095 11994
rect 11147 11942 15784 11994
rect 15836 11942 15848 11994
rect 15900 11942 15912 11994
rect 15964 11942 15976 11994
rect 16028 11942 16040 11994
rect 16092 11942 20729 11994
rect 20781 11942 20793 11994
rect 20845 11942 20857 11994
rect 20909 11942 20921 11994
rect 20973 11942 20985 11994
rect 21037 11942 21043 11994
rect 1104 11920 21043 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 1854 11880 1860 11892
rect 1811 11852 1860 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 1854 11840 1860 11852
rect 1912 11840 1918 11892
rect 13725 11883 13783 11889
rect 13725 11849 13737 11883
rect 13771 11880 13783 11883
rect 14734 11880 14740 11892
rect 13771 11852 14740 11880
rect 13771 11849 13783 11852
rect 13725 11843 13783 11849
rect 14734 11840 14740 11852
rect 14792 11880 14798 11892
rect 15562 11880 15568 11892
rect 14792 11852 15568 11880
rect 14792 11840 14798 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18785 11883 18843 11889
rect 18785 11880 18797 11883
rect 18656 11852 18797 11880
rect 18656 11840 18662 11852
rect 18785 11849 18797 11852
rect 18831 11849 18843 11883
rect 18785 11843 18843 11849
rect 19610 11840 19616 11892
rect 19668 11840 19674 11892
rect 19794 11880 19800 11892
rect 19755 11852 19800 11880
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 3513 11815 3571 11821
rect 3513 11812 3525 11815
rect 1688 11784 3525 11812
rect 1688 11756 1716 11784
rect 3513 11781 3525 11784
rect 3559 11781 3571 11815
rect 19429 11815 19487 11821
rect 19429 11812 19441 11815
rect 3513 11775 3571 11781
rect 18616 11784 19441 11812
rect 18616 11756 18644 11784
rect 19429 11781 19441 11784
rect 19475 11781 19487 11815
rect 19429 11775 19487 11781
rect 19521 11815 19579 11821
rect 19521 11781 19533 11815
rect 19567 11812 19579 11815
rect 19628 11812 19656 11840
rect 19567 11784 19656 11812
rect 19567 11781 19579 11784
rect 19521 11775 19579 11781
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2406 11744 2412 11756
rect 1995 11716 2412 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5534 11744 5540 11756
rect 5215 11716 5540 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 6546 11744 6552 11756
rect 6507 11716 6552 11744
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6822 11753 6828 11756
rect 6816 11707 6828 11753
rect 6880 11744 6886 11756
rect 6880 11716 6916 11744
rect 6822 11704 6828 11707
rect 6880 11704 6886 11716
rect 11698 11704 11704 11756
rect 11756 11744 11762 11756
rect 12250 11744 12256 11756
rect 11756 11716 12256 11744
rect 11756 11704 11762 11716
rect 12250 11704 12256 11716
rect 12308 11744 12314 11756
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 12308 11716 12357 11744
rect 12308 11704 12314 11716
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12612 11747 12670 11753
rect 12612 11713 12624 11747
rect 12658 11744 12670 11747
rect 14918 11744 14924 11756
rect 12658 11716 14924 11744
rect 12658 11713 12670 11716
rect 12612 11707 12670 11713
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 15160 11716 18429 11744
rect 15160 11704 15166 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 18417 11707 18475 11713
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 4893 11679 4951 11685
rect 4893 11676 4905 11679
rect 2280 11648 4905 11676
rect 2280 11636 2286 11648
rect 4893 11645 4905 11648
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11645 15071 11679
rect 15013 11639 15071 11645
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11645 17463 11679
rect 18432 11676 18460 11707
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 18782 11704 18788 11756
rect 18840 11744 18846 11756
rect 19245 11747 19303 11753
rect 19245 11744 19257 11747
rect 18840 11716 19257 11744
rect 18840 11704 18846 11716
rect 19245 11713 19257 11716
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 19659 11716 19748 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 19426 11676 19432 11688
rect 18432 11648 19432 11676
rect 17405 11639 17463 11645
rect 1946 11608 1952 11620
rect 1907 11580 1952 11608
rect 1946 11568 1952 11580
rect 2004 11568 2010 11620
rect 15028 11608 15056 11639
rect 15102 11608 15108 11620
rect 15028 11580 15108 11608
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 15286 11608 15292 11620
rect 15247 11580 15292 11608
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 16724 11580 16865 11608
rect 16724 11568 16730 11580
rect 16853 11577 16865 11580
rect 16899 11577 16911 11611
rect 17310 11608 17316 11620
rect 17271 11580 17316 11608
rect 16853 11571 16911 11577
rect 17310 11568 17316 11580
rect 17368 11568 17374 11620
rect 17420 11608 17448 11639
rect 19426 11636 19432 11648
rect 19484 11676 19490 11688
rect 19720 11676 19748 11716
rect 19484 11648 19748 11676
rect 19484 11636 19490 11648
rect 19794 11608 19800 11620
rect 17420 11580 19800 11608
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7892 11512 7941 11540
rect 7892 11500 7898 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 7929 11503 7987 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 15712 11512 17233 11540
rect 15712 11500 15718 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17678 11540 17684 11552
rect 17639 11512 17684 11540
rect 17221 11503 17279 11509
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 1104 11450 20884 11472
rect 1104 11398 3422 11450
rect 3474 11398 3486 11450
rect 3538 11398 3550 11450
rect 3602 11398 3614 11450
rect 3666 11398 3678 11450
rect 3730 11398 8367 11450
rect 8419 11398 8431 11450
rect 8483 11398 8495 11450
rect 8547 11398 8559 11450
rect 8611 11398 8623 11450
rect 8675 11398 13312 11450
rect 13364 11398 13376 11450
rect 13428 11398 13440 11450
rect 13492 11398 13504 11450
rect 13556 11398 13568 11450
rect 13620 11398 18257 11450
rect 18309 11398 18321 11450
rect 18373 11398 18385 11450
rect 18437 11398 18449 11450
rect 18501 11398 18513 11450
rect 18565 11398 20884 11450
rect 1104 11376 20884 11398
rect 2222 11336 2228 11348
rect 2183 11308 2228 11336
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 16666 11336 16672 11348
rect 16627 11308 16672 11336
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18506 11336 18512 11348
rect 16960 11308 18512 11336
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 6825 11271 6883 11277
rect 6825 11268 6837 11271
rect 6696 11240 6837 11268
rect 6696 11228 6702 11240
rect 6825 11237 6837 11240
rect 6871 11237 6883 11271
rect 6825 11231 6883 11237
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 16960 11268 16988 11308
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 19610 11296 19616 11348
rect 19668 11336 19674 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19668 11308 19717 11336
rect 19668 11296 19674 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 15528 11240 16988 11268
rect 15528 11228 15534 11240
rect 17034 11228 17040 11280
rect 17092 11268 17098 11280
rect 17092 11240 19012 11268
rect 17092 11228 17098 11240
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12526 11200 12532 11212
rect 11664 11172 12532 11200
rect 11664 11160 11670 11172
rect 12526 11160 12532 11172
rect 12584 11200 12590 11212
rect 17310 11200 17316 11212
rect 12584 11172 15332 11200
rect 17271 11172 17316 11200
rect 12584 11160 12590 11172
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 1946 11132 1952 11144
rect 1728 11104 1952 11132
rect 1728 11092 1734 11104
rect 1946 11092 1952 11104
rect 2004 11132 2010 11144
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 2004 11104 2053 11132
rect 2004 11092 2010 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2406 11132 2412 11144
rect 2271 11104 2412 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5534 11132 5540 11144
rect 5491 11104 5540 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5712 11067 5770 11073
rect 5712 11033 5724 11067
rect 5758 11064 5770 11067
rect 5810 11064 5816 11076
rect 5758 11036 5816 11064
rect 5758 11033 5770 11036
rect 5712 11027 5770 11033
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 15013 11067 15071 11073
rect 15013 11033 15025 11067
rect 15059 11064 15071 11067
rect 15102 11064 15108 11076
rect 15059 11036 15108 11064
rect 15059 11033 15071 11036
rect 15013 11027 15071 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 15304 11064 15332 11172
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 17828 11172 18613 11200
rect 17828 11160 17834 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 16206 11132 16212 11144
rect 15427 11104 16212 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16724 11104 17141 11132
rect 16724 11092 16730 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 18138 11092 18144 11144
rect 18196 11132 18202 11144
rect 18782 11132 18788 11144
rect 18196 11104 18788 11132
rect 18196 11092 18202 11104
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11101 18935 11135
rect 18984 11132 19012 11240
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 18984 11104 19625 11132
rect 18877 11095 18935 11101
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 15304 11036 17080 11064
rect 17052 11005 17080 11036
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 18892 11064 18920 11095
rect 18564 11036 18920 11064
rect 18564 11024 18570 11036
rect 17037 10999 17095 11005
rect 17037 10965 17049 10999
rect 17083 10965 17095 10999
rect 18598 10996 18604 11008
rect 18559 10968 18604 10996
rect 17037 10959 17095 10965
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 1104 10906 21043 10928
rect 1104 10854 5894 10906
rect 5946 10854 5958 10906
rect 6010 10854 6022 10906
rect 6074 10854 6086 10906
rect 6138 10854 6150 10906
rect 6202 10854 10839 10906
rect 10891 10854 10903 10906
rect 10955 10854 10967 10906
rect 11019 10854 11031 10906
rect 11083 10854 11095 10906
rect 11147 10854 15784 10906
rect 15836 10854 15848 10906
rect 15900 10854 15912 10906
rect 15964 10854 15976 10906
rect 16028 10854 16040 10906
rect 16092 10854 20729 10906
rect 20781 10854 20793 10906
rect 20845 10854 20857 10906
rect 20909 10854 20921 10906
rect 20973 10854 20985 10906
rect 21037 10854 21043 10906
rect 1104 10832 21043 10854
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 16945 10795 17003 10801
rect 16945 10792 16957 10795
rect 14976 10764 16957 10792
rect 14976 10752 14982 10764
rect 16945 10761 16957 10764
rect 16991 10761 17003 10795
rect 18506 10792 18512 10804
rect 18467 10764 18512 10792
rect 16945 10755 17003 10761
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 1946 10684 1952 10736
rect 2004 10724 2010 10736
rect 17126 10733 17132 10736
rect 12520 10727 12578 10733
rect 2004 10696 2360 10724
rect 2004 10684 2010 10696
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2332 10665 2360 10696
rect 12520 10693 12532 10727
rect 12566 10724 12578 10727
rect 17113 10727 17132 10733
rect 12566 10696 17080 10724
rect 12566 10693 12578 10696
rect 12520 10687 12578 10693
rect 2225 10659 2283 10665
rect 2225 10656 2237 10659
rect 1912 10628 2237 10656
rect 1912 10616 1918 10628
rect 2225 10625 2237 10628
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 4718 10659 4776 10665
rect 4718 10656 4730 10659
rect 2924 10628 4730 10656
rect 2924 10616 2930 10628
rect 4718 10625 4730 10628
rect 4764 10625 4776 10659
rect 4718 10619 4776 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5534 10656 5540 10668
rect 5031 10628 5540 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 6604 10628 8033 10656
rect 6604 10616 6610 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 12250 10656 12256 10668
rect 12211 10628 12256 10656
rect 8021 10619 8079 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 14700 10628 15761 10656
rect 14700 10616 14706 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 2041 10591 2099 10597
rect 2041 10588 2053 10591
rect 1964 10560 2053 10588
rect 1964 10452 1992 10560
rect 2041 10557 2053 10560
rect 2087 10557 2099 10591
rect 2041 10551 2099 10557
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 8297 10591 8355 10597
rect 2179 10560 2728 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2700 10532 2728 10560
rect 8297 10557 8309 10591
rect 8343 10588 8355 10591
rect 9950 10588 9956 10600
rect 8343 10560 9956 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15160 10560 15485 10588
rect 15160 10548 15166 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 17052 10588 17080 10696
rect 17113 10693 17125 10727
rect 17113 10687 17132 10693
rect 17126 10684 17132 10687
rect 17184 10684 17190 10736
rect 17313 10727 17371 10733
rect 17313 10693 17325 10727
rect 17359 10724 17371 10727
rect 17770 10724 17776 10736
rect 17359 10696 17776 10724
rect 17359 10693 17371 10696
rect 17313 10687 17371 10693
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 18598 10684 18604 10736
rect 18656 10724 18662 10736
rect 18693 10727 18751 10733
rect 18693 10724 18705 10727
rect 18656 10696 18705 10724
rect 18656 10684 18662 10696
rect 18693 10693 18705 10696
rect 18739 10693 18751 10727
rect 19886 10724 19892 10736
rect 18693 10687 18751 10693
rect 19536 10696 19892 10724
rect 18138 10616 18144 10668
rect 18196 10656 18202 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18196 10628 18429 10656
rect 18196 10616 18202 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 19426 10656 19432 10668
rect 19387 10628 19432 10656
rect 18417 10619 18475 10625
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19536 10665 19564 10696
rect 19886 10684 19892 10696
rect 19944 10684 19950 10736
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 18598 10588 18604 10600
rect 17052 10560 18604 10588
rect 15473 10551 15531 10557
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19628 10588 19656 10619
rect 19208 10560 19656 10588
rect 19208 10548 19214 10560
rect 2682 10480 2688 10532
rect 2740 10520 2746 10532
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 2740 10492 3617 10520
rect 2740 10480 2746 10492
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 3605 10483 3663 10489
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 18693 10523 18751 10529
rect 18693 10520 18705 10523
rect 13780 10492 18705 10520
rect 13780 10480 13786 10492
rect 18693 10489 18705 10492
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 2406 10452 2412 10464
rect 1964 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2774 10452 2780 10464
rect 2547 10424 2780 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2774 10412 2780 10424
rect 2832 10412 2838 10464
rect 9585 10455 9643 10461
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 11606 10452 11612 10464
rect 9631 10424 11612 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 14550 10452 14556 10464
rect 13679 10424 14556 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 14918 10412 14924 10464
rect 14976 10452 14982 10464
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 14976 10424 15209 10452
rect 14976 10412 14982 10424
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 15197 10415 15255 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 17129 10455 17187 10461
rect 17129 10421 17141 10455
rect 17175 10452 17187 10455
rect 17954 10452 17960 10464
rect 17175 10424 17960 10452
rect 17175 10421 17187 10424
rect 17129 10415 17187 10421
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 19242 10452 19248 10464
rect 19203 10424 19248 10452
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 1104 10362 20884 10384
rect 1104 10310 3422 10362
rect 3474 10310 3486 10362
rect 3538 10310 3550 10362
rect 3602 10310 3614 10362
rect 3666 10310 3678 10362
rect 3730 10310 8367 10362
rect 8419 10310 8431 10362
rect 8483 10310 8495 10362
rect 8547 10310 8559 10362
rect 8611 10310 8623 10362
rect 8675 10310 13312 10362
rect 13364 10310 13376 10362
rect 13428 10310 13440 10362
rect 13492 10310 13504 10362
rect 13556 10310 13568 10362
rect 13620 10310 18257 10362
rect 18309 10310 18321 10362
rect 18373 10310 18385 10362
rect 18437 10310 18449 10362
rect 18501 10310 18513 10362
rect 18565 10310 20884 10362
rect 1104 10288 20884 10310
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2866 10248 2872 10260
rect 2823 10220 2872 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 15286 10257 15292 10260
rect 15243 10251 15292 10257
rect 15243 10217 15255 10251
rect 15289 10217 15292 10251
rect 15243 10211 15292 10217
rect 15286 10208 15292 10211
rect 15344 10208 15350 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 16209 10251 16267 10257
rect 16209 10248 16221 10251
rect 15620 10220 16221 10248
rect 15620 10208 15626 10220
rect 16209 10217 16221 10220
rect 16255 10217 16267 10251
rect 16209 10211 16267 10217
rect 17589 10251 17647 10257
rect 17589 10217 17601 10251
rect 17635 10248 17647 10251
rect 18138 10248 18144 10260
rect 17635 10220 18144 10248
rect 17635 10217 17647 10220
rect 17589 10211 17647 10217
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 2133 10183 2191 10189
rect 2133 10149 2145 10183
rect 2179 10149 2191 10183
rect 2133 10143 2191 10149
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 1946 10044 1952 10056
rect 1903 10016 1952 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2148 10044 2176 10143
rect 15102 10140 15108 10192
rect 15160 10180 15166 10192
rect 15160 10152 15424 10180
rect 15160 10140 15166 10152
rect 12161 10115 12219 10121
rect 12161 10081 12173 10115
rect 12207 10112 12219 10115
rect 12250 10112 12256 10124
rect 12207 10084 12256 10112
rect 12207 10081 12219 10084
rect 12161 10075 12219 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 2148 10016 2605 10044
rect 2593 10013 2605 10016
rect 2639 10013 2651 10047
rect 2593 10007 2651 10013
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 7742 10044 7748 10056
rect 2832 10016 2877 10044
rect 7703 10016 7748 10044
rect 2832 10004 2838 10016
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 14918 10044 14924 10056
rect 14879 10016 14924 10044
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15102 10044 15108 10056
rect 15063 10016 15108 10044
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15396 10053 15424 10152
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 17037 10183 17095 10189
rect 17037 10180 17049 10183
rect 16908 10152 17049 10180
rect 16908 10140 16914 10152
rect 17037 10149 17049 10152
rect 17083 10149 17095 10183
rect 17037 10143 17095 10149
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16868 10044 16896 10140
rect 18138 10112 18144 10124
rect 17328 10084 18144 10112
rect 17328 10053 17356 10084
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19484 10084 20116 10112
rect 19484 10072 19490 10084
rect 16623 10016 16896 10044
rect 17313 10047 17371 10053
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 2133 9979 2191 9985
rect 2133 9945 2145 9979
rect 2179 9976 2191 9979
rect 2682 9976 2688 9988
rect 2179 9948 2688 9976
rect 2179 9945 2191 9948
rect 2133 9939 2191 9945
rect 2682 9936 2688 9948
rect 2740 9936 2746 9988
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 9582 9976 9588 9988
rect 7055 9948 9588 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 9582 9936 9588 9948
rect 9640 9976 9646 9988
rect 10413 9979 10471 9985
rect 10413 9976 10425 9979
rect 9640 9948 10425 9976
rect 9640 9936 9646 9948
rect 10413 9945 10425 9948
rect 10459 9945 10471 9979
rect 10413 9939 10471 9945
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 15396 9976 15424 10007
rect 13964 9948 15424 9976
rect 16316 9976 16344 10007
rect 18046 10004 18052 10056
rect 18104 10044 18110 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18104 10016 18613 10044
rect 18104 10004 18110 10016
rect 18601 10013 18613 10016
rect 18647 10013 18659 10047
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 18601 10007 18659 10013
rect 19168 10016 19625 10044
rect 16316 9948 18828 9976
rect 13964 9936 13970 9948
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 1949 9911 2007 9917
rect 1949 9908 1961 9911
rect 1912 9880 1961 9908
rect 1912 9868 1918 9880
rect 1949 9877 1961 9880
rect 1995 9908 2007 9911
rect 2222 9908 2228 9920
rect 1995 9880 2228 9908
rect 1995 9877 2007 9880
rect 1949 9871 2007 9877
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 7837 9911 7895 9917
rect 7837 9877 7849 9911
rect 7883 9908 7895 9911
rect 7926 9908 7932 9920
rect 7883 9880 7932 9908
rect 7883 9877 7895 9880
rect 7837 9871 7895 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 15010 9908 15016 9920
rect 14971 9880 15016 9908
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15252 9880 16037 9908
rect 15252 9868 15258 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 17218 9908 17224 9920
rect 17179 9880 17224 9908
rect 16025 9871 16083 9877
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 17402 9868 17408 9920
rect 17460 9908 17466 9920
rect 18800 9917 18828 9948
rect 19168 9920 19196 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 19702 10004 19708 10056
rect 19760 10044 19766 10056
rect 19886 10044 19892 10056
rect 19760 10016 19892 10044
rect 19760 10004 19766 10016
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 20088 10053 20116 10084
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 18785 9911 18843 9917
rect 17460 9880 17505 9908
rect 17460 9868 17466 9880
rect 18785 9877 18797 9911
rect 18831 9908 18843 9911
rect 19150 9908 19156 9920
rect 18831 9880 19156 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 19426 9908 19432 9920
rect 19387 9880 19432 9908
rect 19426 9868 19432 9880
rect 19484 9868 19490 9920
rect 1104 9818 21043 9840
rect 1104 9766 5894 9818
rect 5946 9766 5958 9818
rect 6010 9766 6022 9818
rect 6074 9766 6086 9818
rect 6138 9766 6150 9818
rect 6202 9766 10839 9818
rect 10891 9766 10903 9818
rect 10955 9766 10967 9818
rect 11019 9766 11031 9818
rect 11083 9766 11095 9818
rect 11147 9766 15784 9818
rect 15836 9766 15848 9818
rect 15900 9766 15912 9818
rect 15964 9766 15976 9818
rect 16028 9766 16040 9818
rect 16092 9766 20729 9818
rect 20781 9766 20793 9818
rect 20845 9766 20857 9818
rect 20909 9766 20921 9818
rect 20973 9766 20985 9818
rect 21037 9766 21043 9818
rect 1104 9744 21043 9766
rect 14918 9664 14924 9716
rect 14976 9704 14982 9716
rect 15378 9704 15384 9716
rect 14976 9676 15384 9704
rect 14976 9664 14982 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17313 9707 17371 9713
rect 17313 9704 17325 9707
rect 17276 9676 17325 9704
rect 17276 9664 17282 9676
rect 17313 9673 17325 9676
rect 17359 9673 17371 9707
rect 17313 9667 17371 9673
rect 12520 9639 12578 9645
rect 9784 9608 12296 9636
rect 9784 9580 9812 9608
rect 12268 9580 12296 9608
rect 12520 9605 12532 9639
rect 12566 9636 12578 9639
rect 13722 9636 13728 9648
rect 12566 9608 13728 9636
rect 12566 9605 12578 9608
rect 12520 9599 12578 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 17954 9636 17960 9648
rect 17915 9608 17960 9636
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 19521 9639 19579 9645
rect 19521 9636 19533 9639
rect 19484 9608 19533 9636
rect 19484 9596 19490 9608
rect 19521 9605 19533 9608
rect 19567 9605 19579 9639
rect 19521 9599 19579 9605
rect 4614 9568 4620 9580
rect 4672 9577 4678 9580
rect 4584 9540 4620 9568
rect 4614 9528 4620 9540
rect 4672 9531 4684 9577
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5718 9568 5724 9580
rect 4939 9540 5724 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 4672 9528 4678 9531
rect 5718 9528 5724 9540
rect 5776 9568 5782 9580
rect 6546 9568 6552 9580
rect 5776 9540 6552 9568
rect 5776 9528 5782 9540
rect 6546 9528 6552 9540
rect 6604 9568 6610 9580
rect 8018 9577 8024 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 6604 9540 7757 9568
rect 6604 9528 6610 9540
rect 7745 9537 7757 9540
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 8012 9531 8024 9577
rect 8076 9568 8082 9580
rect 9766 9568 9772 9580
rect 8076 9540 8112 9568
rect 9679 9540 9772 9568
rect 8018 9528 8024 9531
rect 8076 9528 8082 9540
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10036 9571 10094 9577
rect 10036 9537 10048 9571
rect 10082 9568 10094 9571
rect 11974 9568 11980 9580
rect 10082 9540 11980 9568
rect 10082 9537 10094 9540
rect 10036 9531 10094 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12250 9568 12256 9580
rect 12211 9540 12256 9568
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 14090 9568 14096 9580
rect 12360 9540 14096 9568
rect 12360 9500 12388 9540
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14734 9528 14740 9580
rect 14792 9568 14798 9580
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14792 9540 14933 9568
rect 14792 9528 14798 9540
rect 14921 9537 14933 9540
rect 14967 9568 14979 9571
rect 17218 9568 17224 9580
rect 14967 9540 17224 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 17310 9528 17316 9580
rect 17368 9568 17374 9580
rect 17405 9571 17463 9577
rect 17405 9568 17417 9571
rect 17368 9540 17417 9568
rect 17368 9528 17374 9540
rect 17405 9537 17417 9540
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17552 9540 17877 9568
rect 17552 9528 17558 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18138 9568 18144 9580
rect 18095 9540 18144 9568
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18138 9528 18144 9540
rect 18196 9568 18202 9580
rect 18874 9568 18880 9580
rect 18196 9540 18880 9568
rect 18196 9528 18202 9540
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 19300 9540 19349 9568
rect 19300 9528 19306 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19610 9568 19616 9580
rect 19571 9540 19616 9568
rect 19337 9531 19395 9537
rect 19610 9528 19616 9540
rect 19668 9528 19674 9580
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 19886 9568 19892 9580
rect 19751 9540 19892 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 15194 9500 15200 9512
rect 11072 9472 12388 9500
rect 15155 9472 15200 9500
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 2832 9336 3525 9364
rect 2832 9324 2838 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 9125 9367 9183 9373
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 11072 9364 11100 9472
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15286 9460 15292 9512
rect 15344 9460 15350 9512
rect 13633 9435 13691 9441
rect 13633 9401 13645 9435
rect 13679 9432 13691 9435
rect 15304 9432 15332 9460
rect 13679 9404 15332 9432
rect 13679 9401 13691 9404
rect 13633 9395 13691 9401
rect 19794 9392 19800 9444
rect 19852 9432 19858 9444
rect 19889 9435 19947 9441
rect 19889 9432 19901 9435
rect 19852 9404 19901 9432
rect 19852 9392 19858 9404
rect 19889 9401 19901 9404
rect 19935 9401 19947 9435
rect 19889 9395 19947 9401
rect 9171 9336 11100 9364
rect 11149 9367 11207 9373
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11882 9364 11888 9376
rect 11195 9336 11888 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 13044 9336 15025 9364
rect 13044 9324 13050 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15013 9327 15071 9333
rect 15105 9367 15163 9373
rect 15105 9333 15117 9367
rect 15151 9364 15163 9367
rect 15286 9364 15292 9376
rect 15151 9336 15292 9364
rect 15151 9333 15163 9336
rect 15105 9327 15163 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 1104 9274 20884 9296
rect 1104 9222 3422 9274
rect 3474 9222 3486 9274
rect 3538 9222 3550 9274
rect 3602 9222 3614 9274
rect 3666 9222 3678 9274
rect 3730 9222 8367 9274
rect 8419 9222 8431 9274
rect 8483 9222 8495 9274
rect 8547 9222 8559 9274
rect 8611 9222 8623 9274
rect 8675 9222 13312 9274
rect 13364 9222 13376 9274
rect 13428 9222 13440 9274
rect 13492 9222 13504 9274
rect 13556 9222 13568 9274
rect 13620 9222 18257 9274
rect 18309 9222 18321 9274
rect 18373 9222 18385 9274
rect 18437 9222 18449 9274
rect 18501 9222 18513 9274
rect 18565 9222 20884 9274
rect 1104 9200 20884 9222
rect 4246 9160 4252 9172
rect 4207 9132 4252 9160
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 7742 9160 7748 9172
rect 6595 9132 7748 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13814 9160 13820 9172
rect 13587 9132 13820 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 14458 9120 14464 9172
rect 14516 9160 14522 9172
rect 14918 9160 14924 9172
rect 14516 9132 14924 9160
rect 14516 9120 14522 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15010 9120 15016 9172
rect 15068 9169 15074 9172
rect 15068 9163 15117 9169
rect 15068 9129 15071 9163
rect 15105 9129 15117 9163
rect 17218 9160 17224 9172
rect 17179 9132 17224 9160
rect 15068 9123 15117 9129
rect 15068 9120 15074 9123
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17402 9160 17408 9172
rect 17363 9132 17408 9160
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 19886 9160 19892 9172
rect 19847 9132 19892 9160
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 2682 9092 2688 9104
rect 2608 9064 2688 9092
rect 2608 9033 2636 9064
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9061 8539 9095
rect 8481 9055 8539 9061
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 8993 2651 9027
rect 2593 8987 2651 8993
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3142 8956 3148 8968
rect 2731 8928 3148 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 4120 8928 4169 8956
rect 4120 8916 4126 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 4430 8956 4436 8968
rect 4387 8928 4436 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5718 8956 5724 8968
rect 5215 8928 5724 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5718 8916 5724 8928
rect 5776 8956 5782 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 5776 8928 7113 8956
rect 5776 8916 5782 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 8496 8956 8524 9055
rect 14734 9052 14740 9104
rect 14792 9092 14798 9104
rect 15197 9095 15255 9101
rect 15197 9092 15209 9095
rect 14792 9064 15209 9092
rect 14792 9052 14798 9064
rect 15197 9061 15209 9064
rect 15243 9061 15255 9095
rect 15197 9055 15255 9061
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17310 9092 17316 9104
rect 17092 9064 17316 9092
rect 17092 9052 17098 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 15286 9024 15292 9036
rect 15247 8996 15292 9024
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 19150 9024 19156 9036
rect 16960 8996 19156 9024
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8496 8928 9137 8956
rect 7101 8919 7159 8925
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8956 12219 8959
rect 12250 8956 12256 8968
rect 12207 8928 12256 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12360 8928 14780 8956
rect 5414 8891 5472 8897
rect 5414 8888 5426 8891
rect 4356 8860 5426 8888
rect 4356 8832 4384 8860
rect 5414 8857 5426 8860
rect 5460 8857 5472 8891
rect 5414 8851 5472 8857
rect 7368 8891 7426 8897
rect 7368 8857 7380 8891
rect 7414 8888 7426 8891
rect 8110 8888 8116 8900
rect 7414 8860 8116 8888
rect 7414 8857 7426 8860
rect 7368 8851 7426 8857
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 10036 8891 10094 8897
rect 10036 8857 10048 8891
rect 10082 8888 10094 8891
rect 10686 8888 10692 8900
rect 10082 8860 10692 8888
rect 10082 8857 10094 8860
rect 10036 8851 10094 8857
rect 10686 8848 10692 8860
rect 10744 8848 10750 8900
rect 11606 8848 11612 8900
rect 11664 8888 11670 8900
rect 12360 8888 12388 8928
rect 11664 8860 12388 8888
rect 12428 8891 12486 8897
rect 11664 8848 11670 8860
rect 12428 8857 12440 8891
rect 12474 8888 12486 8891
rect 12802 8888 12808 8900
rect 12474 8860 12808 8888
rect 12474 8857 12486 8860
rect 12428 8851 12486 8857
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 14752 8888 14780 8928
rect 14826 8916 14832 8968
rect 14884 8956 14890 8968
rect 14921 8959 14979 8965
rect 14921 8956 14933 8959
rect 14884 8928 14933 8956
rect 14884 8916 14890 8928
rect 14921 8925 14933 8928
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 16960 8888 16988 8996
rect 19150 8984 19156 8996
rect 19208 9024 19214 9036
rect 19208 8996 19656 9024
rect 19208 8984 19214 8996
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19628 8965 19656 8996
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19300 8928 19533 8956
rect 19300 8916 19306 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 14752 8860 16988 8888
rect 17034 8848 17040 8900
rect 17092 8888 17098 8900
rect 19720 8888 19748 8919
rect 17092 8860 19748 8888
rect 17092 8848 17098 8860
rect 1854 8820 1860 8832
rect 1815 8792 1860 8820
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 4338 8780 4344 8832
rect 4396 8780 4402 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 9180 8792 9229 8820
rect 9180 8780 9186 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8820 11207 8823
rect 14458 8820 14464 8832
rect 11195 8792 14464 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 15010 8820 15016 8832
rect 14608 8792 15016 8820
rect 14608 8780 14614 8792
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 15562 8820 15568 8832
rect 15523 8792 15568 8820
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 17237 8823 17295 8829
rect 17237 8820 17249 8823
rect 16816 8792 17249 8820
rect 16816 8780 16822 8792
rect 17237 8789 17249 8792
rect 17283 8789 17295 8823
rect 17237 8783 17295 8789
rect 1104 8730 21043 8752
rect 1104 8678 5894 8730
rect 5946 8678 5958 8730
rect 6010 8678 6022 8730
rect 6074 8678 6086 8730
rect 6138 8678 6150 8730
rect 6202 8678 10839 8730
rect 10891 8678 10903 8730
rect 10955 8678 10967 8730
rect 11019 8678 11031 8730
rect 11083 8678 11095 8730
rect 11147 8678 15784 8730
rect 15836 8678 15848 8730
rect 15900 8678 15912 8730
rect 15964 8678 15976 8730
rect 16028 8678 16040 8730
rect 16092 8678 20729 8730
rect 20781 8678 20793 8730
rect 20845 8678 20857 8730
rect 20909 8678 20921 8730
rect 20973 8678 20985 8730
rect 21037 8678 21043 8730
rect 1104 8656 21043 8678
rect 4614 8616 4620 8628
rect 4575 8588 4620 8616
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5810 8616 5816 8628
rect 5767 8588 5816 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6822 8616 6828 8628
rect 6779 8588 6828 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7616 8588 7941 8616
rect 7616 8576 7622 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10744 8588 10793 8616
rect 10744 8576 10750 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 12897 8619 12955 8625
rect 12897 8616 12909 8619
rect 10928 8588 12909 8616
rect 10928 8576 10934 8588
rect 12897 8585 12909 8588
rect 12943 8585 12955 8619
rect 14734 8616 14740 8628
rect 14695 8588 14740 8616
rect 12897 8579 12955 8585
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 17034 8616 17040 8628
rect 15068 8588 17040 8616
rect 15068 8576 15074 8588
rect 3148 8560 3200 8566
rect 8846 8548 8852 8560
rect 8807 8520 8852 8548
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 9858 8548 9864 8560
rect 9815 8520 9864 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 10318 8548 10324 8560
rect 10183 8520 10324 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 10318 8508 10324 8520
rect 10376 8548 10382 8560
rect 10376 8520 11284 8548
rect 10376 8508 10382 8520
rect 3148 8502 3200 8508
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5592 8452 5641 8480
rect 5592 8440 5598 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5776 8452 6561 8480
rect 5776 8440 5782 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6730 8480 6736 8492
rect 6691 8452 6736 8480
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7650 8480 7656 8492
rect 7515 8452 7656 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4062 8412 4068 8424
rect 4019 8384 4068 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4338 8412 4344 8424
rect 4299 8384 4344 8412
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4522 8412 4528 8424
rect 4479 8384 4528 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 4522 8372 4528 8384
rect 4580 8412 4586 8424
rect 5442 8412 5448 8424
rect 4580 8384 5448 8412
rect 4580 8372 4586 8384
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 7300 8412 7328 8443
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 8110 8480 8116 8492
rect 7791 8452 8116 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 6236 8384 7328 8412
rect 6236 8372 6242 8384
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8260 8384 8953 8412
rect 8260 8372 8266 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 9232 8412 9260 8443
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 10229 8483 10287 8489
rect 9364 8452 9409 8480
rect 9364 8440 9370 8452
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10410 8480 10416 8492
rect 10275 8452 10416 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10410 8440 10416 8452
rect 10468 8480 10474 8492
rect 10870 8480 10876 8492
rect 10468 8452 10876 8480
rect 10468 8440 10474 8452
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 11146 8480 11152 8492
rect 11107 8452 11152 8480
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11256 8480 11284 8520
rect 11698 8508 11704 8560
rect 11756 8548 11762 8560
rect 11853 8551 11911 8557
rect 11853 8548 11865 8551
rect 11756 8520 11865 8548
rect 11756 8508 11762 8520
rect 11853 8517 11865 8520
rect 11899 8517 11911 8551
rect 12066 8548 12072 8560
rect 12027 8520 12072 8548
rect 11853 8511 11911 8517
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 14001 8551 14059 8557
rect 14001 8548 14013 8551
rect 13372 8520 14013 8548
rect 12434 8480 12440 8492
rect 11256 8452 12440 8480
rect 12434 8440 12440 8452
rect 12492 8480 12498 8492
rect 13372 8489 13400 8520
rect 14001 8517 14013 8520
rect 14047 8548 14059 8551
rect 15102 8548 15108 8560
rect 14047 8520 15108 8548
rect 14047 8517 14059 8520
rect 14001 8511 14059 8517
rect 15102 8508 15108 8520
rect 15160 8548 15166 8560
rect 15289 8551 15347 8557
rect 15289 8548 15301 8551
rect 15160 8520 15301 8548
rect 15160 8508 15166 8520
rect 15289 8517 15301 8520
rect 15335 8517 15347 8551
rect 15289 8511 15347 8517
rect 15381 8551 15439 8557
rect 15381 8517 15393 8551
rect 15427 8548 15439 8551
rect 15470 8548 15476 8560
rect 15427 8520 15476 8548
rect 15427 8517 15439 8520
rect 15381 8511 15439 8517
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 12838 8483 12896 8489
rect 12838 8480 12850 8483
rect 12492 8452 12850 8480
rect 12492 8440 12498 8452
rect 12838 8449 12850 8452
rect 12884 8449 12896 8483
rect 12838 8443 12896 8449
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8449 13415 8483
rect 13357 8443 13415 8449
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 15010 8480 15016 8492
rect 14971 8452 15016 8480
rect 13909 8443 13967 8449
rect 9861 8415 9919 8421
rect 9232 8384 9628 8412
rect 8941 8375 8999 8381
rect 9600 8356 9628 8384
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 9907 8384 11069 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 11057 8381 11069 8384
rect 11103 8412 11115 8415
rect 11330 8412 11336 8424
rect 11103 8384 11336 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 13924 8412 13952 8443
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 16132 8489 16160 8588
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17184 8588 17509 8616
rect 17184 8576 17190 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 19521 8619 19579 8625
rect 19521 8585 19533 8619
rect 19567 8616 19579 8619
rect 19610 8616 19616 8628
rect 19567 8588 19616 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8548 17003 8551
rect 17402 8548 17408 8560
rect 16991 8520 17408 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16758 8480 16764 8492
rect 16347 8452 16764 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8480 16911 8483
rect 17126 8480 17132 8492
rect 16899 8452 17132 8480
rect 16899 8449 16911 8452
rect 16853 8443 16911 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8481 17279 8483
rect 17267 8480 17280 8481
rect 17954 8480 17960 8492
rect 17267 8452 17960 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 19150 8480 19156 8492
rect 19111 8452 19156 8480
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 11940 8384 13952 8412
rect 11940 8372 11946 8384
rect 9582 8304 9588 8356
rect 9640 8344 9646 8356
rect 11238 8344 11244 8356
rect 9640 8316 11244 8344
rect 9640 8304 9646 8316
rect 11238 8304 11244 8316
rect 11296 8344 11302 8356
rect 12066 8344 12072 8356
rect 11296 8316 12072 8344
rect 11296 8304 11302 8316
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 13265 8347 13323 8353
rect 13265 8313 13277 8347
rect 13311 8344 13323 8347
rect 13924 8344 13952 8384
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14700 8384 14933 8412
rect 14700 8372 14706 8384
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 16114 8344 16120 8356
rect 13311 8316 13860 8344
rect 13924 8316 16120 8344
rect 13311 8313 13323 8316
rect 13265 8307 13323 8313
rect 9030 8276 9036 8288
rect 8991 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10042 8276 10048 8288
rect 9999 8248 10048 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 11149 8279 11207 8285
rect 11149 8245 11161 8279
rect 11195 8276 11207 8279
rect 11701 8279 11759 8285
rect 11701 8276 11713 8279
rect 11195 8248 11713 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 11701 8245 11713 8248
rect 11747 8245 11759 8279
rect 11882 8276 11888 8288
rect 11843 8248 11888 8276
rect 11701 8239 11759 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12710 8276 12716 8288
rect 12671 8248 12716 8276
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 13832 8276 13860 8316
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8344 16267 8347
rect 17034 8344 17040 8356
rect 16255 8316 17040 8344
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 17034 8304 17040 8316
rect 17092 8344 17098 8356
rect 17328 8344 17356 8375
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 19242 8412 19248 8424
rect 18196 8384 19248 8412
rect 18196 8372 18202 8384
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 17092 8316 17356 8344
rect 17092 8304 17098 8316
rect 13906 8276 13912 8288
rect 13832 8248 13912 8276
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 16942 8236 16948 8288
rect 17000 8276 17006 8288
rect 19153 8279 19211 8285
rect 19153 8276 19165 8279
rect 17000 8248 19165 8276
rect 17000 8236 17006 8248
rect 19153 8245 19165 8248
rect 19199 8245 19211 8279
rect 19153 8239 19211 8245
rect 1104 8186 20884 8208
rect 1104 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 3550 8186
rect 3602 8134 3614 8186
rect 3666 8134 3678 8186
rect 3730 8134 8367 8186
rect 8419 8134 8431 8186
rect 8483 8134 8495 8186
rect 8547 8134 8559 8186
rect 8611 8134 8623 8186
rect 8675 8134 13312 8186
rect 13364 8134 13376 8186
rect 13428 8134 13440 8186
rect 13492 8134 13504 8186
rect 13556 8134 13568 8186
rect 13620 8134 18257 8186
rect 18309 8134 18321 8186
rect 18373 8134 18385 8186
rect 18437 8134 18449 8186
rect 18501 8134 18513 8186
rect 18565 8134 20884 8186
rect 1104 8112 20884 8134
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6512 8044 6653 8072
rect 6512 8032 6518 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 7653 8075 7711 8081
rect 7653 8041 7665 8075
rect 7699 8072 7711 8075
rect 8018 8072 8024 8084
rect 7699 8044 8024 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 9088 8044 9321 8072
rect 9088 8032 9094 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 11204 8044 11345 8072
rect 11204 8032 11210 8044
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 12710 8072 12716 8084
rect 12115 8044 12716 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 12897 8075 12955 8081
rect 12897 8041 12909 8075
rect 12943 8072 12955 8075
rect 14182 8072 14188 8084
rect 12943 8044 14188 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 4430 7964 4436 8016
rect 4488 8004 4494 8016
rect 4525 8007 4583 8013
rect 4525 8004 4537 8007
rect 4488 7976 4537 8004
rect 4488 7964 4494 7976
rect 4525 7973 4537 7976
rect 4571 7973 4583 8007
rect 4525 7967 4583 7973
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12161 8007 12219 8013
rect 12161 8004 12173 8007
rect 12032 7976 12173 8004
rect 12032 7964 12038 7976
rect 12161 7973 12173 7976
rect 12207 7973 12219 8007
rect 12161 7967 12219 7973
rect 2038 7936 2044 7948
rect 1999 7908 2044 7936
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 5736 7908 7573 7936
rect 5736 7880 5764 7908
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7708 7908 7757 7936
rect 7708 7896 7714 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 12253 7939 12311 7945
rect 7745 7899 7803 7905
rect 9324 7908 11100 7936
rect 9324 7880 9352 7908
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4522 7868 4528 7880
rect 4387 7840 4528 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5166 7868 5172 7880
rect 5031 7840 5172 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 4632 7800 4660 7831
rect 5166 7828 5172 7840
rect 5224 7868 5230 7880
rect 5718 7868 5724 7880
rect 5224 7840 5724 7868
rect 5224 7828 5230 7840
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5868 7840 6009 7868
rect 5868 7828 5874 7840
rect 5997 7837 6009 7840
rect 6043 7837 6055 7871
rect 6178 7868 6184 7880
rect 6139 7840 6184 7868
rect 5997 7831 6055 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 6871 7840 7849 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7837 7837 7849 7840
rect 7883 7868 7895 7871
rect 8110 7868 8116 7880
rect 7883 7840 8116 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 5350 7800 5356 7812
rect 4632 7772 5356 7800
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 6840 7800 6868 7831
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 9306 7868 9312 7880
rect 9267 7840 9312 7868
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9582 7868 9588 7880
rect 9543 7840 9588 7868
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 11072 7877 11100 7908
rect 12253 7905 12265 7939
rect 12299 7936 12311 7939
rect 12912 7936 12940 8035
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 17000 8044 17233 8072
rect 17000 8032 17006 8044
rect 17221 8041 17233 8044
rect 17267 8041 17279 8075
rect 17221 8035 17279 8041
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 18831 8044 19625 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 12299 7908 12940 7936
rect 12299 7905 12311 7908
rect 12253 7899 12311 7905
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 15562 7936 15568 7948
rect 14240 7908 15568 7936
rect 14240 7896 14246 7908
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17310 7936 17316 7948
rect 16632 7908 17316 7936
rect 16632 7896 16638 7908
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 17828 7908 19840 7936
rect 17828 7896 17834 7908
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11698 7868 11704 7880
rect 11103 7840 11704 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11698 7828 11704 7840
rect 11756 7868 11762 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11756 7840 11989 7868
rect 11756 7828 11762 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 12710 7868 12716 7880
rect 12671 7840 12716 7868
rect 11977 7831 12035 7837
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 13964 7840 14381 7868
rect 13964 7828 13970 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 14918 7868 14924 7880
rect 14875 7840 14924 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 14918 7828 14924 7840
rect 14976 7868 14982 7880
rect 15102 7868 15108 7880
rect 14976 7840 15108 7868
rect 14976 7828 14982 7840
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16684 7840 17049 7868
rect 5500 7772 6868 7800
rect 7009 7803 7067 7809
rect 5500 7760 5506 7772
rect 7009 7769 7021 7803
rect 7055 7769 7067 7803
rect 7009 7763 7067 7769
rect 11149 7803 11207 7809
rect 11149 7769 11161 7803
rect 11195 7800 11207 7803
rect 11238 7800 11244 7812
rect 11195 7772 11244 7800
rect 11195 7769 11207 7772
rect 11149 7763 11207 7769
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 2590 7732 2596 7744
rect 2455 7704 2596 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6730 7732 6736 7744
rect 6227 7704 6736 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6730 7692 6736 7704
rect 6788 7732 6794 7744
rect 7024 7732 7052 7763
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 11333 7803 11391 7809
rect 11333 7769 11345 7803
rect 11379 7800 11391 7803
rect 11882 7800 11888 7812
rect 11379 7772 11888 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 11882 7760 11888 7772
rect 11940 7800 11946 7812
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 11940 7772 14565 7800
rect 11940 7760 11946 7772
rect 14553 7769 14565 7772
rect 14599 7800 14611 7803
rect 15010 7800 15016 7812
rect 14599 7772 15016 7800
rect 14599 7769 14611 7772
rect 14553 7763 14611 7769
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 6788 7704 7052 7732
rect 9493 7735 9551 7741
rect 6788 7692 6794 7704
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9766 7732 9772 7744
rect 9539 7704 9772 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9766 7692 9772 7704
rect 9824 7732 9830 7744
rect 10226 7732 10232 7744
rect 9824 7704 10232 7732
rect 9824 7692 9830 7704
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 16684 7732 16712 7840
rect 17037 7837 17049 7840
rect 17083 7868 17095 7871
rect 17402 7868 17408 7880
rect 17083 7840 17408 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 17402 7828 17408 7840
rect 17460 7868 17466 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17460 7840 17969 7868
rect 17460 7828 17466 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18233 7831 18291 7837
rect 18248 7800 18276 7831
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 19242 7868 19248 7880
rect 18932 7840 19248 7868
rect 18932 7828 18938 7840
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19334 7800 19340 7812
rect 18248 7772 19340 7800
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 19812 7809 19840 7908
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7769 19855 7803
rect 19797 7763 19855 7769
rect 16850 7732 16856 7744
rect 12308 7704 16712 7732
rect 16811 7704 16856 7732
rect 12308 7692 12314 7704
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 19610 7741 19616 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 17000 7704 19441 7732
rect 17000 7692 17006 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 19597 7735 19616 7741
rect 19597 7701 19609 7735
rect 19597 7695 19616 7701
rect 19610 7692 19616 7695
rect 19668 7692 19674 7744
rect 1104 7642 21043 7664
rect 1104 7590 5894 7642
rect 5946 7590 5958 7642
rect 6010 7590 6022 7642
rect 6074 7590 6086 7642
rect 6138 7590 6150 7642
rect 6202 7590 10839 7642
rect 10891 7590 10903 7642
rect 10955 7590 10967 7642
rect 11019 7590 11031 7642
rect 11083 7590 11095 7642
rect 11147 7590 15784 7642
rect 15836 7590 15848 7642
rect 15900 7590 15912 7642
rect 15964 7590 15976 7642
rect 16028 7590 16040 7642
rect 16092 7590 20729 7642
rect 20781 7590 20793 7642
rect 20845 7590 20857 7642
rect 20909 7590 20921 7642
rect 20973 7590 20985 7642
rect 21037 7590 21043 7642
rect 1104 7568 21043 7590
rect 4062 7528 4068 7540
rect 4023 7500 4068 7528
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4522 7528 4528 7540
rect 4479 7500 4528 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5534 7528 5540 7540
rect 5215 7500 5540 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5184 7460 5212 7491
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 10410 7528 10416 7540
rect 10060 7500 10416 7528
rect 5350 7460 5356 7472
rect 4540 7432 5212 7460
rect 5276 7432 5356 7460
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2222 7392 2228 7404
rect 2004 7364 2228 7392
rect 2004 7352 2010 7364
rect 2222 7352 2228 7364
rect 2280 7392 2286 7404
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2280 7364 2421 7392
rect 2280 7352 2286 7364
rect 2409 7361 2421 7364
rect 2455 7361 2467 7395
rect 2590 7392 2596 7404
rect 2551 7364 2596 7392
rect 2409 7355 2467 7361
rect 2590 7352 2596 7364
rect 2648 7352 2654 7404
rect 4540 7401 4568 7432
rect 5276 7401 5304 7432
rect 5350 7420 5356 7432
rect 5408 7460 5414 7472
rect 7650 7460 7656 7472
rect 5408 7432 7656 7460
rect 5408 7420 5414 7432
rect 7650 7420 7656 7432
rect 7708 7420 7714 7472
rect 10060 7469 10088 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 16942 7528 16948 7540
rect 12406 7500 16948 7528
rect 10045 7463 10103 7469
rect 10045 7429 10057 7463
rect 10091 7429 10103 7463
rect 10045 7423 10103 7429
rect 10226 7420 10232 7472
rect 10284 7460 10290 7472
rect 12250 7460 12256 7472
rect 10284 7432 12256 7460
rect 10284 7420 10290 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4525 7355 4583 7361
rect 5000 7364 5089 7392
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7293 2375 7327
rect 2498 7324 2504 7336
rect 2459 7296 2504 7324
rect 2317 7287 2375 7293
rect 2332 7256 2360 7287
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 4264 7324 4292 7355
rect 4338 7324 4344 7336
rect 4251 7296 4344 7324
rect 4338 7284 4344 7296
rect 4396 7324 4402 7336
rect 4890 7324 4896 7336
rect 4396 7296 4896 7324
rect 4396 7284 4402 7296
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 3142 7256 3148 7268
rect 2332 7228 3148 7256
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 2130 7188 2136 7200
rect 2091 7160 2136 7188
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 5000 7188 5028 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7361 5319 7395
rect 5902 7392 5908 7404
rect 5815 7364 5908 7392
rect 5261 7355 5319 7361
rect 5902 7352 5908 7364
rect 5960 7392 5966 7404
rect 6270 7392 6276 7404
rect 5960 7364 6276 7392
rect 5960 7352 5966 7364
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10376 7364 10421 7392
rect 10376 7352 10382 7364
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7293 5871 7327
rect 5813 7287 5871 7293
rect 5074 7216 5080 7268
rect 5132 7256 5138 7268
rect 5828 7256 5856 7287
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 12406 7324 12434 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 19429 7531 19487 7537
rect 17184 7500 17264 7528
rect 17184 7488 17190 7500
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 13541 7463 13599 7469
rect 13541 7460 13553 7463
rect 12584 7432 13553 7460
rect 12584 7420 12590 7432
rect 13541 7429 13553 7432
rect 13587 7429 13599 7463
rect 13541 7423 13599 7429
rect 15562 7420 15568 7472
rect 15620 7460 15626 7472
rect 15620 7432 17172 7460
rect 15620 7420 15626 7432
rect 13814 7392 13820 7404
rect 13775 7364 13820 7392
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 14829 7355 14887 7361
rect 13722 7324 13728 7336
rect 9456 7296 12434 7324
rect 13683 7296 13728 7324
rect 9456 7284 9462 7296
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 14458 7324 14464 7336
rect 14419 7296 14464 7324
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7293 14703 7327
rect 14844 7324 14872 7355
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 15654 7352 15660 7404
rect 15712 7392 15718 7404
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 15712 7364 15761 7392
rect 15712 7352 15718 7364
rect 15749 7361 15761 7364
rect 15795 7361 15807 7395
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 15749 7355 15807 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17034 7392 17040 7404
rect 16995 7364 17040 7392
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 17144 7401 17172 7432
rect 17236 7401 17264 7500
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 19610 7528 19616 7540
rect 19475 7500 19616 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 17862 7460 17868 7472
rect 17368 7432 17868 7460
rect 17368 7420 17374 7432
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7392 17279 7395
rect 17678 7392 17684 7404
rect 17267 7364 17684 7392
rect 17267 7361 17279 7364
rect 17221 7355 17279 7361
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 18690 7392 18696 7404
rect 17972 7364 18696 7392
rect 14844 7296 15608 7324
rect 14645 7287 14703 7293
rect 10042 7256 10048 7268
rect 5132 7228 5856 7256
rect 10003 7228 10048 7256
rect 5132 7216 5138 7228
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 14001 7259 14059 7265
rect 12124 7228 13952 7256
rect 12124 7216 12130 7228
rect 5534 7188 5540 7200
rect 2372 7160 5540 7188
rect 2372 7148 2378 7160
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 13630 7188 13636 7200
rect 11664 7160 13636 7188
rect 11664 7148 11670 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13924 7188 13952 7228
rect 14001 7225 14013 7259
rect 14047 7256 14059 7259
rect 14660 7256 14688 7287
rect 15580 7265 15608 7296
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 17972 7333 18000 7364
rect 18690 7352 18696 7364
rect 18748 7392 18754 7404
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18748 7364 19073 7392
rect 18748 7352 18754 7364
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19242 7392 19248 7404
rect 19203 7364 19248 7392
rect 19061 7355 19119 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 16816 7296 17969 7324
rect 16816 7284 16822 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18196 7296 18429 7324
rect 18196 7284 18202 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 14047 7228 14688 7256
rect 15565 7259 15623 7265
rect 14047 7225 14059 7228
rect 14001 7219 14059 7225
rect 15565 7225 15577 7259
rect 15611 7225 15623 7259
rect 15565 7219 15623 7225
rect 16040 7228 17632 7256
rect 14274 7188 14280 7200
rect 13924 7160 14280 7188
rect 14274 7148 14280 7160
rect 14332 7188 14338 7200
rect 16040 7197 16068 7228
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 14332 7160 16037 7188
rect 14332 7148 14338 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 17494 7188 17500 7200
rect 17455 7160 17500 7188
rect 16025 7151 16083 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 17604 7188 17632 7228
rect 17862 7216 17868 7268
rect 17920 7256 17926 7268
rect 18049 7259 18107 7265
rect 18049 7256 18061 7259
rect 17920 7228 18061 7256
rect 17920 7216 17926 7228
rect 18049 7225 18061 7228
rect 18095 7225 18107 7259
rect 18049 7219 18107 7225
rect 19702 7188 19708 7200
rect 17604 7160 19708 7188
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 1104 7098 20884 7120
rect 1104 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 3550 7098
rect 3602 7046 3614 7098
rect 3666 7046 3678 7098
rect 3730 7046 8367 7098
rect 8419 7046 8431 7098
rect 8483 7046 8495 7098
rect 8547 7046 8559 7098
rect 8611 7046 8623 7098
rect 8675 7046 13312 7098
rect 13364 7046 13376 7098
rect 13428 7046 13440 7098
rect 13492 7046 13504 7098
rect 13556 7046 13568 7098
rect 13620 7046 18257 7098
rect 18309 7046 18321 7098
rect 18373 7046 18385 7098
rect 18437 7046 18449 7098
rect 18501 7046 18513 7098
rect 18565 7046 20884 7098
rect 1104 7024 20884 7046
rect 5166 6984 5172 6996
rect 5127 6956 5172 6984
rect 5166 6944 5172 6956
rect 5224 6944 5230 6996
rect 10321 6987 10379 6993
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 12894 6984 12900 6996
rect 10367 6956 12900 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 6454 6916 6460 6928
rect 5552 6888 6460 6916
rect 5552 6860 5580 6888
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 11698 6916 11704 6928
rect 11659 6888 11704 6916
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 12250 6916 12256 6928
rect 12211 6888 12256 6916
rect 12250 6876 12256 6888
rect 12308 6876 12314 6928
rect 13722 6916 13728 6928
rect 12912 6888 13728 6916
rect 5350 6848 5356 6860
rect 5311 6820 5356 6848
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5902 6848 5908 6860
rect 5675 6820 5908 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 12710 6848 12716 6860
rect 6288 6820 12716 6848
rect 1854 6780 1860 6792
rect 1815 6752 1860 6780
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 2130 6780 2136 6792
rect 2091 6752 2136 6780
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6288 6789 6316 6820
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 12912 6857 12940 6888
rect 13722 6876 13728 6888
rect 13780 6916 13786 6928
rect 16206 6916 16212 6928
rect 13780 6888 16212 6916
rect 13780 6876 13786 6888
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 7650 6780 7656 6792
rect 7611 6752 7656 6780
rect 6273 6743 6331 6749
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 6288 6712 6316 6743
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 2004 6684 6316 6712
rect 2004 6672 2010 6684
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 7760 6712 7788 6743
rect 7616 6684 7788 6712
rect 7852 6712 7880 6743
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 7984 6752 8029 6780
rect 7984 6740 7990 6752
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10468 6752 11192 6780
rect 10468 6740 10474 6752
rect 8018 6712 8024 6724
rect 7852 6684 8024 6712
rect 7616 6672 7622 6684
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 10505 6715 10563 6721
rect 10505 6712 10517 6715
rect 8996 6684 10517 6712
rect 8996 6672 9002 6684
rect 10505 6681 10517 6684
rect 10551 6681 10563 6715
rect 10505 6675 10563 6681
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3694 6644 3700 6656
rect 2915 6616 3700 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 7742 6644 7748 6656
rect 7515 6616 7748 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 10137 6647 10195 6653
rect 10137 6644 10149 6647
rect 10008 6616 10149 6644
rect 10008 6604 10014 6616
rect 10137 6613 10149 6616
rect 10183 6613 10195 6647
rect 10137 6607 10195 6613
rect 10305 6647 10363 6653
rect 10305 6613 10317 6647
rect 10351 6644 10363 6647
rect 10686 6644 10692 6656
rect 10351 6616 10692 6644
rect 10351 6613 10363 6616
rect 10305 6607 10363 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11164 6644 11192 6752
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11848 6752 11989 6780
rect 11848 6740 11854 6752
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12434 6780 12440 6792
rect 12115 6752 12440 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 12434 6740 12440 6752
rect 12492 6780 12498 6792
rect 13173 6783 13231 6789
rect 12492 6752 13124 6780
rect 12492 6740 12498 6752
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 12986 6712 12992 6724
rect 11296 6684 12992 6712
rect 11296 6672 11302 6684
rect 12986 6672 12992 6684
rect 13044 6672 13050 6724
rect 13096 6712 13124 6752
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13906 6780 13912 6792
rect 13219 6752 13912 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6780 14427 6783
rect 14553 6783 14611 6789
rect 14415 6752 14504 6780
rect 14415 6749 14427 6752
rect 14369 6743 14427 6749
rect 14476 6712 14504 6752
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14660 6780 14688 6888
rect 16206 6876 16212 6888
rect 16264 6876 16270 6928
rect 17405 6919 17463 6925
rect 17405 6885 17417 6919
rect 17451 6885 17463 6919
rect 17405 6879 17463 6885
rect 17420 6848 17448 6879
rect 17420 6820 18184 6848
rect 14599 6752 14688 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 16448 6752 17141 6780
rect 16448 6740 16454 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17310 6780 17316 6792
rect 17267 6752 17316 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6780 17463 6783
rect 17494 6780 17500 6792
rect 17451 6752 17500 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17644 6752 17877 6780
rect 17644 6740 17650 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 18046 6780 18052 6792
rect 18007 6752 18052 6780
rect 17865 6743 17923 6749
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 18156 6789 18184 6820
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6749 18199 6783
rect 18141 6743 18199 6749
rect 15010 6712 15016 6724
rect 13096 6684 14504 6712
rect 14971 6684 15016 6712
rect 11885 6647 11943 6653
rect 11885 6644 11897 6647
rect 11164 6616 11897 6644
rect 11885 6613 11897 6616
rect 11931 6644 11943 6647
rect 11974 6644 11980 6656
rect 11931 6616 11980 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12526 6644 12532 6656
rect 12124 6616 12532 6644
rect 12124 6604 12130 6616
rect 12526 6604 12532 6616
rect 12584 6644 12590 6656
rect 13722 6644 13728 6656
rect 12584 6616 13728 6644
rect 12584 6604 12590 6616
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14476 6644 14504 6684
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15654 6644 15660 6656
rect 14476 6616 15660 6644
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 18141 6647 18199 6653
rect 18141 6613 18153 6647
rect 18187 6644 18199 6647
rect 18598 6644 18604 6656
rect 18187 6616 18604 6644
rect 18187 6613 18199 6616
rect 18141 6607 18199 6613
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 1104 6554 21043 6576
rect 1104 6502 5894 6554
rect 5946 6502 5958 6554
rect 6010 6502 6022 6554
rect 6074 6502 6086 6554
rect 6138 6502 6150 6554
rect 6202 6502 10839 6554
rect 10891 6502 10903 6554
rect 10955 6502 10967 6554
rect 11019 6502 11031 6554
rect 11083 6502 11095 6554
rect 11147 6502 15784 6554
rect 15836 6502 15848 6554
rect 15900 6502 15912 6554
rect 15964 6502 15976 6554
rect 16028 6502 16040 6554
rect 16092 6502 20729 6554
rect 20781 6502 20793 6554
rect 20845 6502 20857 6554
rect 20909 6502 20921 6554
rect 20973 6502 20985 6554
rect 21037 6502 21043 6554
rect 1104 6480 21043 6502
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 8938 6440 8944 6452
rect 6512 6412 8944 6440
rect 6512 6400 6518 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9272 6412 9597 6440
rect 9272 6400 9278 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 11330 6440 11336 6452
rect 9585 6403 9643 6409
rect 9968 6412 11336 6440
rect 3053 6375 3111 6381
rect 3053 6341 3065 6375
rect 3099 6372 3111 6375
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3099 6344 3801 6372
rect 3099 6341 3111 6344
rect 3053 6335 3111 6341
rect 3789 6341 3801 6344
rect 3835 6372 3847 6375
rect 4801 6375 4859 6381
rect 4801 6372 4813 6375
rect 3835 6344 4813 6372
rect 3835 6341 3847 6344
rect 3789 6335 3847 6341
rect 4801 6341 4813 6344
rect 4847 6341 4859 6375
rect 4801 6335 4859 6341
rect 5166 6332 5172 6384
rect 5224 6372 5230 6384
rect 5224 6344 6224 6372
rect 5224 6332 5230 6344
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2041 6267 2099 6273
rect 2884 6276 2973 6304
rect 2056 6168 2084 6267
rect 2884 6236 2912 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 3142 6304 3148 6316
rect 3103 6276 3148 6304
rect 2961 6267 3019 6273
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3970 6304 3976 6316
rect 3252 6276 3976 6304
rect 3252 6236 3280 6276
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5031 6276 5641 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5810 6304 5816 6316
rect 5771 6276 5816 6304
rect 5629 6267 5687 6273
rect 3694 6236 3700 6248
rect 2884 6208 3280 6236
rect 3655 6208 3700 6236
rect 3694 6196 3700 6208
rect 3752 6236 3758 6248
rect 5000 6236 5028 6267
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6196 6304 6224 6344
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 7377 6375 7435 6381
rect 7377 6372 7389 6375
rect 6328 6344 7389 6372
rect 6328 6332 6334 6344
rect 7377 6341 7389 6344
rect 7423 6341 7435 6375
rect 7377 6335 7435 6341
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 8846 6372 8852 6384
rect 7708 6344 8852 6372
rect 7708 6332 7714 6344
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 6822 6304 6828 6316
rect 6196 6276 6684 6304
rect 6783 6276 6828 6304
rect 3752 6208 5028 6236
rect 5721 6239 5779 6245
rect 3752 6196 3758 6208
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 5767 6208 6561 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6656 6236 6684 6276
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7742 6304 7748 6316
rect 7703 6276 7748 6304
rect 7009 6267 7067 6273
rect 7024 6236 7052 6267
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8202 6304 8208 6316
rect 7975 6276 8208 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 6656 6208 7052 6236
rect 6549 6199 6607 6205
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7944 6236 7972 6267
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 8864 6304 8892 6332
rect 8956 6313 8984 6400
rect 9490 6332 9496 6384
rect 9548 6372 9554 6384
rect 9548 6344 9904 6372
rect 9548 6332 9554 6344
rect 8711 6276 8892 6304
rect 8941 6307 8999 6313
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 9122 6304 9128 6316
rect 9083 6276 9128 6304
rect 8941 6267 8999 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9766 6304 9772 6316
rect 9727 6276 9772 6304
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 9876 6313 9904 6344
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6273 9919 6307
rect 9968 6304 9996 6412
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 11974 6440 11980 6452
rect 11931 6412 11980 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 13170 6440 13176 6452
rect 12115 6412 13176 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 13780 6412 16436 6440
rect 13780 6400 13786 6412
rect 16298 6372 16304 6384
rect 10888 6344 16304 6372
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9968 6276 10057 6304
rect 9861 6267 9919 6273
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10226 6304 10232 6316
rect 10183 6276 10232 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 7156 6208 7972 6236
rect 7156 6196 7162 6208
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8076 6208 8861 6236
rect 8076 6196 8082 6208
rect 8849 6205 8861 6208
rect 8895 6236 8907 6239
rect 9950 6236 9956 6248
rect 8895 6208 9956 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 9950 6196 9956 6208
rect 10008 6236 10014 6248
rect 10152 6236 10180 6267
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10888 6313 10916 6344
rect 16298 6332 16304 6344
rect 16356 6332 16362 6384
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11238 6304 11244 6316
rect 11195 6276 11244 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11664 6276 11713 6304
rect 11664 6264 11670 6276
rect 11701 6273 11713 6276
rect 11747 6304 11759 6307
rect 11790 6304 11796 6316
rect 11747 6276 11796 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 16408 6304 16436 6412
rect 17494 6400 17500 6452
rect 17552 6440 17558 6452
rect 17881 6443 17939 6449
rect 17881 6440 17893 6443
rect 17552 6412 17893 6440
rect 17552 6400 17558 6412
rect 17881 6409 17893 6412
rect 17927 6409 17939 6443
rect 18046 6440 18052 6452
rect 18007 6412 18052 6440
rect 17881 6403 17939 6409
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 19334 6440 19340 6452
rect 19295 6412 19340 6440
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 17310 6332 17316 6384
rect 17368 6372 17374 6384
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 17368 6344 17693 6372
rect 17368 6332 17374 6344
rect 17681 6341 17693 6344
rect 17727 6341 17739 6375
rect 17681 6335 17739 6341
rect 16482 6304 16488 6316
rect 12032 6276 12077 6304
rect 12176 6276 15424 6304
rect 16395 6276 16488 6304
rect 12032 6264 12038 6276
rect 10008 6208 10180 6236
rect 10008 6196 10014 6208
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 10744 6208 11069 6236
rect 10744 6196 10750 6208
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 2406 6168 2412 6180
rect 2056 6140 2412 6168
rect 2406 6128 2412 6140
rect 2464 6168 2470 6180
rect 7116 6168 7144 6196
rect 2464 6140 7144 6168
rect 2464 6128 2470 6140
rect 7558 6128 7564 6180
rect 7616 6168 7622 6180
rect 8757 6171 8815 6177
rect 8757 6168 8769 6171
rect 7616 6140 8769 6168
rect 7616 6128 7622 6140
rect 8757 6137 8769 6140
rect 8803 6168 8815 6171
rect 10042 6168 10048 6180
rect 8803 6140 10048 6168
rect 8803 6137 8815 6140
rect 8757 6131 8815 6137
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 12176 6168 12204 6276
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12308 6208 12353 6236
rect 12308 6196 12314 6208
rect 13078 6196 13084 6248
rect 13136 6236 13142 6248
rect 13906 6236 13912 6248
rect 13136 6208 13912 6236
rect 13136 6196 13142 6208
rect 13906 6196 13912 6208
rect 13964 6236 13970 6248
rect 15286 6236 15292 6248
rect 13964 6208 15292 6236
rect 13964 6196 13970 6208
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 15396 6236 15424 6276
rect 16482 6264 16488 6276
rect 16540 6304 16546 6316
rect 17067 6307 17125 6313
rect 17067 6304 17079 6307
rect 16540 6276 17079 6304
rect 16540 6264 16546 6276
rect 17067 6273 17079 6276
rect 17113 6273 17125 6307
rect 17218 6304 17224 6316
rect 17179 6276 17224 6304
rect 17067 6267 17125 6273
rect 17218 6264 17224 6276
rect 17276 6304 17282 6316
rect 18138 6304 18144 6316
rect 17276 6276 18144 6304
rect 17276 6264 17282 6276
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18598 6264 18604 6316
rect 18656 6304 18662 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 18656 6276 19257 6304
rect 18656 6264 18662 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 19886 6236 19892 6248
rect 15396 6208 19892 6236
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 13633 6171 13691 6177
rect 10612 6140 12204 6168
rect 12268 6140 13584 6168
rect 4246 6100 4252 6112
rect 4207 6072 4252 6100
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 8260 6072 8493 6100
rect 8260 6060 8266 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 8481 6063 8539 6069
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 10612 6100 10640 6140
rect 9548 6072 10640 6100
rect 10689 6103 10747 6109
rect 9548 6060 9554 6072
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 10778 6100 10784 6112
rect 10735 6072 10784 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 12066 6100 12072 6112
rect 11388 6072 12072 6100
rect 11388 6060 11394 6072
rect 12066 6060 12072 6072
rect 12124 6100 12130 6112
rect 12268 6100 12296 6140
rect 12124 6072 12296 6100
rect 12124 6060 12130 6072
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 13044 6072 13461 6100
rect 13044 6060 13050 6072
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 13556 6100 13584 6140
rect 13633 6137 13645 6171
rect 13679 6168 13691 6171
rect 13814 6168 13820 6180
rect 13679 6140 13820 6168
rect 13679 6137 13691 6140
rect 13633 6131 13691 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 16298 6128 16304 6180
rect 16356 6168 16362 6180
rect 16666 6168 16672 6180
rect 16356 6140 16672 6168
rect 16356 6128 16362 6140
rect 16666 6128 16672 6140
rect 16724 6168 16730 6180
rect 16853 6171 16911 6177
rect 16853 6168 16865 6171
rect 16724 6140 16865 6168
rect 16724 6128 16730 6140
rect 16853 6137 16865 6140
rect 16899 6137 16911 6171
rect 16853 6131 16911 6137
rect 17586 6100 17592 6112
rect 13556 6072 17592 6100
rect 13449 6063 13507 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17862 6100 17868 6112
rect 17823 6072 17868 6100
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 1104 6010 20884 6032
rect 1104 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 3550 6010
rect 3602 5958 3614 6010
rect 3666 5958 3678 6010
rect 3730 5958 8367 6010
rect 8419 5958 8431 6010
rect 8483 5958 8495 6010
rect 8547 5958 8559 6010
rect 8611 5958 8623 6010
rect 8675 5958 13312 6010
rect 13364 5958 13376 6010
rect 13428 5958 13440 6010
rect 13492 5958 13504 6010
rect 13556 5958 13568 6010
rect 13620 5958 18257 6010
rect 18309 5958 18321 6010
rect 18373 5958 18385 6010
rect 18437 5958 18449 6010
rect 18501 5958 18513 6010
rect 18565 5958 20884 6010
rect 1104 5936 20884 5958
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3970 5896 3976 5908
rect 3007 5868 3976 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10652 5868 10701 5896
rect 10652 5856 10658 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 12894 5896 12900 5908
rect 12855 5868 12900 5896
rect 10689 5859 10747 5865
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13630 5896 13636 5908
rect 13311 5868 13636 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13630 5856 13636 5868
rect 13688 5896 13694 5908
rect 13688 5868 14964 5896
rect 13688 5856 13694 5868
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 5997 5831 6055 5837
rect 5997 5828 6009 5831
rect 5408 5800 6009 5828
rect 5408 5788 5414 5800
rect 5997 5797 6009 5800
rect 6043 5797 6055 5831
rect 5997 5791 6055 5797
rect 8110 5788 8116 5840
rect 8168 5828 8174 5840
rect 8297 5831 8355 5837
rect 8297 5828 8309 5831
rect 8168 5800 8309 5828
rect 8168 5788 8174 5800
rect 8297 5797 8309 5800
rect 8343 5797 8355 5831
rect 10778 5828 10784 5840
rect 10739 5800 10784 5828
rect 8297 5791 8355 5797
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 4304 5732 7880 5760
rect 4304 5720 4310 5732
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2222 5692 2228 5704
rect 2179 5664 2228 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2406 5692 2412 5704
rect 2363 5664 2412 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 2866 5692 2872 5704
rect 2547 5664 2872 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 2866 5652 2872 5664
rect 2924 5692 2930 5704
rect 3145 5695 3203 5701
rect 3145 5692 3157 5695
rect 2924 5664 3157 5692
rect 2924 5652 2930 5664
rect 3145 5661 3157 5664
rect 3191 5661 3203 5695
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 3145 5655 3203 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6270 5692 6276 5704
rect 6227 5664 6276 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7852 5701 7880 5732
rect 13078 5720 13084 5772
rect 13136 5760 13142 5772
rect 14936 5769 14964 5868
rect 15286 5828 15292 5840
rect 15028 5800 15292 5828
rect 15028 5769 15056 5800
rect 15286 5788 15292 5800
rect 15344 5828 15350 5840
rect 18598 5828 18604 5840
rect 15344 5800 18604 5828
rect 15344 5788 15350 5800
rect 18598 5788 18604 5800
rect 18656 5788 18662 5840
rect 14921 5763 14979 5769
rect 13136 5732 13216 5760
rect 13136 5720 13142 5732
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7432 5664 7573 5692
rect 7432 5652 7438 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 8352 5664 8401 5692
rect 8352 5652 8358 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9398 5692 9404 5704
rect 8904 5664 9404 5692
rect 8904 5652 8910 5664
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9950 5701 9956 5704
rect 9907 5695 9956 5701
rect 9907 5661 9919 5695
rect 9953 5661 9956 5695
rect 9907 5655 9956 5661
rect 9950 5652 9956 5655
rect 10008 5652 10014 5704
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 10100 5664 10149 5692
rect 10100 5652 10106 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 6549 5627 6607 5633
rect 6549 5593 6561 5627
rect 6595 5624 6607 5627
rect 7282 5624 7288 5636
rect 6595 5596 7288 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 10152 5624 10180 5655
rect 10410 5652 10416 5704
rect 10468 5692 10474 5704
rect 13188 5701 13216 5732
rect 14921 5729 14933 5763
rect 14967 5729 14979 5763
rect 14921 5723 14979 5729
rect 15013 5763 15071 5769
rect 15013 5729 15025 5763
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 15102 5720 15108 5772
rect 15160 5760 15166 5772
rect 15473 5763 15531 5769
rect 15160 5732 15332 5760
rect 15160 5720 15166 5732
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10468 5664 10701 5692
rect 10468 5652 10474 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 13173 5695 13231 5701
rect 10689 5655 10747 5661
rect 10796 5664 13124 5692
rect 10796 5624 10824 5664
rect 10152 5596 10824 5624
rect 10965 5627 11023 5633
rect 10965 5593 10977 5627
rect 11011 5624 11023 5627
rect 11330 5624 11336 5636
rect 11011 5596 11336 5624
rect 11011 5593 11023 5596
rect 10965 5587 11023 5593
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 13096 5624 13124 5664
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 14182 5692 14188 5704
rect 13320 5664 13365 5692
rect 13556 5664 14188 5692
rect 13320 5652 13326 5664
rect 13556 5624 13584 5664
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 15304 5692 15332 5732
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 16114 5760 16120 5772
rect 15519 5732 16120 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16393 5763 16451 5769
rect 16393 5729 16405 5763
rect 16439 5760 16451 5763
rect 17218 5760 17224 5772
rect 16439 5732 17224 5760
rect 16439 5729 16451 5732
rect 16393 5723 16451 5729
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15304 5664 15945 5692
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 15933 5655 15991 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 17313 5695 17371 5701
rect 17313 5661 17325 5695
rect 17359 5661 17371 5695
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 17313 5655 17371 5661
rect 13096 5596 13584 5624
rect 13630 5584 13636 5636
rect 13688 5624 13694 5636
rect 17328 5624 17356 5655
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 13688 5596 17356 5624
rect 13688 5584 13694 5596
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 5224 5528 6285 5556
rect 5224 5516 5230 5528
rect 6273 5525 6285 5528
rect 6319 5525 6331 5559
rect 6273 5519 6331 5525
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6822 5556 6828 5568
rect 6411 5528 6828 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6822 5516 6828 5528
rect 6880 5556 6886 5568
rect 10229 5559 10287 5565
rect 10229 5556 10241 5559
rect 6880 5528 10241 5556
rect 6880 5516 6886 5528
rect 10229 5525 10241 5528
rect 10275 5556 10287 5559
rect 13648 5556 13676 5584
rect 10275 5528 13676 5556
rect 15289 5559 15347 5565
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 15289 5525 15301 5559
rect 15335 5556 15347 5559
rect 15654 5556 15660 5568
rect 15335 5528 15660 5556
rect 15335 5525 15347 5528
rect 15289 5519 15347 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16114 5556 16120 5568
rect 16075 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 17770 5556 17776 5568
rect 17731 5528 17776 5556
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 1104 5466 21043 5488
rect 1104 5414 5894 5466
rect 5946 5414 5958 5466
rect 6010 5414 6022 5466
rect 6074 5414 6086 5466
rect 6138 5414 6150 5466
rect 6202 5414 10839 5466
rect 10891 5414 10903 5466
rect 10955 5414 10967 5466
rect 11019 5414 11031 5466
rect 11083 5414 11095 5466
rect 11147 5414 15784 5466
rect 15836 5414 15848 5466
rect 15900 5414 15912 5466
rect 15964 5414 15976 5466
rect 16028 5414 16040 5466
rect 16092 5414 20729 5466
rect 20781 5414 20793 5466
rect 20845 5414 20857 5466
rect 20909 5414 20921 5466
rect 20973 5414 20985 5466
rect 21037 5414 21043 5466
rect 1104 5392 21043 5414
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6270 5352 6276 5364
rect 6043 5324 6276 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 7282 5352 7288 5364
rect 7243 5324 7288 5352
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 11793 5355 11851 5361
rect 11793 5321 11805 5355
rect 11839 5352 11851 5355
rect 11974 5352 11980 5364
rect 11839 5324 11980 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13320 5324 13553 5352
rect 13320 5312 13326 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5321 13967 5355
rect 13909 5315 13967 5321
rect 2222 5284 2228 5296
rect 1872 5256 2228 5284
rect 1872 5225 1900 5256
rect 2222 5244 2228 5256
rect 2280 5244 2286 5296
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3007 5256 5856 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2406 5216 2412 5228
rect 2087 5188 2412 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2866 5216 2872 5228
rect 2827 5188 2872 5216
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 5828 5225 5856 5256
rect 6638 5244 6644 5296
rect 6696 5284 6702 5296
rect 6696 5256 7788 5284
rect 6696 5244 6702 5256
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5994 5216 6000 5228
rect 5955 5188 6000 5216
rect 5813 5179 5871 5185
rect 2133 5151 2191 5157
rect 2133 5117 2145 5151
rect 2179 5117 2191 5151
rect 2133 5111 2191 5117
rect 2148 5080 2176 5111
rect 3068 5080 3096 5179
rect 5828 5148 5856 5179
rect 5994 5176 6000 5188
rect 6052 5176 6058 5228
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 6638 5148 6644 5160
rect 5828 5120 6644 5148
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 7484 5148 7512 5179
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 7760 5225 7788 5256
rect 12986 5244 12992 5296
rect 13044 5284 13050 5296
rect 13924 5284 13952 5315
rect 16114 5284 16120 5296
rect 13044 5256 15332 5284
rect 13044 5244 13050 5256
rect 7745 5219 7803 5225
rect 7616 5188 7661 5216
rect 7616 5176 7622 5188
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11296 5188 11713 5216
rect 11296 5176 11302 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 13998 5216 14004 5228
rect 13959 5188 14004 5216
rect 11701 5179 11759 5185
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 14093 5219 14151 5225
rect 14093 5185 14105 5219
rect 14139 5216 14151 5219
rect 14182 5216 14188 5228
rect 14139 5188 14188 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 15010 5216 15016 5228
rect 14971 5188 15016 5216
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15304 5225 15332 5256
rect 15856 5256 16120 5284
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 15562 5216 15568 5228
rect 15335 5188 15568 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 15856 5225 15884 5256
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 16390 5284 16396 5296
rect 16347 5256 16396 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 16390 5244 16396 5256
rect 16448 5244 16454 5296
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 7653 5151 7711 5157
rect 7484 5120 7604 5148
rect 3326 5080 3332 5092
rect 2148 5052 3332 5080
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 7576 5080 7604 5120
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 8018 5148 8024 5160
rect 7699 5120 8024 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 9456 5120 13369 5148
rect 9456 5108 9462 5120
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 7926 5080 7932 5092
rect 7576 5052 7932 5080
rect 7926 5040 7932 5052
rect 7984 5080 7990 5092
rect 9416 5080 9444 5108
rect 7984 5052 9444 5080
rect 13372 5080 13400 5111
rect 15654 5108 15660 5160
rect 15712 5148 15718 5160
rect 16040 5148 16068 5179
rect 15712 5120 16068 5148
rect 15712 5108 15718 5120
rect 17126 5080 17132 5092
rect 13372 5052 17132 5080
rect 7984 5040 7990 5052
rect 17126 5040 17132 5052
rect 17184 5040 17190 5092
rect 1104 4922 20884 4944
rect 1104 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 3550 4922
rect 3602 4870 3614 4922
rect 3666 4870 3678 4922
rect 3730 4870 8367 4922
rect 8419 4870 8431 4922
rect 8483 4870 8495 4922
rect 8547 4870 8559 4922
rect 8611 4870 8623 4922
rect 8675 4870 13312 4922
rect 13364 4870 13376 4922
rect 13428 4870 13440 4922
rect 13492 4870 13504 4922
rect 13556 4870 13568 4922
rect 13620 4870 18257 4922
rect 18309 4870 18321 4922
rect 18373 4870 18385 4922
rect 18437 4870 18449 4922
rect 18501 4870 18513 4922
rect 18565 4870 20884 4922
rect 1104 4848 20884 4870
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10192 4780 10885 4808
rect 10192 4768 10198 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 12802 4808 12808 4820
rect 12763 4780 12808 4808
rect 10873 4771 10931 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13173 4811 13231 4817
rect 13173 4777 13185 4811
rect 13219 4808 13231 4811
rect 13630 4808 13636 4820
rect 13219 4780 13636 4808
rect 13219 4777 13231 4780
rect 13173 4771 13231 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13998 4768 14004 4820
rect 14056 4808 14062 4820
rect 15197 4811 15255 4817
rect 15197 4808 15209 4811
rect 14056 4780 15209 4808
rect 14056 4768 14062 4780
rect 15197 4777 15209 4780
rect 15243 4808 15255 4811
rect 15243 4780 15700 4808
rect 15243 4777 15255 4780
rect 15197 4771 15255 4777
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 7098 4740 7104 4752
rect 6328 4712 7104 4740
rect 6328 4700 6334 4712
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 11974 4700 11980 4752
rect 12032 4700 12038 4752
rect 12986 4700 12992 4752
rect 13044 4700 13050 4752
rect 15562 4740 15568 4752
rect 15523 4712 15568 4740
rect 15562 4700 15568 4712
rect 15620 4700 15626 4752
rect 15672 4740 15700 4780
rect 19242 4740 19248 4752
rect 15672 4712 19248 4740
rect 19242 4700 19248 4712
rect 19300 4700 19306 4752
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 5077 4675 5135 4681
rect 3384 4644 4200 4672
rect 3384 4632 3390 4644
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3200 4576 4077 4604
rect 3200 4564 3206 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4172 4590 4200 4644
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 5994 4672 6000 4684
rect 5123 4644 6000 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 5994 4632 6000 4644
rect 6052 4672 6058 4684
rect 7374 4672 7380 4684
rect 6052 4644 6592 4672
rect 7335 4644 7380 4672
rect 6052 4632 6058 4644
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 4065 4567 4123 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6564 4613 6592 4644
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 10888 4644 11529 4672
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6380 4468 6408 4567
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6825 4607 6883 4613
rect 6696 4576 6741 4604
rect 6696 4564 6702 4576
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 6871 4576 7573 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7926 4604 7932 4616
rect 7708 4576 7753 4604
rect 7887 4576 7932 4604
rect 7708 4564 7714 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 10594 4604 10600 4616
rect 10555 4576 10600 4604
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 10888 4613 10916 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 11992 4672 12020 4700
rect 11839 4644 12020 4672
rect 13004 4672 13032 4700
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 13004 4644 13277 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 13265 4641 13277 4644
rect 13311 4641 13323 4675
rect 13265 4635 13323 4641
rect 15010 4632 15016 4684
rect 15068 4672 15074 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15068 4644 15485 4672
rect 15068 4632 15074 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 15694 4675 15752 4681
rect 15694 4641 15706 4675
rect 15740 4672 15752 4675
rect 16114 4672 16120 4684
rect 15740 4644 16120 4672
rect 15740 4641 15752 4644
rect 15694 4635 15752 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11882 4604 11888 4616
rect 11843 4576 11888 4604
rect 11701 4567 11759 4573
rect 10689 4539 10747 4545
rect 10689 4505 10701 4539
rect 10735 4536 10747 4539
rect 11238 4536 11244 4548
rect 10735 4508 11244 4536
rect 10735 4505 10747 4508
rect 10689 4499 10747 4505
rect 11238 4496 11244 4508
rect 11296 4496 11302 4548
rect 11716 4536 11744 4567
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 12066 4604 12072 4616
rect 12023 4576 12072 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12986 4604 12992 4616
rect 12947 4576 12992 4604
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15672 4576 15853 4604
rect 15672 4548 15700 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 12158 4536 12164 4548
rect 11716 4508 12164 4536
rect 12158 4496 12164 4508
rect 12216 4536 12222 4548
rect 13170 4536 13176 4548
rect 12216 4508 13176 4536
rect 12216 4496 12222 4508
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 15654 4496 15660 4548
rect 15712 4496 15718 4548
rect 14458 4468 14464 4480
rect 6380 4440 14464 4468
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 1104 4378 21043 4400
rect 1104 4326 5894 4378
rect 5946 4326 5958 4378
rect 6010 4326 6022 4378
rect 6074 4326 6086 4378
rect 6138 4326 6150 4378
rect 6202 4326 10839 4378
rect 10891 4326 10903 4378
rect 10955 4326 10967 4378
rect 11019 4326 11031 4378
rect 11083 4326 11095 4378
rect 11147 4326 15784 4378
rect 15836 4326 15848 4378
rect 15900 4326 15912 4378
rect 15964 4326 15976 4378
rect 16028 4326 16040 4378
rect 16092 4326 20729 4378
rect 20781 4326 20793 4378
rect 20845 4326 20857 4378
rect 20909 4326 20921 4378
rect 20973 4326 20985 4378
rect 21037 4326 21043 4378
rect 1104 4304 21043 4326
rect 12897 4267 12955 4273
rect 12897 4233 12909 4267
rect 12943 4264 12955 4267
rect 12986 4264 12992 4276
rect 12943 4236 12992 4264
rect 12943 4233 12955 4236
rect 12897 4227 12955 4233
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 11882 4196 11888 4208
rect 11808 4168 11888 4196
rect 11808 4137 11836 4168
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 12158 4196 12164 4208
rect 11992 4168 12164 4196
rect 11992 4137 12020 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12805 4131 12863 4137
rect 12805 4128 12817 4131
rect 12124 4100 12817 4128
rect 12124 4088 12130 4100
rect 12805 4097 12817 4100
rect 12851 4097 12863 4131
rect 12805 4091 12863 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4128 13047 4131
rect 13170 4128 13176 4140
rect 13035 4100 13176 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 10652 4032 11897 4060
rect 10652 4020 10658 4032
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 11885 4023 11943 4029
rect 1104 3834 20884 3856
rect 1104 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 3550 3834
rect 3602 3782 3614 3834
rect 3666 3782 3678 3834
rect 3730 3782 8367 3834
rect 8419 3782 8431 3834
rect 8483 3782 8495 3834
rect 8547 3782 8559 3834
rect 8611 3782 8623 3834
rect 8675 3782 13312 3834
rect 13364 3782 13376 3834
rect 13428 3782 13440 3834
rect 13492 3782 13504 3834
rect 13556 3782 13568 3834
rect 13620 3782 18257 3834
rect 18309 3782 18321 3834
rect 18373 3782 18385 3834
rect 18437 3782 18449 3834
rect 18501 3782 18513 3834
rect 18565 3782 20884 3834
rect 1104 3760 20884 3782
rect 1104 3290 21043 3312
rect 1104 3238 5894 3290
rect 5946 3238 5958 3290
rect 6010 3238 6022 3290
rect 6074 3238 6086 3290
rect 6138 3238 6150 3290
rect 6202 3238 10839 3290
rect 10891 3238 10903 3290
rect 10955 3238 10967 3290
rect 11019 3238 11031 3290
rect 11083 3238 11095 3290
rect 11147 3238 15784 3290
rect 15836 3238 15848 3290
rect 15900 3238 15912 3290
rect 15964 3238 15976 3290
rect 16028 3238 16040 3290
rect 16092 3238 20729 3290
rect 20781 3238 20793 3290
rect 20845 3238 20857 3290
rect 20909 3238 20921 3290
rect 20973 3238 20985 3290
rect 21037 3238 21043 3290
rect 1104 3216 21043 3238
rect 1104 2746 20884 2768
rect 1104 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 3550 2746
rect 3602 2694 3614 2746
rect 3666 2694 3678 2746
rect 3730 2694 8367 2746
rect 8419 2694 8431 2746
rect 8483 2694 8495 2746
rect 8547 2694 8559 2746
rect 8611 2694 8623 2746
rect 8675 2694 13312 2746
rect 13364 2694 13376 2746
rect 13428 2694 13440 2746
rect 13492 2694 13504 2746
rect 13556 2694 13568 2746
rect 13620 2694 18257 2746
rect 18309 2694 18321 2746
rect 18373 2694 18385 2746
rect 18437 2694 18449 2746
rect 18501 2694 18513 2746
rect 18565 2694 20884 2746
rect 1104 2672 20884 2694
rect 7926 2524 7932 2576
rect 7984 2564 7990 2576
rect 7984 2536 16574 2564
rect 7984 2524 7990 2536
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 8812 2468 12388 2496
rect 8812 2456 8818 2468
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2774 2428 2780 2440
rect 2179 2400 2780 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 5534 2428 5540 2440
rect 4847 2400 5540 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 7466 2428 7472 2440
rect 7427 2400 7472 2428
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 12360 2437 12388 2468
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14148 2400 15025 2428
rect 14148 2388 14154 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 16546 2428 16574 2536
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 16546 2400 17693 2428
rect 15013 2391 15071 2397
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 19886 2428 19892 2440
rect 19847 2400 19892 2428
rect 17681 2391 17739 2397
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 1636 2332 1869 2360
rect 1636 2320 1642 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 4246 2320 4252 2372
rect 4304 2360 4310 2372
rect 4525 2363 4583 2369
rect 4525 2360 4537 2363
rect 4304 2332 4537 2360
rect 4304 2320 4310 2332
rect 4525 2329 4537 2332
rect 4571 2329 4583 2363
rect 4525 2323 4583 2329
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 7193 2363 7251 2369
rect 7193 2360 7205 2363
rect 6972 2332 7205 2360
rect 6972 2320 6978 2332
rect 7193 2329 7205 2332
rect 7239 2329 7251 2363
rect 7193 2323 7251 2329
rect 9582 2320 9588 2372
rect 9640 2360 9646 2372
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 9640 2332 9965 2360
rect 9640 2320 9646 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 9953 2323 10011 2329
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 12308 2332 12633 2360
rect 12308 2320 12314 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 12621 2323 12679 2329
rect 14918 2320 14924 2372
rect 14976 2360 14982 2372
rect 15289 2363 15347 2369
rect 15289 2360 15301 2363
rect 14976 2332 15301 2360
rect 14976 2320 14982 2332
rect 15289 2329 15301 2332
rect 15335 2329 15347 2363
rect 15289 2323 15347 2329
rect 17586 2320 17592 2372
rect 17644 2360 17650 2372
rect 17957 2363 18015 2369
rect 17957 2360 17969 2363
rect 17644 2332 17969 2360
rect 17644 2320 17650 2332
rect 17957 2329 17969 2332
rect 18003 2329 18015 2363
rect 17957 2323 18015 2329
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 20254 2360 20260 2372
rect 20211 2332 20260 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 1104 2202 21043 2224
rect 1104 2150 5894 2202
rect 5946 2150 5958 2202
rect 6010 2150 6022 2202
rect 6074 2150 6086 2202
rect 6138 2150 6150 2202
rect 6202 2150 10839 2202
rect 10891 2150 10903 2202
rect 10955 2150 10967 2202
rect 11019 2150 11031 2202
rect 11083 2150 11095 2202
rect 11147 2150 15784 2202
rect 15836 2150 15848 2202
rect 15900 2150 15912 2202
rect 15964 2150 15976 2202
rect 16028 2150 16040 2202
rect 16092 2150 20729 2202
rect 20781 2150 20793 2202
rect 20845 2150 20857 2202
rect 20909 2150 20921 2202
rect 20973 2150 20985 2202
rect 21037 2150 21043 2202
rect 1104 2128 21043 2150
<< via1 >>
rect 11244 19660 11296 19712
rect 14372 19660 14424 19712
rect 5894 19558 5946 19610
rect 5958 19558 6010 19610
rect 6022 19558 6074 19610
rect 6086 19558 6138 19610
rect 6150 19558 6202 19610
rect 10839 19558 10891 19610
rect 10903 19558 10955 19610
rect 10967 19558 11019 19610
rect 11031 19558 11083 19610
rect 11095 19558 11147 19610
rect 15784 19558 15836 19610
rect 15848 19558 15900 19610
rect 15912 19558 15964 19610
rect 15976 19558 16028 19610
rect 16040 19558 16092 19610
rect 20729 19558 20781 19610
rect 20793 19558 20845 19610
rect 20857 19558 20909 19610
rect 20921 19558 20973 19610
rect 20985 19558 21037 19610
rect 13728 19456 13780 19508
rect 10692 19388 10744 19440
rect 14188 19388 14240 19440
rect 14372 19431 14424 19440
rect 14372 19397 14381 19431
rect 14381 19397 14415 19431
rect 14415 19397 14424 19431
rect 14372 19388 14424 19397
rect 2412 19320 2464 19372
rect 6828 19320 6880 19372
rect 11704 19252 11756 19304
rect 4896 19116 4948 19168
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 16212 19320 16264 19372
rect 18236 19388 18288 19440
rect 19340 19252 19392 19304
rect 14096 19184 14148 19236
rect 16580 19184 16632 19236
rect 14740 19159 14792 19168
rect 14740 19125 14749 19159
rect 14749 19125 14783 19159
rect 14783 19125 14792 19159
rect 14740 19116 14792 19125
rect 15384 19159 15436 19168
rect 15384 19125 15393 19159
rect 15393 19125 15427 19159
rect 15427 19125 15436 19159
rect 15384 19116 15436 19125
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 17500 19116 17552 19168
rect 3422 19014 3474 19066
rect 3486 19014 3538 19066
rect 3550 19014 3602 19066
rect 3614 19014 3666 19066
rect 3678 19014 3730 19066
rect 8367 19014 8419 19066
rect 8431 19014 8483 19066
rect 8495 19014 8547 19066
rect 8559 19014 8611 19066
rect 8623 19014 8675 19066
rect 13312 19014 13364 19066
rect 13376 19014 13428 19066
rect 13440 19014 13492 19066
rect 13504 19014 13556 19066
rect 13568 19014 13620 19066
rect 18257 19014 18309 19066
rect 18321 19014 18373 19066
rect 18385 19014 18437 19066
rect 18449 19014 18501 19066
rect 18513 19014 18565 19066
rect 6828 18912 6880 18964
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 7564 18708 7616 18760
rect 2320 18683 2372 18692
rect 2320 18649 2329 18683
rect 2329 18649 2363 18683
rect 2363 18649 2372 18683
rect 2320 18640 2372 18649
rect 2412 18640 2464 18692
rect 4160 18640 4212 18692
rect 14740 18912 14792 18964
rect 15016 18912 15068 18964
rect 11244 18844 11296 18896
rect 14096 18844 14148 18896
rect 14188 18844 14240 18896
rect 9220 18708 9272 18760
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 14556 18708 14608 18760
rect 2964 18572 3016 18624
rect 13636 18640 13688 18692
rect 14740 18683 14792 18692
rect 14740 18649 14749 18683
rect 14749 18649 14783 18683
rect 14783 18649 14792 18683
rect 14740 18640 14792 18649
rect 13912 18572 13964 18624
rect 15660 18640 15712 18692
rect 17224 18708 17276 18760
rect 16580 18640 16632 18692
rect 17040 18640 17092 18692
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 19340 18640 19392 18692
rect 15200 18572 15252 18624
rect 5894 18470 5946 18522
rect 5958 18470 6010 18522
rect 6022 18470 6074 18522
rect 6086 18470 6138 18522
rect 6150 18470 6202 18522
rect 10839 18470 10891 18522
rect 10903 18470 10955 18522
rect 10967 18470 11019 18522
rect 11031 18470 11083 18522
rect 11095 18470 11147 18522
rect 15784 18470 15836 18522
rect 15848 18470 15900 18522
rect 15912 18470 15964 18522
rect 15976 18470 16028 18522
rect 16040 18470 16092 18522
rect 20729 18470 20781 18522
rect 20793 18470 20845 18522
rect 20857 18470 20909 18522
rect 20921 18470 20973 18522
rect 20985 18470 21037 18522
rect 14740 18368 14792 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 4896 18343 4948 18352
rect 4896 18309 4914 18343
rect 4914 18309 4948 18343
rect 4896 18300 4948 18309
rect 8208 18300 8260 18352
rect 2964 18275 3016 18284
rect 2964 18241 2973 18275
rect 2973 18241 3007 18275
rect 3007 18241 3016 18275
rect 2964 18232 3016 18241
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 16580 18300 16632 18352
rect 17868 18300 17920 18352
rect 5356 18164 5408 18216
rect 9220 18164 9272 18216
rect 11704 18164 11756 18216
rect 3056 18028 3108 18080
rect 6184 18028 6236 18080
rect 13912 18096 13964 18148
rect 14924 18275 14976 18284
rect 14924 18241 14933 18275
rect 14933 18241 14967 18275
rect 14967 18241 14976 18275
rect 14924 18232 14976 18241
rect 15016 18275 15068 18284
rect 15016 18241 15025 18275
rect 15025 18241 15059 18275
rect 15059 18241 15068 18275
rect 15568 18275 15620 18284
rect 15016 18232 15068 18241
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 14832 18028 14884 18080
rect 16672 18232 16724 18284
rect 16948 18232 17000 18284
rect 16212 18164 16264 18216
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 19340 18028 19392 18080
rect 3422 17926 3474 17978
rect 3486 17926 3538 17978
rect 3550 17926 3602 17978
rect 3614 17926 3666 17978
rect 3678 17926 3730 17978
rect 8367 17926 8419 17978
rect 8431 17926 8483 17978
rect 8495 17926 8547 17978
rect 8559 17926 8611 17978
rect 8623 17926 8675 17978
rect 13312 17926 13364 17978
rect 13376 17926 13428 17978
rect 13440 17926 13492 17978
rect 13504 17926 13556 17978
rect 13568 17926 13620 17978
rect 18257 17926 18309 17978
rect 18321 17926 18373 17978
rect 18385 17926 18437 17978
rect 18449 17926 18501 17978
rect 18513 17926 18565 17978
rect 1768 17620 1820 17672
rect 2320 17824 2372 17876
rect 13636 17824 13688 17876
rect 14924 17756 14976 17808
rect 1952 17620 2004 17672
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 3056 17620 3108 17672
rect 5356 17620 5408 17672
rect 7564 17620 7616 17672
rect 6184 17595 6236 17604
rect 6184 17561 6218 17595
rect 6218 17561 6236 17595
rect 6184 17552 6236 17561
rect 14188 17688 14240 17740
rect 15016 17731 15068 17740
rect 15016 17697 15025 17731
rect 15025 17697 15059 17731
rect 15059 17697 15068 17731
rect 15016 17688 15068 17697
rect 15568 17688 15620 17740
rect 17040 17756 17092 17808
rect 13728 17620 13780 17672
rect 16948 17620 17000 17672
rect 15384 17552 15436 17604
rect 15844 17552 15896 17604
rect 16304 17552 16356 17604
rect 16672 17595 16724 17604
rect 16672 17561 16681 17595
rect 16681 17561 16715 17595
rect 16715 17561 16724 17595
rect 16672 17552 16724 17561
rect 17868 17552 17920 17604
rect 19340 17552 19392 17604
rect 19800 17595 19852 17604
rect 19800 17561 19809 17595
rect 19809 17561 19843 17595
rect 19843 17561 19852 17595
rect 19800 17552 19852 17561
rect 1952 17527 2004 17536
rect 1952 17493 1967 17527
rect 1967 17493 2001 17527
rect 2001 17493 2004 17527
rect 1952 17484 2004 17493
rect 3148 17484 3200 17536
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 5894 17382 5946 17434
rect 5958 17382 6010 17434
rect 6022 17382 6074 17434
rect 6086 17382 6138 17434
rect 6150 17382 6202 17434
rect 10839 17382 10891 17434
rect 10903 17382 10955 17434
rect 10967 17382 11019 17434
rect 11031 17382 11083 17434
rect 11095 17382 11147 17434
rect 15784 17382 15836 17434
rect 15848 17382 15900 17434
rect 15912 17382 15964 17434
rect 15976 17382 16028 17434
rect 16040 17382 16092 17434
rect 20729 17382 20781 17434
rect 20793 17382 20845 17434
rect 20857 17382 20909 17434
rect 20921 17382 20973 17434
rect 20985 17382 21037 17434
rect 1952 17144 2004 17196
rect 4252 17144 4304 17196
rect 5356 17144 5408 17196
rect 11152 17144 11204 17196
rect 13728 17144 13780 17196
rect 15384 17144 15436 17196
rect 19524 17144 19576 17196
rect 19708 17144 19760 17196
rect 1860 17119 1912 17128
rect 1860 17085 1869 17119
rect 1869 17085 1903 17119
rect 1903 17085 1912 17119
rect 1860 17076 1912 17085
rect 9220 17076 9272 17128
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 17500 17119 17552 17128
rect 17500 17085 17509 17119
rect 17509 17085 17543 17119
rect 17543 17085 17552 17119
rect 17500 17076 17552 17085
rect 2136 17008 2188 17060
rect 3884 16940 3936 16992
rect 16856 17008 16908 17060
rect 14280 16940 14332 16992
rect 15108 16940 15160 16992
rect 19616 16940 19668 16992
rect 3422 16838 3474 16890
rect 3486 16838 3538 16890
rect 3550 16838 3602 16890
rect 3614 16838 3666 16890
rect 3678 16838 3730 16890
rect 8367 16838 8419 16890
rect 8431 16838 8483 16890
rect 8495 16838 8547 16890
rect 8559 16838 8611 16890
rect 8623 16838 8675 16890
rect 13312 16838 13364 16890
rect 13376 16838 13428 16890
rect 13440 16838 13492 16890
rect 13504 16838 13556 16890
rect 13568 16838 13620 16890
rect 18257 16838 18309 16890
rect 18321 16838 18373 16890
rect 18385 16838 18437 16890
rect 18449 16838 18501 16890
rect 18513 16838 18565 16890
rect 3976 16736 4028 16788
rect 8300 16736 8352 16788
rect 10600 16779 10652 16788
rect 10600 16745 10609 16779
rect 10609 16745 10643 16779
rect 10643 16745 10652 16779
rect 10600 16736 10652 16745
rect 11152 16736 11204 16788
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2780 16668 2832 16720
rect 13636 16668 13688 16720
rect 16580 16668 16632 16720
rect 5448 16600 5500 16652
rect 9220 16643 9272 16652
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 11704 16600 11756 16652
rect 2228 16464 2280 16516
rect 5264 16439 5316 16448
rect 5264 16405 5273 16439
rect 5273 16405 5307 16439
rect 5307 16405 5316 16439
rect 5264 16396 5316 16405
rect 7564 16464 7616 16516
rect 10508 16532 10560 16584
rect 9312 16464 9364 16516
rect 14924 16532 14976 16584
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 16948 16532 17000 16584
rect 18144 16532 18196 16584
rect 19340 16532 19392 16584
rect 19800 16668 19852 16720
rect 19524 16600 19576 16652
rect 19616 16575 19668 16584
rect 19616 16541 19625 16575
rect 19625 16541 19659 16575
rect 19659 16541 19668 16575
rect 19616 16532 19668 16541
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 14740 16464 14792 16516
rect 16580 16507 16632 16516
rect 16580 16473 16589 16507
rect 16589 16473 16623 16507
rect 16623 16473 16632 16507
rect 16580 16464 16632 16473
rect 17408 16507 17460 16516
rect 17408 16473 17417 16507
rect 17417 16473 17451 16507
rect 17451 16473 17460 16507
rect 17408 16464 17460 16473
rect 16856 16396 16908 16448
rect 17684 16439 17736 16448
rect 17684 16405 17693 16439
rect 17693 16405 17727 16439
rect 17727 16405 17736 16439
rect 18052 16464 18104 16516
rect 17684 16396 17736 16405
rect 19524 16396 19576 16448
rect 5894 16294 5946 16346
rect 5958 16294 6010 16346
rect 6022 16294 6074 16346
rect 6086 16294 6138 16346
rect 6150 16294 6202 16346
rect 10839 16294 10891 16346
rect 10903 16294 10955 16346
rect 10967 16294 11019 16346
rect 11031 16294 11083 16346
rect 11095 16294 11147 16346
rect 15784 16294 15836 16346
rect 15848 16294 15900 16346
rect 15912 16294 15964 16346
rect 15976 16294 16028 16346
rect 16040 16294 16092 16346
rect 20729 16294 20781 16346
rect 20793 16294 20845 16346
rect 20857 16294 20909 16346
rect 20921 16294 20973 16346
rect 20985 16294 21037 16346
rect 2228 16235 2280 16244
rect 2228 16201 2237 16235
rect 2237 16201 2271 16235
rect 2271 16201 2280 16235
rect 2228 16192 2280 16201
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 2780 16192 2832 16201
rect 10600 16192 10652 16244
rect 11888 16192 11940 16244
rect 19800 16235 19852 16244
rect 3884 16167 3936 16176
rect 3884 16133 3902 16167
rect 3902 16133 3936 16167
rect 3884 16124 3936 16133
rect 1952 16099 2004 16108
rect 1952 16065 1961 16099
rect 1961 16065 1995 16099
rect 1995 16065 2004 16099
rect 1952 16056 2004 16065
rect 2136 16056 2188 16108
rect 19800 16201 19809 16235
rect 19809 16201 19843 16235
rect 19843 16201 19852 16235
rect 19800 16192 19852 16201
rect 5448 16056 5500 16108
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 6000 16056 6052 16065
rect 7564 16056 7616 16108
rect 9128 16056 9180 16108
rect 11704 16056 11756 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 15568 16056 15620 16108
rect 15200 16031 15252 16040
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 2412 15852 2464 15904
rect 13728 15920 13780 15972
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 17592 16099 17644 16108
rect 17592 16065 17601 16099
rect 17601 16065 17635 16099
rect 17635 16065 17644 16099
rect 17592 16056 17644 16065
rect 17684 16056 17736 16108
rect 16580 15988 16632 16040
rect 17500 15988 17552 16040
rect 9496 15852 9548 15904
rect 15108 15852 15160 15904
rect 16764 15920 16816 15972
rect 17316 15852 17368 15904
rect 19524 16056 19576 16108
rect 19708 16124 19760 16176
rect 19432 16031 19484 16040
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 3422 15750 3474 15802
rect 3486 15750 3538 15802
rect 3550 15750 3602 15802
rect 3614 15750 3666 15802
rect 3678 15750 3730 15802
rect 8367 15750 8419 15802
rect 8431 15750 8483 15802
rect 8495 15750 8547 15802
rect 8559 15750 8611 15802
rect 8623 15750 8675 15802
rect 13312 15750 13364 15802
rect 13376 15750 13428 15802
rect 13440 15750 13492 15802
rect 13504 15750 13556 15802
rect 13568 15750 13620 15802
rect 18257 15750 18309 15802
rect 18321 15750 18373 15802
rect 18385 15750 18437 15802
rect 18449 15750 18501 15802
rect 18513 15750 18565 15802
rect 5632 15648 5684 15700
rect 6000 15648 6052 15700
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 17592 15691 17644 15700
rect 2320 15580 2372 15632
rect 14464 15580 14516 15632
rect 17040 15580 17092 15632
rect 17592 15657 17601 15691
rect 17601 15657 17635 15691
rect 17635 15657 17644 15691
rect 17592 15648 17644 15657
rect 17868 15648 17920 15700
rect 19432 15648 19484 15700
rect 17684 15580 17736 15632
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15292 15512 15344 15564
rect 16948 15512 17000 15564
rect 17868 15512 17920 15564
rect 2412 15444 2464 15496
rect 15108 15444 15160 15496
rect 2504 15376 2556 15428
rect 9588 15376 9640 15428
rect 13636 15376 13688 15428
rect 16672 15376 16724 15428
rect 17316 15376 17368 15428
rect 19524 15376 19576 15428
rect 2044 15308 2096 15360
rect 5894 15206 5946 15258
rect 5958 15206 6010 15258
rect 6022 15206 6074 15258
rect 6086 15206 6138 15258
rect 6150 15206 6202 15258
rect 10839 15206 10891 15258
rect 10903 15206 10955 15258
rect 10967 15206 11019 15258
rect 11031 15206 11083 15258
rect 11095 15206 11147 15258
rect 15784 15206 15836 15258
rect 15848 15206 15900 15258
rect 15912 15206 15964 15258
rect 15976 15206 16028 15258
rect 16040 15206 16092 15258
rect 20729 15206 20781 15258
rect 20793 15206 20845 15258
rect 20857 15206 20909 15258
rect 20921 15206 20973 15258
rect 20985 15206 21037 15258
rect 4160 15104 4212 15156
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 8300 15079 8352 15088
rect 8300 15045 8309 15079
rect 8309 15045 8343 15079
rect 8343 15045 8352 15079
rect 8300 15036 8352 15045
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 9220 14968 9272 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 16948 14968 17000 15020
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 1952 14900 2004 14952
rect 2412 14900 2464 14952
rect 16856 14900 16908 14952
rect 15476 14832 15528 14884
rect 15384 14807 15436 14816
rect 15384 14773 15393 14807
rect 15393 14773 15427 14807
rect 15427 14773 15436 14807
rect 15384 14764 15436 14773
rect 19708 14764 19760 14816
rect 3422 14662 3474 14714
rect 3486 14662 3538 14714
rect 3550 14662 3602 14714
rect 3614 14662 3666 14714
rect 3678 14662 3730 14714
rect 8367 14662 8419 14714
rect 8431 14662 8483 14714
rect 8495 14662 8547 14714
rect 8559 14662 8611 14714
rect 8623 14662 8675 14714
rect 13312 14662 13364 14714
rect 13376 14662 13428 14714
rect 13440 14662 13492 14714
rect 13504 14662 13556 14714
rect 13568 14662 13620 14714
rect 18257 14662 18309 14714
rect 18321 14662 18373 14714
rect 18385 14662 18437 14714
rect 18449 14662 18501 14714
rect 18513 14662 18565 14714
rect 15476 14560 15528 14612
rect 16764 14560 16816 14612
rect 17132 14560 17184 14612
rect 19524 14560 19576 14612
rect 14924 14492 14976 14544
rect 15384 14492 15436 14544
rect 1952 14424 2004 14476
rect 5632 14467 5684 14476
rect 5632 14433 5641 14467
rect 5641 14433 5675 14467
rect 5675 14433 5684 14467
rect 5632 14424 5684 14433
rect 9220 14424 9272 14476
rect 14648 14424 14700 14476
rect 18420 14492 18472 14544
rect 19156 14492 19208 14544
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 5264 14356 5316 14408
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 7932 14356 7984 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 16672 14356 16724 14408
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17776 14399 17828 14408
rect 17040 14356 17092 14365
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 18696 14424 18748 14476
rect 18604 14356 18656 14408
rect 2320 14288 2372 14340
rect 7564 14288 7616 14340
rect 19340 14288 19392 14340
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 8760 14220 8812 14272
rect 14648 14220 14700 14272
rect 14832 14263 14884 14272
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 15200 14220 15252 14272
rect 16120 14220 16172 14272
rect 17316 14263 17368 14272
rect 17316 14229 17325 14263
rect 17325 14229 17359 14263
rect 17359 14229 17368 14263
rect 17316 14220 17368 14229
rect 19524 14220 19576 14272
rect 5894 14118 5946 14170
rect 5958 14118 6010 14170
rect 6022 14118 6074 14170
rect 6086 14118 6138 14170
rect 6150 14118 6202 14170
rect 10839 14118 10891 14170
rect 10903 14118 10955 14170
rect 10967 14118 11019 14170
rect 11031 14118 11083 14170
rect 11095 14118 11147 14170
rect 15784 14118 15836 14170
rect 15848 14118 15900 14170
rect 15912 14118 15964 14170
rect 15976 14118 16028 14170
rect 16040 14118 16092 14170
rect 20729 14118 20781 14170
rect 20793 14118 20845 14170
rect 20857 14118 20909 14170
rect 20921 14118 20973 14170
rect 20985 14118 21037 14170
rect 2412 14016 2464 14068
rect 1860 13880 1912 13932
rect 2412 13880 2464 13932
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2136 13812 2188 13864
rect 3148 13880 3200 13932
rect 3608 13880 3660 13932
rect 2872 13744 2924 13796
rect 3976 13880 4028 13932
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 10140 13923 10192 13932
rect 10140 13889 10158 13923
rect 10158 13889 10192 13923
rect 10140 13880 10192 13889
rect 16580 14016 16632 14068
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 17132 13991 17184 14000
rect 14924 13923 14976 13932
rect 5540 13812 5592 13864
rect 11704 13812 11756 13864
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15292 13880 15344 13932
rect 17132 13957 17141 13991
rect 17141 13957 17175 13991
rect 17175 13957 17184 13991
rect 17132 13948 17184 13957
rect 18420 13991 18472 14000
rect 18420 13957 18429 13991
rect 18429 13957 18463 13991
rect 18463 13957 18472 13991
rect 18420 13948 18472 13957
rect 18604 13991 18656 14000
rect 18604 13957 18629 13991
rect 18629 13957 18656 13991
rect 18604 13948 18656 13957
rect 19524 13923 19576 13932
rect 15200 13812 15252 13864
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 19524 13889 19533 13923
rect 19533 13889 19567 13923
rect 19567 13889 19576 13923
rect 19524 13880 19576 13889
rect 19984 13948 20036 14000
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 3976 13787 4028 13796
rect 3976 13753 3985 13787
rect 3985 13753 4019 13787
rect 4019 13753 4028 13787
rect 3976 13744 4028 13753
rect 14280 13744 14332 13796
rect 15292 13787 15344 13796
rect 15292 13753 15301 13787
rect 15301 13753 15335 13787
rect 15335 13753 15344 13787
rect 15292 13744 15344 13753
rect 17776 13744 17828 13796
rect 15200 13719 15252 13728
rect 15200 13685 15209 13719
rect 15209 13685 15243 13719
rect 15243 13685 15252 13719
rect 15200 13676 15252 13685
rect 17224 13676 17276 13728
rect 19708 13744 19760 13796
rect 18696 13676 18748 13728
rect 3422 13574 3474 13626
rect 3486 13574 3538 13626
rect 3550 13574 3602 13626
rect 3614 13574 3666 13626
rect 3678 13574 3730 13626
rect 8367 13574 8419 13626
rect 8431 13574 8483 13626
rect 8495 13574 8547 13626
rect 8559 13574 8611 13626
rect 8623 13574 8675 13626
rect 13312 13574 13364 13626
rect 13376 13574 13428 13626
rect 13440 13574 13492 13626
rect 13504 13574 13556 13626
rect 13568 13574 13620 13626
rect 18257 13574 18309 13626
rect 18321 13574 18373 13626
rect 18385 13574 18437 13626
rect 18449 13574 18501 13626
rect 18513 13574 18565 13626
rect 5356 13472 5408 13524
rect 17132 13472 17184 13524
rect 19340 13472 19392 13524
rect 19616 13515 19668 13524
rect 19616 13481 19625 13515
rect 19625 13481 19659 13515
rect 19659 13481 19668 13515
rect 19616 13472 19668 13481
rect 2872 13404 2924 13456
rect 4252 13404 4304 13456
rect 19984 13447 20036 13456
rect 19984 13413 19993 13447
rect 19993 13413 20027 13447
rect 20027 13413 20036 13447
rect 19984 13404 20036 13413
rect 3976 13336 4028 13388
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 2320 13268 2372 13320
rect 5540 13268 5592 13320
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 17960 13268 18012 13320
rect 6460 13200 6512 13252
rect 7472 13132 7524 13184
rect 17776 13132 17828 13184
rect 19248 13132 19300 13184
rect 19708 13132 19760 13184
rect 5894 13030 5946 13082
rect 5958 13030 6010 13082
rect 6022 13030 6074 13082
rect 6086 13030 6138 13082
rect 6150 13030 6202 13082
rect 10839 13030 10891 13082
rect 10903 13030 10955 13082
rect 10967 13030 11019 13082
rect 11031 13030 11083 13082
rect 11095 13030 11147 13082
rect 15784 13030 15836 13082
rect 15848 13030 15900 13082
rect 15912 13030 15964 13082
rect 15976 13030 16028 13082
rect 16040 13030 16092 13082
rect 20729 13030 20781 13082
rect 20793 13030 20845 13082
rect 20857 13030 20909 13082
rect 20921 13030 20973 13082
rect 20985 13030 21037 13082
rect 19616 12971 19668 12980
rect 19616 12937 19625 12971
rect 19625 12937 19659 12971
rect 19659 12937 19668 12971
rect 19616 12928 19668 12937
rect 1768 12860 1820 12912
rect 1952 12860 2004 12912
rect 2504 12860 2556 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 5540 12860 5592 12912
rect 17224 12903 17276 12912
rect 17224 12869 17233 12903
rect 17233 12869 17267 12903
rect 17267 12869 17276 12903
rect 17224 12860 17276 12869
rect 17776 12860 17828 12912
rect 19340 12860 19392 12912
rect 4436 12835 4488 12844
rect 4436 12801 4470 12835
rect 4470 12801 4488 12835
rect 4436 12792 4488 12801
rect 7932 12792 7984 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 8852 12724 8904 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 17960 12656 18012 12708
rect 18604 12792 18656 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 18696 12724 18748 12776
rect 19616 12724 19668 12776
rect 19984 12656 20036 12708
rect 5632 12588 5684 12640
rect 11244 12588 11296 12640
rect 14740 12588 14792 12640
rect 15384 12588 15436 12640
rect 18696 12588 18748 12640
rect 3422 12486 3474 12538
rect 3486 12486 3538 12538
rect 3550 12486 3602 12538
rect 3614 12486 3666 12538
rect 3678 12486 3730 12538
rect 8367 12486 8419 12538
rect 8431 12486 8483 12538
rect 8495 12486 8547 12538
rect 8559 12486 8611 12538
rect 8623 12486 8675 12538
rect 13312 12486 13364 12538
rect 13376 12486 13428 12538
rect 13440 12486 13492 12538
rect 13504 12486 13556 12538
rect 13568 12486 13620 12538
rect 18257 12486 18309 12538
rect 18321 12486 18373 12538
rect 18385 12486 18437 12538
rect 18449 12486 18501 12538
rect 18513 12486 18565 12538
rect 11888 12384 11940 12436
rect 15200 12427 15252 12436
rect 1860 12248 1912 12300
rect 1952 12223 2004 12232
rect 1676 12112 1728 12164
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 5540 12180 5592 12232
rect 6552 12180 6604 12232
rect 7932 12180 7984 12232
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 15200 12393 15209 12427
rect 15209 12393 15243 12427
rect 15243 12393 15252 12427
rect 15200 12384 15252 12393
rect 15292 12384 15344 12436
rect 17960 12427 18012 12436
rect 17960 12393 17969 12427
rect 17969 12393 18003 12427
rect 18003 12393 18012 12427
rect 17960 12384 18012 12393
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 19708 12384 19760 12436
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 13820 12248 13872 12300
rect 15568 12316 15620 12368
rect 16212 12316 16264 12368
rect 16120 12223 16172 12232
rect 4252 12044 4304 12096
rect 10600 12112 10652 12164
rect 9680 12044 9732 12096
rect 11612 12044 11664 12096
rect 14740 12112 14792 12164
rect 15108 12112 15160 12164
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 18052 12316 18104 12368
rect 19340 12316 19392 12368
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 16580 12112 16632 12164
rect 17224 12155 17276 12164
rect 17224 12121 17233 12155
rect 17233 12121 17267 12155
rect 17267 12121 17276 12155
rect 17224 12112 17276 12121
rect 15384 12044 15436 12096
rect 17776 12044 17828 12096
rect 19708 12112 19760 12164
rect 19800 12087 19852 12096
rect 19800 12053 19809 12087
rect 19809 12053 19843 12087
rect 19843 12053 19852 12087
rect 19800 12044 19852 12053
rect 5894 11942 5946 11994
rect 5958 11942 6010 11994
rect 6022 11942 6074 11994
rect 6086 11942 6138 11994
rect 6150 11942 6202 11994
rect 10839 11942 10891 11994
rect 10903 11942 10955 11994
rect 10967 11942 11019 11994
rect 11031 11942 11083 11994
rect 11095 11942 11147 11994
rect 15784 11942 15836 11994
rect 15848 11942 15900 11994
rect 15912 11942 15964 11994
rect 15976 11942 16028 11994
rect 16040 11942 16092 11994
rect 20729 11942 20781 11994
rect 20793 11942 20845 11994
rect 20857 11942 20909 11994
rect 20921 11942 20973 11994
rect 20985 11942 21037 11994
rect 1860 11840 1912 11892
rect 14740 11840 14792 11892
rect 15568 11840 15620 11892
rect 18604 11840 18656 11892
rect 19616 11840 19668 11892
rect 19800 11883 19852 11892
rect 19800 11849 19809 11883
rect 19809 11849 19843 11883
rect 19843 11849 19852 11883
rect 19800 11840 19852 11849
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 2412 11704 2464 11756
rect 5540 11704 5592 11756
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 6828 11747 6880 11756
rect 6828 11713 6862 11747
rect 6862 11713 6880 11747
rect 6828 11704 6880 11713
rect 11704 11704 11756 11756
rect 12256 11704 12308 11756
rect 14924 11704 14976 11756
rect 15108 11704 15160 11756
rect 18604 11747 18656 11756
rect 2228 11636 2280 11688
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 18788 11704 18840 11756
rect 1952 11611 2004 11620
rect 1952 11577 1961 11611
rect 1961 11577 1995 11611
rect 1995 11577 2004 11611
rect 1952 11568 2004 11577
rect 15108 11568 15160 11620
rect 15292 11611 15344 11620
rect 15292 11577 15301 11611
rect 15301 11577 15335 11611
rect 15335 11577 15344 11611
rect 15292 11568 15344 11577
rect 16672 11568 16724 11620
rect 17316 11611 17368 11620
rect 17316 11577 17325 11611
rect 17325 11577 17359 11611
rect 17359 11577 17368 11611
rect 17316 11568 17368 11577
rect 19432 11636 19484 11688
rect 19800 11568 19852 11620
rect 7840 11500 7892 11552
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 15660 11500 15712 11552
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 3422 11398 3474 11450
rect 3486 11398 3538 11450
rect 3550 11398 3602 11450
rect 3614 11398 3666 11450
rect 3678 11398 3730 11450
rect 8367 11398 8419 11450
rect 8431 11398 8483 11450
rect 8495 11398 8547 11450
rect 8559 11398 8611 11450
rect 8623 11398 8675 11450
rect 13312 11398 13364 11450
rect 13376 11398 13428 11450
rect 13440 11398 13492 11450
rect 13504 11398 13556 11450
rect 13568 11398 13620 11450
rect 18257 11398 18309 11450
rect 18321 11398 18373 11450
rect 18385 11398 18437 11450
rect 18449 11398 18501 11450
rect 18513 11398 18565 11450
rect 2228 11339 2280 11348
rect 2228 11305 2237 11339
rect 2237 11305 2271 11339
rect 2271 11305 2280 11339
rect 2228 11296 2280 11305
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 6644 11228 6696 11280
rect 15476 11228 15528 11280
rect 18512 11296 18564 11348
rect 19616 11296 19668 11348
rect 17040 11228 17092 11280
rect 11612 11160 11664 11212
rect 12532 11160 12584 11212
rect 17316 11203 17368 11212
rect 1676 11092 1728 11144
rect 1952 11092 2004 11144
rect 2412 11092 2464 11144
rect 5540 11092 5592 11144
rect 5816 11024 5868 11076
rect 15108 11024 15160 11076
rect 17316 11169 17325 11203
rect 17325 11169 17359 11203
rect 17359 11169 17368 11203
rect 17316 11160 17368 11169
rect 17776 11160 17828 11212
rect 16212 11092 16264 11144
rect 16672 11092 16724 11144
rect 18144 11092 18196 11144
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 18512 11024 18564 11076
rect 18604 10999 18656 11008
rect 18604 10965 18613 10999
rect 18613 10965 18647 10999
rect 18647 10965 18656 10999
rect 18604 10956 18656 10965
rect 5894 10854 5946 10906
rect 5958 10854 6010 10906
rect 6022 10854 6074 10906
rect 6086 10854 6138 10906
rect 6150 10854 6202 10906
rect 10839 10854 10891 10906
rect 10903 10854 10955 10906
rect 10967 10854 11019 10906
rect 11031 10854 11083 10906
rect 11095 10854 11147 10906
rect 15784 10854 15836 10906
rect 15848 10854 15900 10906
rect 15912 10854 15964 10906
rect 15976 10854 16028 10906
rect 16040 10854 16092 10906
rect 20729 10854 20781 10906
rect 20793 10854 20845 10906
rect 20857 10854 20909 10906
rect 20921 10854 20973 10906
rect 20985 10854 21037 10906
rect 14924 10752 14976 10804
rect 18512 10795 18564 10804
rect 18512 10761 18521 10795
rect 18521 10761 18555 10795
rect 18555 10761 18564 10795
rect 18512 10752 18564 10761
rect 1952 10684 2004 10736
rect 1860 10616 1912 10668
rect 17132 10727 17184 10736
rect 2872 10616 2924 10668
rect 5540 10616 5592 10668
rect 6552 10616 6604 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 14648 10616 14700 10668
rect 9956 10548 10008 10600
rect 15108 10548 15160 10600
rect 17132 10693 17159 10727
rect 17159 10693 17184 10727
rect 17132 10684 17184 10693
rect 17776 10684 17828 10736
rect 18604 10684 18656 10736
rect 18144 10616 18196 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19892 10684 19944 10736
rect 18604 10548 18656 10600
rect 19156 10548 19208 10600
rect 2688 10480 2740 10532
rect 13728 10480 13780 10532
rect 2412 10412 2464 10464
rect 2780 10412 2832 10464
rect 11612 10412 11664 10464
rect 14556 10412 14608 10464
rect 14924 10412 14976 10464
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 17960 10412 18012 10464
rect 19248 10455 19300 10464
rect 19248 10421 19257 10455
rect 19257 10421 19291 10455
rect 19291 10421 19300 10455
rect 19248 10412 19300 10421
rect 3422 10310 3474 10362
rect 3486 10310 3538 10362
rect 3550 10310 3602 10362
rect 3614 10310 3666 10362
rect 3678 10310 3730 10362
rect 8367 10310 8419 10362
rect 8431 10310 8483 10362
rect 8495 10310 8547 10362
rect 8559 10310 8611 10362
rect 8623 10310 8675 10362
rect 13312 10310 13364 10362
rect 13376 10310 13428 10362
rect 13440 10310 13492 10362
rect 13504 10310 13556 10362
rect 13568 10310 13620 10362
rect 18257 10310 18309 10362
rect 18321 10310 18373 10362
rect 18385 10310 18437 10362
rect 18449 10310 18501 10362
rect 18513 10310 18565 10362
rect 2872 10208 2924 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 15292 10208 15344 10260
rect 15568 10208 15620 10260
rect 18144 10208 18196 10260
rect 1952 10004 2004 10056
rect 15108 10140 15160 10192
rect 12256 10072 12308 10124
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 7748 10047 7800 10056
rect 2780 10004 2832 10013
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 16856 10140 16908 10192
rect 18144 10072 18196 10124
rect 19432 10072 19484 10124
rect 2688 9936 2740 9988
rect 9588 9936 9640 9988
rect 13912 9936 13964 9988
rect 18052 10004 18104 10056
rect 1860 9868 1912 9920
rect 2228 9868 2280 9920
rect 7932 9868 7984 9920
rect 15016 9911 15068 9920
rect 15016 9877 15025 9911
rect 15025 9877 15059 9911
rect 15059 9877 15068 9911
rect 15016 9868 15068 9877
rect 15200 9868 15252 9920
rect 17224 9911 17276 9920
rect 17224 9877 17233 9911
rect 17233 9877 17267 9911
rect 17267 9877 17276 9911
rect 17224 9868 17276 9877
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 19708 10004 19760 10056
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 17408 9868 17460 9877
rect 19156 9868 19208 9920
rect 19432 9911 19484 9920
rect 19432 9877 19441 9911
rect 19441 9877 19475 9911
rect 19475 9877 19484 9911
rect 19432 9868 19484 9877
rect 5894 9766 5946 9818
rect 5958 9766 6010 9818
rect 6022 9766 6074 9818
rect 6086 9766 6138 9818
rect 6150 9766 6202 9818
rect 10839 9766 10891 9818
rect 10903 9766 10955 9818
rect 10967 9766 11019 9818
rect 11031 9766 11083 9818
rect 11095 9766 11147 9818
rect 15784 9766 15836 9818
rect 15848 9766 15900 9818
rect 15912 9766 15964 9818
rect 15976 9766 16028 9818
rect 16040 9766 16092 9818
rect 20729 9766 20781 9818
rect 20793 9766 20845 9818
rect 20857 9766 20909 9818
rect 20921 9766 20973 9818
rect 20985 9766 21037 9818
rect 14924 9664 14976 9716
rect 15384 9664 15436 9716
rect 17224 9664 17276 9716
rect 13728 9596 13780 9648
rect 17960 9639 18012 9648
rect 17960 9605 17969 9639
rect 17969 9605 18003 9639
rect 18003 9605 18012 9639
rect 17960 9596 18012 9605
rect 19432 9596 19484 9648
rect 4620 9571 4672 9580
rect 4620 9537 4638 9571
rect 4638 9537 4672 9571
rect 4620 9528 4672 9537
rect 5724 9528 5776 9580
rect 6552 9528 6604 9580
rect 8024 9571 8076 9580
rect 8024 9537 8058 9571
rect 8058 9537 8076 9571
rect 9772 9571 9824 9580
rect 8024 9528 8076 9537
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 11980 9528 12032 9580
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 14096 9528 14148 9580
rect 14740 9528 14792 9580
rect 17224 9528 17276 9580
rect 17316 9528 17368 9580
rect 17500 9528 17552 9580
rect 18144 9528 18196 9580
rect 18880 9528 18932 9580
rect 19248 9528 19300 9580
rect 19616 9571 19668 9580
rect 19616 9537 19625 9571
rect 19625 9537 19659 9571
rect 19659 9537 19668 9571
rect 19616 9528 19668 9537
rect 19892 9528 19944 9580
rect 15200 9503 15252 9512
rect 2780 9324 2832 9376
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 15292 9460 15344 9512
rect 19800 9392 19852 9444
rect 11888 9324 11940 9376
rect 12992 9324 13044 9376
rect 15292 9324 15344 9376
rect 3422 9222 3474 9274
rect 3486 9222 3538 9274
rect 3550 9222 3602 9274
rect 3614 9222 3666 9274
rect 3678 9222 3730 9274
rect 8367 9222 8419 9274
rect 8431 9222 8483 9274
rect 8495 9222 8547 9274
rect 8559 9222 8611 9274
rect 8623 9222 8675 9274
rect 13312 9222 13364 9274
rect 13376 9222 13428 9274
rect 13440 9222 13492 9274
rect 13504 9222 13556 9274
rect 13568 9222 13620 9274
rect 18257 9222 18309 9274
rect 18321 9222 18373 9274
rect 18385 9222 18437 9274
rect 18449 9222 18501 9274
rect 18513 9222 18565 9274
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 7748 9120 7800 9172
rect 13820 9120 13872 9172
rect 14464 9120 14516 9172
rect 14924 9120 14976 9172
rect 15016 9120 15068 9172
rect 17224 9163 17276 9172
rect 17224 9129 17233 9163
rect 17233 9129 17267 9163
rect 17267 9129 17276 9163
rect 17224 9120 17276 9129
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 19892 9163 19944 9172
rect 19892 9129 19901 9163
rect 19901 9129 19935 9163
rect 19935 9129 19944 9163
rect 19892 9120 19944 9129
rect 2688 9052 2740 9104
rect 3148 8916 3200 8968
rect 4068 8916 4120 8968
rect 4436 8916 4488 8968
rect 5724 8916 5776 8968
rect 14740 9052 14792 9104
rect 17040 9052 17092 9104
rect 17316 9052 17368 9104
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 12256 8916 12308 8968
rect 8116 8848 8168 8900
rect 10692 8848 10744 8900
rect 11612 8848 11664 8900
rect 12808 8848 12860 8900
rect 14832 8916 14884 8968
rect 19156 8984 19208 9036
rect 19248 8916 19300 8968
rect 17040 8891 17092 8900
rect 17040 8857 17049 8891
rect 17049 8857 17083 8891
rect 17083 8857 17092 8891
rect 17040 8848 17092 8857
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 4344 8780 4396 8832
rect 9128 8780 9180 8832
rect 14464 8780 14516 8832
rect 14556 8780 14608 8832
rect 15016 8780 15068 8832
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 16764 8780 16816 8832
rect 5894 8678 5946 8730
rect 5958 8678 6010 8730
rect 6022 8678 6074 8730
rect 6086 8678 6138 8730
rect 6150 8678 6202 8730
rect 10839 8678 10891 8730
rect 10903 8678 10955 8730
rect 10967 8678 11019 8730
rect 11031 8678 11083 8730
rect 11095 8678 11147 8730
rect 15784 8678 15836 8730
rect 15848 8678 15900 8730
rect 15912 8678 15964 8730
rect 15976 8678 16028 8730
rect 16040 8678 16092 8730
rect 20729 8678 20781 8730
rect 20793 8678 20845 8730
rect 20857 8678 20909 8730
rect 20921 8678 20973 8730
rect 20985 8678 21037 8730
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 5816 8576 5868 8628
rect 6828 8576 6880 8628
rect 7564 8576 7616 8628
rect 10692 8576 10744 8628
rect 10876 8576 10928 8628
rect 14740 8619 14792 8628
rect 14740 8585 14749 8619
rect 14749 8585 14783 8619
rect 14783 8585 14792 8619
rect 14740 8576 14792 8585
rect 15016 8576 15068 8628
rect 3148 8508 3200 8560
rect 8852 8551 8904 8560
rect 8852 8517 8861 8551
rect 8861 8517 8895 8551
rect 8895 8517 8904 8551
rect 8852 8508 8904 8517
rect 9864 8508 9916 8560
rect 10324 8508 10376 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 5540 8440 5592 8492
rect 5724 8440 5776 8492
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 4068 8372 4120 8424
rect 4344 8415 4396 8424
rect 4344 8381 4353 8415
rect 4353 8381 4387 8415
rect 4387 8381 4396 8415
rect 4344 8372 4396 8381
rect 4528 8372 4580 8424
rect 5448 8372 5500 8424
rect 6184 8372 6236 8424
rect 7656 8440 7708 8492
rect 8116 8440 8168 8492
rect 8208 8372 8260 8424
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 10416 8440 10468 8492
rect 10876 8440 10928 8492
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 11704 8508 11756 8560
rect 12072 8551 12124 8560
rect 12072 8517 12081 8551
rect 12081 8517 12115 8551
rect 12115 8517 12124 8551
rect 12072 8508 12124 8517
rect 12440 8440 12492 8492
rect 15108 8508 15160 8560
rect 15476 8508 15528 8560
rect 15016 8483 15068 8492
rect 11336 8372 11388 8424
rect 11888 8372 11940 8424
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 17040 8576 17092 8628
rect 17132 8576 17184 8628
rect 19616 8576 19668 8628
rect 17408 8508 17460 8560
rect 16764 8440 16816 8492
rect 17132 8440 17184 8492
rect 17960 8440 18012 8492
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 9588 8304 9640 8356
rect 11244 8304 11296 8356
rect 12072 8304 12124 8356
rect 14648 8372 14700 8424
rect 9036 8279 9088 8288
rect 9036 8245 9045 8279
rect 9045 8245 9079 8279
rect 9079 8245 9088 8279
rect 9036 8236 9088 8245
rect 10048 8236 10100 8288
rect 11888 8279 11940 8288
rect 11888 8245 11897 8279
rect 11897 8245 11931 8279
rect 11931 8245 11940 8279
rect 11888 8236 11940 8245
rect 12716 8279 12768 8288
rect 12716 8245 12725 8279
rect 12725 8245 12759 8279
rect 12759 8245 12768 8279
rect 12716 8236 12768 8245
rect 16120 8304 16172 8356
rect 17040 8304 17092 8356
rect 18144 8372 18196 8424
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 13912 8236 13964 8288
rect 16948 8236 17000 8288
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 3550 8134 3602 8186
rect 3614 8134 3666 8186
rect 3678 8134 3730 8186
rect 8367 8134 8419 8186
rect 8431 8134 8483 8186
rect 8495 8134 8547 8186
rect 8559 8134 8611 8186
rect 8623 8134 8675 8186
rect 13312 8134 13364 8186
rect 13376 8134 13428 8186
rect 13440 8134 13492 8186
rect 13504 8134 13556 8186
rect 13568 8134 13620 8186
rect 18257 8134 18309 8186
rect 18321 8134 18373 8186
rect 18385 8134 18437 8186
rect 18449 8134 18501 8186
rect 18513 8134 18565 8186
rect 6460 8032 6512 8084
rect 8024 8032 8076 8084
rect 9036 8032 9088 8084
rect 11152 8032 11204 8084
rect 12716 8032 12768 8084
rect 4436 7964 4488 8016
rect 11980 7964 12032 8016
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 7656 7896 7708 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 4528 7828 4580 7880
rect 5172 7828 5224 7880
rect 5724 7828 5776 7880
rect 5816 7828 5868 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 5356 7760 5408 7812
rect 5448 7760 5500 7812
rect 8116 7828 8168 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 14188 8032 14240 8084
rect 16948 8032 17000 8084
rect 14188 7896 14240 7948
rect 15568 7896 15620 7948
rect 16580 7896 16632 7948
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 17776 7896 17828 7948
rect 11704 7828 11756 7880
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 13912 7828 13964 7880
rect 14924 7828 14976 7880
rect 15108 7828 15160 7880
rect 2596 7692 2648 7744
rect 6736 7692 6788 7744
rect 11244 7760 11296 7812
rect 11888 7760 11940 7812
rect 15016 7760 15068 7812
rect 9772 7692 9824 7744
rect 10232 7692 10284 7744
rect 12256 7692 12308 7744
rect 17408 7828 17460 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 19248 7828 19300 7880
rect 19340 7760 19392 7812
rect 16856 7735 16908 7744
rect 16856 7701 16865 7735
rect 16865 7701 16899 7735
rect 16899 7701 16908 7735
rect 16856 7692 16908 7701
rect 16948 7692 17000 7744
rect 19616 7735 19668 7744
rect 19616 7701 19643 7735
rect 19643 7701 19668 7735
rect 19616 7692 19668 7701
rect 5894 7590 5946 7642
rect 5958 7590 6010 7642
rect 6022 7590 6074 7642
rect 6086 7590 6138 7642
rect 6150 7590 6202 7642
rect 10839 7590 10891 7642
rect 10903 7590 10955 7642
rect 10967 7590 11019 7642
rect 11031 7590 11083 7642
rect 11095 7590 11147 7642
rect 15784 7590 15836 7642
rect 15848 7590 15900 7642
rect 15912 7590 15964 7642
rect 15976 7590 16028 7642
rect 16040 7590 16092 7642
rect 20729 7590 20781 7642
rect 20793 7590 20845 7642
rect 20857 7590 20909 7642
rect 20921 7590 20973 7642
rect 20985 7590 21037 7642
rect 4068 7531 4120 7540
rect 4068 7497 4077 7531
rect 4077 7497 4111 7531
rect 4111 7497 4120 7531
rect 4068 7488 4120 7497
rect 4528 7488 4580 7540
rect 5540 7488 5592 7540
rect 1952 7352 2004 7404
rect 2228 7352 2280 7404
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 5356 7420 5408 7472
rect 7656 7420 7708 7472
rect 10416 7488 10468 7540
rect 10232 7463 10284 7472
rect 10232 7429 10241 7463
rect 10241 7429 10275 7463
rect 10275 7429 10284 7463
rect 10232 7420 10284 7429
rect 12256 7420 12308 7472
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 4344 7284 4396 7336
rect 4896 7284 4948 7336
rect 3148 7216 3200 7268
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 2320 7148 2372 7200
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6276 7352 6328 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 5080 7216 5132 7268
rect 9404 7284 9456 7336
rect 16948 7488 17000 7540
rect 17132 7488 17184 7540
rect 12532 7420 12584 7472
rect 15568 7420 15620 7472
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 15016 7395 15068 7404
rect 13728 7327 13780 7336
rect 13728 7293 13737 7327
rect 13737 7293 13771 7327
rect 13771 7293 13780 7327
rect 13728 7284 13780 7293
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 15660 7352 15712 7404
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 19616 7488 19668 7540
rect 17316 7420 17368 7472
rect 17868 7420 17920 7472
rect 17684 7352 17736 7404
rect 10048 7259 10100 7268
rect 10048 7225 10057 7259
rect 10057 7225 10091 7259
rect 10091 7225 10100 7259
rect 10048 7216 10100 7225
rect 12072 7216 12124 7268
rect 5540 7148 5592 7200
rect 11612 7148 11664 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 16764 7284 16816 7336
rect 18696 7352 18748 7404
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 18144 7284 18196 7336
rect 14280 7148 14332 7200
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 17868 7216 17920 7268
rect 19708 7148 19760 7200
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 3550 7046 3602 7098
rect 3614 7046 3666 7098
rect 3678 7046 3730 7098
rect 8367 7046 8419 7098
rect 8431 7046 8483 7098
rect 8495 7046 8547 7098
rect 8559 7046 8611 7098
rect 8623 7046 8675 7098
rect 13312 7046 13364 7098
rect 13376 7046 13428 7098
rect 13440 7046 13492 7098
rect 13504 7046 13556 7098
rect 13568 7046 13620 7098
rect 18257 7046 18309 7098
rect 18321 7046 18373 7098
rect 18385 7046 18437 7098
rect 18449 7046 18501 7098
rect 18513 7046 18565 7098
rect 5172 6987 5224 6996
rect 5172 6953 5181 6987
rect 5181 6953 5215 6987
rect 5215 6953 5224 6987
rect 5172 6944 5224 6953
rect 12900 6944 12952 6996
rect 6460 6919 6512 6928
rect 6460 6885 6469 6919
rect 6469 6885 6503 6919
rect 6503 6885 6512 6919
rect 6460 6876 6512 6885
rect 11704 6919 11756 6928
rect 11704 6885 11713 6919
rect 11713 6885 11747 6919
rect 11747 6885 11756 6919
rect 11704 6876 11756 6885
rect 12256 6919 12308 6928
rect 12256 6885 12265 6919
rect 12265 6885 12299 6919
rect 12299 6885 12308 6919
rect 12256 6876 12308 6885
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 5908 6808 5960 6860
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 12716 6808 12768 6860
rect 13728 6876 13780 6928
rect 7656 6783 7708 6792
rect 1952 6672 2004 6724
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 7564 6672 7616 6724
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 10416 6740 10468 6792
rect 8024 6672 8076 6724
rect 8944 6672 8996 6724
rect 3700 6604 3752 6656
rect 7748 6604 7800 6656
rect 9956 6604 10008 6656
rect 10692 6604 10744 6656
rect 11796 6740 11848 6792
rect 12440 6740 12492 6792
rect 11244 6672 11296 6724
rect 12992 6715 13044 6724
rect 12992 6681 13001 6715
rect 13001 6681 13035 6715
rect 13035 6681 13044 6715
rect 12992 6672 13044 6681
rect 13912 6740 13964 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 16212 6876 16264 6928
rect 16396 6740 16448 6792
rect 17316 6740 17368 6792
rect 17500 6740 17552 6792
rect 17592 6740 17644 6792
rect 18052 6783 18104 6792
rect 18052 6749 18061 6783
rect 18061 6749 18095 6783
rect 18095 6749 18104 6783
rect 18052 6740 18104 6749
rect 15016 6715 15068 6724
rect 11980 6604 12032 6656
rect 12072 6604 12124 6656
rect 12532 6604 12584 6656
rect 13728 6604 13780 6656
rect 15016 6681 15025 6715
rect 15025 6681 15059 6715
rect 15059 6681 15068 6715
rect 15016 6672 15068 6681
rect 15660 6604 15712 6656
rect 18604 6604 18656 6656
rect 5894 6502 5946 6554
rect 5958 6502 6010 6554
rect 6022 6502 6074 6554
rect 6086 6502 6138 6554
rect 6150 6502 6202 6554
rect 10839 6502 10891 6554
rect 10903 6502 10955 6554
rect 10967 6502 11019 6554
rect 11031 6502 11083 6554
rect 11095 6502 11147 6554
rect 15784 6502 15836 6554
rect 15848 6502 15900 6554
rect 15912 6502 15964 6554
rect 15976 6502 16028 6554
rect 16040 6502 16092 6554
rect 20729 6502 20781 6554
rect 20793 6502 20845 6554
rect 20857 6502 20909 6554
rect 20921 6502 20973 6554
rect 20985 6502 21037 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 6460 6400 6512 6452
rect 8944 6400 8996 6452
rect 9220 6400 9272 6452
rect 5172 6332 5224 6384
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 5816 6307 5868 6316
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6276 6332 6328 6384
rect 7656 6332 7708 6384
rect 8852 6332 8904 6384
rect 6828 6307 6880 6316
rect 3700 6196 3752 6205
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 7104 6196 7156 6248
rect 8208 6264 8260 6316
rect 9496 6332 9548 6384
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 11336 6400 11388 6452
rect 11980 6400 12032 6452
rect 13176 6400 13228 6452
rect 13728 6400 13780 6452
rect 8024 6196 8076 6248
rect 9956 6196 10008 6248
rect 10232 6264 10284 6316
rect 16304 6332 16356 6384
rect 11244 6264 11296 6316
rect 11612 6264 11664 6316
rect 11796 6264 11848 6316
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 17500 6400 17552 6452
rect 18052 6443 18104 6452
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 19340 6443 19392 6452
rect 19340 6409 19349 6443
rect 19349 6409 19383 6443
rect 19383 6409 19392 6443
rect 19340 6400 19392 6409
rect 17316 6332 17368 6384
rect 11980 6264 12032 6273
rect 10692 6196 10744 6248
rect 2412 6128 2464 6180
rect 7564 6128 7616 6180
rect 10048 6128 10100 6180
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 13084 6196 13136 6248
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 15292 6196 15344 6248
rect 16488 6264 16540 6316
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 18144 6264 18196 6316
rect 18604 6264 18656 6316
rect 19892 6196 19944 6248
rect 4252 6103 4304 6112
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 8208 6060 8260 6112
rect 9496 6060 9548 6112
rect 10784 6060 10836 6112
rect 11336 6060 11388 6112
rect 12072 6060 12124 6112
rect 12992 6060 13044 6112
rect 13820 6128 13872 6180
rect 16304 6128 16356 6180
rect 16672 6128 16724 6180
rect 17592 6060 17644 6112
rect 17868 6103 17920 6112
rect 17868 6069 17877 6103
rect 17877 6069 17911 6103
rect 17911 6069 17920 6103
rect 17868 6060 17920 6069
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 3550 5958 3602 6010
rect 3614 5958 3666 6010
rect 3678 5958 3730 6010
rect 8367 5958 8419 6010
rect 8431 5958 8483 6010
rect 8495 5958 8547 6010
rect 8559 5958 8611 6010
rect 8623 5958 8675 6010
rect 13312 5958 13364 6010
rect 13376 5958 13428 6010
rect 13440 5958 13492 6010
rect 13504 5958 13556 6010
rect 13568 5958 13620 6010
rect 18257 5958 18309 6010
rect 18321 5958 18373 6010
rect 18385 5958 18437 6010
rect 18449 5958 18501 6010
rect 18513 5958 18565 6010
rect 3976 5856 4028 5908
rect 10600 5856 10652 5908
rect 12900 5899 12952 5908
rect 12900 5865 12909 5899
rect 12909 5865 12943 5899
rect 12943 5865 12952 5899
rect 12900 5856 12952 5865
rect 13636 5856 13688 5908
rect 5356 5788 5408 5840
rect 8116 5788 8168 5840
rect 10784 5831 10836 5840
rect 10784 5797 10793 5831
rect 10793 5797 10827 5831
rect 10827 5797 10836 5831
rect 10784 5788 10836 5797
rect 4252 5720 4304 5772
rect 2228 5652 2280 5704
rect 2412 5652 2464 5704
rect 2872 5652 2924 5704
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 6276 5652 6328 5704
rect 7380 5652 7432 5704
rect 13084 5720 13136 5772
rect 15292 5788 15344 5840
rect 18604 5788 18656 5840
rect 8300 5652 8352 5704
rect 8852 5652 8904 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9956 5652 10008 5704
rect 10048 5652 10100 5704
rect 7288 5584 7340 5636
rect 10416 5652 10468 5704
rect 15108 5720 15160 5772
rect 11336 5584 11388 5636
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 14188 5652 14240 5704
rect 16120 5720 16172 5772
rect 17224 5720 17276 5772
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 17592 5695 17644 5704
rect 13636 5584 13688 5636
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 5172 5516 5224 5568
rect 6828 5516 6880 5568
rect 15660 5516 15712 5568
rect 16120 5559 16172 5568
rect 16120 5525 16129 5559
rect 16129 5525 16163 5559
rect 16163 5525 16172 5559
rect 16120 5516 16172 5525
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 5894 5414 5946 5466
rect 5958 5414 6010 5466
rect 6022 5414 6074 5466
rect 6086 5414 6138 5466
rect 6150 5414 6202 5466
rect 10839 5414 10891 5466
rect 10903 5414 10955 5466
rect 10967 5414 11019 5466
rect 11031 5414 11083 5466
rect 11095 5414 11147 5466
rect 15784 5414 15836 5466
rect 15848 5414 15900 5466
rect 15912 5414 15964 5466
rect 15976 5414 16028 5466
rect 16040 5414 16092 5466
rect 20729 5414 20781 5466
rect 20793 5414 20845 5466
rect 20857 5414 20909 5466
rect 20921 5414 20973 5466
rect 20985 5414 21037 5466
rect 6276 5312 6328 5364
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 11980 5312 12032 5364
rect 13268 5312 13320 5364
rect 2228 5244 2280 5296
rect 2412 5176 2464 5228
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 6644 5244 6696 5296
rect 6000 5219 6052 5228
rect 6000 5185 6009 5219
rect 6009 5185 6043 5219
rect 6043 5185 6052 5219
rect 6000 5176 6052 5185
rect 6644 5108 6696 5160
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 12992 5244 13044 5296
rect 7564 5176 7616 5185
rect 11244 5176 11296 5228
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 14188 5176 14240 5228
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 15568 5176 15620 5228
rect 16120 5244 16172 5296
rect 16396 5244 16448 5296
rect 3332 5040 3384 5092
rect 8024 5108 8076 5160
rect 9404 5108 9456 5160
rect 7932 5040 7984 5092
rect 15660 5108 15712 5160
rect 17132 5040 17184 5092
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 3550 4870 3602 4922
rect 3614 4870 3666 4922
rect 3678 4870 3730 4922
rect 8367 4870 8419 4922
rect 8431 4870 8483 4922
rect 8495 4870 8547 4922
rect 8559 4870 8611 4922
rect 8623 4870 8675 4922
rect 13312 4870 13364 4922
rect 13376 4870 13428 4922
rect 13440 4870 13492 4922
rect 13504 4870 13556 4922
rect 13568 4870 13620 4922
rect 18257 4870 18309 4922
rect 18321 4870 18373 4922
rect 18385 4870 18437 4922
rect 18449 4870 18501 4922
rect 18513 4870 18565 4922
rect 10140 4768 10192 4820
rect 12808 4811 12860 4820
rect 12808 4777 12817 4811
rect 12817 4777 12851 4811
rect 12851 4777 12860 4811
rect 12808 4768 12860 4777
rect 13636 4768 13688 4820
rect 14004 4768 14056 4820
rect 6276 4700 6328 4752
rect 7104 4700 7156 4752
rect 11980 4700 12032 4752
rect 12992 4700 13044 4752
rect 15568 4743 15620 4752
rect 15568 4709 15577 4743
rect 15577 4709 15611 4743
rect 15611 4709 15620 4743
rect 15568 4700 15620 4709
rect 19248 4700 19300 4752
rect 3332 4632 3384 4684
rect 3148 4564 3200 4616
rect 6000 4632 6052 4684
rect 7380 4675 7432 4684
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7932 4607 7984 4616
rect 7656 4564 7708 4573
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 15016 4632 15068 4684
rect 16120 4632 16172 4684
rect 11888 4607 11940 4616
rect 11244 4496 11296 4548
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 12072 4564 12124 4616
rect 12992 4607 13044 4616
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 12164 4496 12216 4548
rect 13176 4496 13228 4548
rect 15660 4496 15712 4548
rect 14464 4428 14516 4480
rect 5894 4326 5946 4378
rect 5958 4326 6010 4378
rect 6022 4326 6074 4378
rect 6086 4326 6138 4378
rect 6150 4326 6202 4378
rect 10839 4326 10891 4378
rect 10903 4326 10955 4378
rect 10967 4326 11019 4378
rect 11031 4326 11083 4378
rect 11095 4326 11147 4378
rect 15784 4326 15836 4378
rect 15848 4326 15900 4378
rect 15912 4326 15964 4378
rect 15976 4326 16028 4378
rect 16040 4326 16092 4378
rect 20729 4326 20781 4378
rect 20793 4326 20845 4378
rect 20857 4326 20909 4378
rect 20921 4326 20973 4378
rect 20985 4326 21037 4378
rect 12992 4224 13044 4276
rect 11888 4156 11940 4208
rect 12164 4156 12216 4208
rect 12072 4088 12124 4140
rect 13176 4088 13228 4140
rect 10600 4020 10652 4072
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 3550 3782 3602 3834
rect 3614 3782 3666 3834
rect 3678 3782 3730 3834
rect 8367 3782 8419 3834
rect 8431 3782 8483 3834
rect 8495 3782 8547 3834
rect 8559 3782 8611 3834
rect 8623 3782 8675 3834
rect 13312 3782 13364 3834
rect 13376 3782 13428 3834
rect 13440 3782 13492 3834
rect 13504 3782 13556 3834
rect 13568 3782 13620 3834
rect 18257 3782 18309 3834
rect 18321 3782 18373 3834
rect 18385 3782 18437 3834
rect 18449 3782 18501 3834
rect 18513 3782 18565 3834
rect 5894 3238 5946 3290
rect 5958 3238 6010 3290
rect 6022 3238 6074 3290
rect 6086 3238 6138 3290
rect 6150 3238 6202 3290
rect 10839 3238 10891 3290
rect 10903 3238 10955 3290
rect 10967 3238 11019 3290
rect 11031 3238 11083 3290
rect 11095 3238 11147 3290
rect 15784 3238 15836 3290
rect 15848 3238 15900 3290
rect 15912 3238 15964 3290
rect 15976 3238 16028 3290
rect 16040 3238 16092 3290
rect 20729 3238 20781 3290
rect 20793 3238 20845 3290
rect 20857 3238 20909 3290
rect 20921 3238 20973 3290
rect 20985 3238 21037 3290
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 3550 2694 3602 2746
rect 3614 2694 3666 2746
rect 3678 2694 3730 2746
rect 8367 2694 8419 2746
rect 8431 2694 8483 2746
rect 8495 2694 8547 2746
rect 8559 2694 8611 2746
rect 8623 2694 8675 2746
rect 13312 2694 13364 2746
rect 13376 2694 13428 2746
rect 13440 2694 13492 2746
rect 13504 2694 13556 2746
rect 13568 2694 13620 2746
rect 18257 2694 18309 2746
rect 18321 2694 18373 2746
rect 18385 2694 18437 2746
rect 18449 2694 18501 2746
rect 18513 2694 18565 2746
rect 7932 2524 7984 2576
rect 8760 2456 8812 2508
rect 2780 2388 2832 2440
rect 5540 2388 5592 2440
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 14096 2388 14148 2440
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 1584 2320 1636 2372
rect 4252 2320 4304 2372
rect 6920 2320 6972 2372
rect 9588 2320 9640 2372
rect 12256 2320 12308 2372
rect 14924 2320 14976 2372
rect 17592 2320 17644 2372
rect 20260 2320 20312 2372
rect 5894 2150 5946 2202
rect 5958 2150 6010 2202
rect 6022 2150 6074 2202
rect 6086 2150 6138 2202
rect 6150 2150 6202 2202
rect 10839 2150 10891 2202
rect 10903 2150 10955 2202
rect 10967 2150 11019 2202
rect 11031 2150 11083 2202
rect 11095 2150 11147 2202
rect 15784 2150 15836 2202
rect 15848 2150 15900 2202
rect 15912 2150 15964 2202
rect 15976 2150 16028 2202
rect 16040 2150 16092 2202
rect 20729 2150 20781 2202
rect 20793 2150 20845 2202
rect 20857 2150 20909 2202
rect 20921 2150 20973 2202
rect 20985 2150 21037 2202
<< metal2 >>
rect 3698 21298 3754 22000
rect 3698 21270 4016 21298
rect 3698 21200 3754 21270
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2424 18698 2452 19314
rect 3422 19068 3730 19077
rect 3422 19066 3428 19068
rect 3484 19066 3508 19068
rect 3564 19066 3588 19068
rect 3644 19066 3668 19068
rect 3724 19066 3730 19068
rect 3484 19014 3486 19066
rect 3666 19014 3668 19066
rect 3422 19012 3428 19014
rect 3484 19012 3508 19014
rect 3564 19012 3588 19014
rect 3644 19012 3668 19014
rect 3724 19012 3730 19014
rect 3422 19003 3730 19012
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2412 18692 2464 18698
rect 2412 18634 2464 18640
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1768 17672 1820 17678
rect 1952 17672 2004 17678
rect 1768 17614 1820 17620
rect 1872 17620 1952 17626
rect 1872 17614 2004 17620
rect 1780 12918 1808 17614
rect 1872 17598 1992 17614
rect 1872 17134 1900 17598
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17202 1992 17478
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1872 16574 1900 17070
rect 2056 16590 2084 18226
rect 2332 17882 2360 18634
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2148 17066 2176 17614
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2044 16584 2096 16590
rect 1872 16546 1992 16574
rect 1964 16114 1992 16546
rect 2424 16574 2452 18634
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 18290 3004 18566
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3068 17678 3096 18022
rect 3422 17980 3730 17989
rect 3422 17978 3428 17980
rect 3484 17978 3508 17980
rect 3564 17978 3588 17980
rect 3644 17978 3668 17980
rect 3724 17978 3730 17980
rect 3484 17926 3486 17978
rect 3666 17926 3668 17978
rect 3422 17924 3428 17926
rect 3484 17924 3508 17926
rect 3564 17924 3588 17926
rect 3644 17924 3668 17926
rect 3724 17924 3730 17926
rect 3422 17915 3730 17924
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2424 16546 2544 16574
rect 2044 16526 2096 16532
rect 2056 16130 2084 16526
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2240 16250 2268 16458
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2056 16114 2176 16130
rect 1952 16108 2004 16114
rect 2056 16108 2188 16114
rect 2056 16102 2136 16108
rect 1952 16050 2004 16056
rect 2136 16050 2188 16056
rect 1964 15314 1992 16050
rect 2044 15360 2096 15366
rect 1964 15308 2044 15314
rect 1964 15302 2096 15308
rect 1964 15286 2084 15302
rect 1964 14958 1992 15286
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1964 14482 1992 14894
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1872 12714 1900 13874
rect 1964 13870 1992 14418
rect 2148 14414 2176 16050
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2332 15026 2360 15574
rect 2424 15502 2452 15846
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2424 14958 2452 15438
rect 2516 15434 2544 16546
rect 2792 16250 2820 16662
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1964 12918 1992 13806
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1952 12912 2004 12918
rect 1952 12854 2004 12860
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 11762 1716 12106
rect 1872 11898 1900 12242
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1688 11150 1716 11698
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1872 10674 1900 11834
rect 1964 11626 1992 12174
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1964 10742 1992 11086
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1872 9926 1900 10610
rect 1964 10062 1992 10678
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 6798 1900 8774
rect 1964 7410 1992 9998
rect 2056 8498 2084 13262
rect 2148 12850 2176 13806
rect 2332 13326 2360 14282
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 14074 2452 14214
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2516 13954 2544 15370
rect 2424 13938 2544 13954
rect 3160 13938 3188 17478
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3422 16892 3730 16901
rect 3422 16890 3428 16892
rect 3484 16890 3508 16892
rect 3564 16890 3588 16892
rect 3644 16890 3668 16892
rect 3724 16890 3730 16892
rect 3484 16838 3486 16890
rect 3666 16838 3668 16890
rect 3422 16836 3428 16838
rect 3484 16836 3508 16838
rect 3564 16836 3588 16838
rect 3644 16836 3668 16838
rect 3724 16836 3730 16838
rect 3422 16827 3730 16836
rect 3896 16182 3924 16934
rect 3988 16794 4016 21270
rect 10704 21270 10916 21298
rect 5894 19612 6202 19621
rect 5894 19610 5900 19612
rect 5956 19610 5980 19612
rect 6036 19610 6060 19612
rect 6116 19610 6140 19612
rect 6196 19610 6202 19612
rect 5956 19558 5958 19610
rect 6138 19558 6140 19610
rect 5894 19556 5900 19558
rect 5956 19556 5980 19558
rect 6036 19556 6060 19558
rect 6116 19556 6140 19558
rect 6196 19556 6202 19558
rect 5894 19547 6202 19556
rect 10704 19446 10732 21270
rect 10888 21162 10916 21270
rect 10966 21200 11022 22000
rect 18234 21200 18290 22000
rect 10980 21162 11008 21200
rect 10888 21134 11008 21162
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 10839 19612 11147 19621
rect 10839 19610 10845 19612
rect 10901 19610 10925 19612
rect 10981 19610 11005 19612
rect 11061 19610 11085 19612
rect 11141 19610 11147 19612
rect 10901 19558 10903 19610
rect 11083 19558 11085 19610
rect 10839 19556 10845 19558
rect 10901 19556 10925 19558
rect 10981 19556 11005 19558
rect 11061 19556 11085 19558
rect 11141 19556 11147 19558
rect 10839 19547 11147 19556
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3422 15804 3730 15813
rect 3422 15802 3428 15804
rect 3484 15802 3508 15804
rect 3564 15802 3588 15804
rect 3644 15802 3668 15804
rect 3724 15802 3730 15804
rect 3484 15750 3486 15802
rect 3666 15750 3668 15802
rect 3422 15748 3428 15750
rect 3484 15748 3508 15750
rect 3564 15748 3588 15750
rect 3644 15748 3668 15750
rect 3724 15748 3730 15750
rect 3422 15739 3730 15748
rect 4172 15162 4200 18634
rect 4908 18358 4936 19110
rect 6840 18970 6868 19314
rect 8367 19068 8675 19077
rect 8367 19066 8373 19068
rect 8429 19066 8453 19068
rect 8509 19066 8533 19068
rect 8589 19066 8613 19068
rect 8669 19066 8675 19068
rect 8429 19014 8431 19066
rect 8611 19014 8613 19066
rect 8367 19012 8373 19014
rect 8429 19012 8453 19014
rect 8509 19012 8533 19014
rect 8589 19012 8613 19014
rect 8669 19012 8675 19014
rect 8367 19003 8675 19012
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 11256 18902 11284 19654
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 11716 18766 11744 19246
rect 13312 19068 13620 19077
rect 13312 19066 13318 19068
rect 13374 19066 13398 19068
rect 13454 19066 13478 19068
rect 13534 19066 13558 19068
rect 13614 19066 13620 19068
rect 13374 19014 13376 19066
rect 13556 19014 13558 19066
rect 13312 19012 13318 19014
rect 13374 19012 13398 19014
rect 13454 19012 13478 19014
rect 13534 19012 13558 19014
rect 13614 19012 13620 19014
rect 13312 19003 13620 19012
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 5368 18222 5396 18702
rect 5894 18524 6202 18533
rect 5894 18522 5900 18524
rect 5956 18522 5980 18524
rect 6036 18522 6060 18524
rect 6116 18522 6140 18524
rect 6196 18522 6202 18524
rect 5956 18470 5958 18522
rect 6138 18470 6140 18522
rect 5894 18468 5900 18470
rect 5956 18468 5980 18470
rect 6036 18468 6060 18470
rect 6116 18468 6140 18470
rect 6196 18468 6202 18470
rect 5894 18459 6202 18468
rect 7576 18290 7604 18702
rect 8208 18352 8260 18358
rect 8206 18320 8208 18329
rect 8260 18320 8262 18329
rect 7564 18284 7616 18290
rect 8206 18255 8262 18264
rect 7564 18226 7616 18232
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5368 17678 5396 18158
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5368 17202 5396 17614
rect 6196 17610 6224 18022
rect 7576 17678 7604 18226
rect 9232 18222 9260 18702
rect 10839 18524 11147 18533
rect 10839 18522 10845 18524
rect 10901 18522 10925 18524
rect 10981 18522 11005 18524
rect 11061 18522 11085 18524
rect 11141 18522 11147 18524
rect 10901 18470 10903 18522
rect 11083 18470 11085 18522
rect 10839 18468 10845 18470
rect 10901 18468 10925 18470
rect 10981 18468 11005 18470
rect 11061 18468 11085 18470
rect 11141 18468 11147 18470
rect 10839 18459 11147 18468
rect 11716 18222 11744 18702
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 8367 17980 8675 17989
rect 8367 17978 8373 17980
rect 8429 17978 8453 17980
rect 8509 17978 8533 17980
rect 8589 17978 8613 17980
rect 8669 17978 8675 17980
rect 8429 17926 8431 17978
rect 8611 17926 8613 17978
rect 8367 17924 8373 17926
rect 8429 17924 8453 17926
rect 8509 17924 8533 17926
rect 8589 17924 8613 17926
rect 8669 17924 8675 17926
rect 8367 17915 8675 17924
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 6184 17604 6236 17610
rect 6184 17546 6236 17552
rect 5894 17436 6202 17445
rect 5894 17434 5900 17436
rect 5956 17434 5980 17436
rect 6036 17434 6060 17436
rect 6116 17434 6140 17436
rect 6196 17434 6202 17436
rect 5956 17382 5958 17434
rect 6138 17382 6140 17434
rect 5894 17380 5900 17382
rect 5956 17380 5980 17382
rect 6036 17380 6060 17382
rect 6116 17380 6140 17382
rect 6196 17380 6202 17382
rect 5894 17371 6202 17380
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3422 14716 3730 14725
rect 3422 14714 3428 14716
rect 3484 14714 3508 14716
rect 3564 14714 3588 14716
rect 3644 14714 3668 14716
rect 3724 14714 3730 14716
rect 3484 14662 3486 14714
rect 3666 14662 3668 14714
rect 3422 14660 3428 14662
rect 3484 14660 3508 14662
rect 3564 14660 3588 14662
rect 3644 14660 3668 14662
rect 3724 14660 3730 14662
rect 3422 14651 3730 14660
rect 2412 13932 2544 13938
rect 2464 13926 2544 13932
rect 3148 13932 3200 13938
rect 2412 13874 2464 13880
rect 3148 13874 3200 13880
rect 3608 13932 3660 13938
rect 3976 13932 4028 13938
rect 3660 13892 3976 13920
rect 3608 13874 3660 13880
rect 3976 13874 4028 13880
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11354 2268 11630
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2240 8498 2268 9862
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2056 7954 2084 8434
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2240 7886 2268 8434
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2148 6798 2176 7142
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1964 6458 1992 6666
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2240 5710 2268 7346
rect 2332 7206 2360 13262
rect 2424 11762 2452 13874
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2884 13462 2912 13738
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2424 11150 2452 11698
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2424 10470 2452 11086
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2424 6186 2452 10406
rect 2516 7342 2544 12854
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2700 9994 2728 10474
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10062 2820 10406
rect 2884 10266 2912 10610
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2700 9110 2728 9930
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7410 2636 7686
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2516 5794 2544 7278
rect 2424 5766 2544 5794
rect 2424 5710 2452 5766
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2240 5302 2268 5646
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2424 5234 2452 5646
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2792 2446 2820 9318
rect 3160 8974 3188 13874
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3422 13628 3730 13637
rect 3422 13626 3428 13628
rect 3484 13626 3508 13628
rect 3564 13626 3588 13628
rect 3644 13626 3668 13628
rect 3724 13626 3730 13628
rect 3484 13574 3486 13626
rect 3666 13574 3668 13626
rect 3422 13572 3428 13574
rect 3484 13572 3508 13574
rect 3564 13572 3588 13574
rect 3644 13572 3668 13574
rect 3724 13572 3730 13574
rect 3422 13563 3730 13572
rect 3988 13394 4016 13738
rect 4264 13462 4292 17138
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 14414 5304 16390
rect 5460 16114 5488 16594
rect 7576 16522 7604 17614
rect 9232 17134 9260 18158
rect 10839 17436 11147 17445
rect 10839 17434 10845 17436
rect 10901 17434 10925 17436
rect 10981 17434 11005 17436
rect 11061 17434 11085 17436
rect 11141 17434 11147 17436
rect 10901 17382 10903 17434
rect 11083 17382 11085 17434
rect 10839 17380 10845 17382
rect 10901 17380 10925 17382
rect 10981 17380 11005 17382
rect 11061 17380 11085 17382
rect 11141 17380 11147 17382
rect 10839 17371 11147 17380
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 8367 16892 8675 16901
rect 8367 16890 8373 16892
rect 8429 16890 8453 16892
rect 8509 16890 8533 16892
rect 8589 16890 8613 16892
rect 8669 16890 8675 16892
rect 8429 16838 8431 16890
rect 8611 16838 8613 16890
rect 8367 16836 8373 16838
rect 8429 16836 8453 16838
rect 8509 16836 8533 16838
rect 8589 16836 8613 16838
rect 8669 16836 8675 16838
rect 8367 16827 8675 16836
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 5894 16348 6202 16357
rect 5894 16346 5900 16348
rect 5956 16346 5980 16348
rect 6036 16346 6060 16348
rect 6116 16346 6140 16348
rect 6196 16346 6202 16348
rect 5956 16294 5958 16346
rect 6138 16294 6140 16346
rect 5894 16292 5900 16294
rect 5956 16292 5980 16294
rect 6036 16292 6060 16294
rect 6116 16292 6140 16294
rect 6196 16292 6202 16294
rect 5894 16283 6202 16292
rect 7576 16114 7604 16458
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 6012 15706 6040 16050
rect 8312 15858 8340 16730
rect 9232 16658 9260 17070
rect 11164 16794 11192 17138
rect 11716 17134 11744 18158
rect 13312 17980 13620 17989
rect 13312 17978 13318 17980
rect 13374 17978 13398 17980
rect 13454 17978 13478 17980
rect 13534 17978 13558 17980
rect 13614 17978 13620 17980
rect 13374 17926 13376 17978
rect 13556 17926 13558 17978
rect 13312 17924 13318 17926
rect 13374 17924 13398 17926
rect 13454 17924 13478 17926
rect 13534 17924 13558 17926
rect 13614 17924 13620 17926
rect 13312 17915 13620 17924
rect 13648 17882 13676 18634
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13740 17678 13768 19450
rect 14384 19446 14412 19654
rect 15784 19612 16092 19621
rect 15784 19610 15790 19612
rect 15846 19610 15870 19612
rect 15926 19610 15950 19612
rect 16006 19610 16030 19612
rect 16086 19610 16092 19612
rect 15846 19558 15848 19610
rect 16028 19558 16030 19610
rect 15784 19556 15790 19558
rect 15846 19556 15870 19558
rect 15926 19556 15950 19558
rect 16006 19556 16030 19558
rect 16086 19556 16092 19558
rect 15784 19547 16092 19556
rect 18248 19446 18276 21200
rect 20729 19612 21037 19621
rect 20729 19610 20735 19612
rect 20791 19610 20815 19612
rect 20871 19610 20895 19612
rect 20951 19610 20975 19612
rect 21031 19610 21037 19612
rect 20791 19558 20793 19610
rect 20973 19558 20975 19610
rect 20729 19556 20735 19558
rect 20791 19556 20815 19558
rect 20871 19556 20895 19558
rect 20951 19556 20975 19558
rect 21031 19556 21037 19558
rect 20729 19547 21037 19556
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14108 18902 14136 19178
rect 14200 18902 14228 19382
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14568 18766 14596 19314
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 14752 18970 14780 19110
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18154 13952 18566
rect 14752 18426 14780 18634
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 15028 18290 15056 18906
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15212 18329 15240 18566
rect 15198 18320 15254 18329
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 15016 18284 15068 18290
rect 15198 18255 15254 18264
rect 15016 18226 15068 18232
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 10506 16688 10562 16697
rect 9220 16652 9272 16658
rect 10506 16623 10562 16632
rect 9220 16594 9272 16600
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8220 15830 8340 15858
rect 8220 15722 8248 15830
rect 8367 15804 8675 15813
rect 8367 15802 8373 15804
rect 8429 15802 8453 15804
rect 8509 15802 8533 15804
rect 8589 15802 8613 15804
rect 8669 15802 8675 15804
rect 8429 15750 8431 15802
rect 8611 15750 8613 15802
rect 8367 15748 8373 15750
rect 8429 15748 8453 15750
rect 8509 15748 8533 15750
rect 8589 15748 8613 15750
rect 8669 15748 8675 15750
rect 8367 15739 8675 15748
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 6000 15700 6052 15706
rect 8220 15694 8340 15722
rect 6000 15642 6052 15648
rect 5644 14482 5672 15642
rect 5894 15260 6202 15269
rect 5894 15258 5900 15260
rect 5956 15258 5980 15260
rect 6036 15258 6060 15260
rect 6116 15258 6140 15260
rect 6196 15258 6202 15260
rect 5956 15206 5958 15258
rect 6138 15206 6140 15258
rect 5894 15204 5900 15206
rect 5956 15204 5980 15206
rect 6036 15204 6060 15206
rect 6116 15204 6140 15206
rect 6196 15204 6202 15206
rect 5894 15195 6202 15204
rect 8312 15094 8340 15694
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8367 14716 8675 14725
rect 8367 14714 8373 14716
rect 8429 14714 8453 14716
rect 8509 14714 8533 14716
rect 8589 14714 8613 14716
rect 8669 14714 8675 14716
rect 8429 14662 8431 14714
rect 8611 14662 8613 14714
rect 8367 14660 8373 14662
rect 8429 14660 8453 14662
rect 8509 14660 8533 14662
rect 8589 14660 8613 14662
rect 8669 14660 8675 14662
rect 8367 14651 8675 14660
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 5368 13530 5396 14350
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 5894 14172 6202 14181
rect 5894 14170 5900 14172
rect 5956 14170 5980 14172
rect 6036 14170 6060 14172
rect 6116 14170 6140 14172
rect 6196 14170 6202 14172
rect 5956 14118 5958 14170
rect 6138 14118 6140 14170
rect 5894 14116 5900 14118
rect 5956 14116 5980 14118
rect 6036 14116 6060 14118
rect 6116 14116 6140 14118
rect 6196 14116 6202 14118
rect 5894 14107 6202 14116
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 5552 13326 5580 13806
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12918 5580 13262
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 5894 13084 6202 13093
rect 5894 13082 5900 13084
rect 5956 13082 5980 13084
rect 6036 13082 6060 13084
rect 6116 13082 6140 13084
rect 6196 13082 6202 13084
rect 5956 13030 5958 13082
rect 6138 13030 6140 13082
rect 5894 13028 5900 13030
rect 5956 13028 5980 13030
rect 6036 13028 6060 13030
rect 6116 13028 6140 13030
rect 6196 13028 6202 13030
rect 5894 13019 6202 13028
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 3422 12540 3730 12549
rect 3422 12538 3428 12540
rect 3484 12538 3508 12540
rect 3564 12538 3588 12540
rect 3644 12538 3668 12540
rect 3724 12538 3730 12540
rect 3484 12486 3486 12538
rect 3666 12486 3668 12538
rect 3422 12484 3428 12486
rect 3484 12484 3508 12486
rect 3564 12484 3588 12486
rect 3644 12484 3668 12486
rect 3724 12484 3730 12486
rect 3422 12475 3730 12484
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 3422 11452 3730 11461
rect 3422 11450 3428 11452
rect 3484 11450 3508 11452
rect 3564 11450 3588 11452
rect 3644 11450 3668 11452
rect 3724 11450 3730 11452
rect 3484 11398 3486 11450
rect 3666 11398 3668 11450
rect 3422 11396 3428 11398
rect 3484 11396 3508 11398
rect 3564 11396 3588 11398
rect 3644 11396 3668 11398
rect 3724 11396 3730 11398
rect 3422 11387 3730 11396
rect 3422 10364 3730 10373
rect 3422 10362 3428 10364
rect 3484 10362 3508 10364
rect 3564 10362 3588 10364
rect 3644 10362 3668 10364
rect 3724 10362 3730 10364
rect 3484 10310 3486 10362
rect 3666 10310 3668 10362
rect 3422 10308 3428 10310
rect 3484 10308 3508 10310
rect 3564 10308 3588 10310
rect 3644 10308 3668 10310
rect 3724 10308 3730 10310
rect 3422 10299 3730 10308
rect 3422 9276 3730 9285
rect 3422 9274 3428 9276
rect 3484 9274 3508 9276
rect 3564 9274 3588 9276
rect 3644 9274 3668 9276
rect 3724 9274 3730 9276
rect 3484 9222 3486 9274
rect 3666 9222 3668 9274
rect 3422 9220 3428 9222
rect 3484 9220 3508 9222
rect 3564 9220 3588 9222
rect 3644 9220 3668 9222
rect 3724 9220 3730 9222
rect 3422 9211 3730 9220
rect 4264 9178 4292 12038
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4448 8974 4476 12786
rect 5552 12238 5580 12854
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11762 5580 12174
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5552 11150 5580 11698
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10674 5580 11086
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 10266 5580 10610
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3160 7274 3188 8502
rect 4080 8430 4108 8910
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8430 4384 8774
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 3422 8188 3730 8197
rect 3422 8186 3428 8188
rect 3484 8186 3508 8188
rect 3564 8186 3588 8188
rect 3644 8186 3668 8188
rect 3724 8186 3730 8188
rect 3484 8134 3486 8186
rect 3666 8134 3668 8186
rect 3422 8132 3428 8134
rect 3484 8132 3508 8134
rect 3564 8132 3588 8134
rect 3644 8132 3668 8134
rect 3724 8132 3730 8134
rect 3422 8123 3730 8132
rect 4080 7546 4108 8366
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4356 7342 4384 8366
rect 4448 8022 4476 8910
rect 4632 8634 4660 9522
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4540 7886 4568 8366
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4540 7546 4568 7822
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4896 7336 4948 7342
rect 4948 7284 5120 7290
rect 4896 7278 5120 7284
rect 4908 7274 5120 7278
rect 3148 7268 3200 7274
rect 4908 7268 5132 7274
rect 4908 7262 5080 7268
rect 3148 7210 3200 7216
rect 5080 7210 5132 7216
rect 3160 6322 3188 7210
rect 3422 7100 3730 7109
rect 3422 7098 3428 7100
rect 3484 7098 3508 7100
rect 3564 7098 3588 7100
rect 3644 7098 3668 7100
rect 3724 7098 3730 7100
rect 3484 7046 3486 7098
rect 3666 7046 3668 7098
rect 3422 7044 3428 7046
rect 3484 7044 3508 7046
rect 3564 7044 3588 7046
rect 3644 7044 3668 7046
rect 3724 7044 3730 7046
rect 3422 7035 3730 7044
rect 5184 7002 5212 7822
rect 5460 7818 5488 8366
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5368 7478 5396 7754
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5368 6866 5396 7414
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5234 2912 5646
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3160 4622 3188 6258
rect 3712 6254 3740 6598
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3422 6012 3730 6021
rect 3422 6010 3428 6012
rect 3484 6010 3508 6012
rect 3564 6010 3588 6012
rect 3644 6010 3668 6012
rect 3724 6010 3730 6012
rect 3484 5958 3486 6010
rect 3666 5958 3668 6010
rect 3422 5956 3428 5958
rect 3484 5956 3508 5958
rect 3564 5956 3588 5958
rect 3644 5956 3668 5958
rect 3724 5956 3730 5958
rect 3422 5947 3730 5956
rect 3988 5914 4016 6258
rect 5184 6118 5212 6326
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4264 5778 4292 6054
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5098 3372 5646
rect 5184 5574 5212 6054
rect 5368 5846 5396 6802
rect 5460 6798 5488 7754
rect 5552 7546 5580 8434
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6866 5580 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3344 4690 3372 5034
rect 3422 4924 3730 4933
rect 3422 4922 3428 4924
rect 3484 4922 3508 4924
rect 3564 4922 3588 4924
rect 3644 4922 3668 4924
rect 3724 4922 3730 4924
rect 3484 4870 3486 4922
rect 3666 4870 3668 4922
rect 3422 4868 3428 4870
rect 3484 4868 3508 4870
rect 3564 4868 3588 4870
rect 3644 4868 3668 4870
rect 3724 4868 3730 4870
rect 3422 4859 3730 4868
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3422 3836 3730 3845
rect 3422 3834 3428 3836
rect 3484 3834 3508 3836
rect 3564 3834 3588 3836
rect 3644 3834 3668 3836
rect 3724 3834 3730 3836
rect 3484 3782 3486 3834
rect 3666 3782 3668 3834
rect 3422 3780 3428 3782
rect 3484 3780 3508 3782
rect 3564 3780 3588 3782
rect 3644 3780 3668 3782
rect 3724 3780 3730 3782
rect 3422 3771 3730 3780
rect 5644 2774 5672 12582
rect 5894 11996 6202 12005
rect 5894 11994 5900 11996
rect 5956 11994 5980 11996
rect 6036 11994 6060 11996
rect 6116 11994 6140 11996
rect 6196 11994 6202 11996
rect 5956 11942 5958 11994
rect 6138 11942 6140 11994
rect 5894 11940 5900 11942
rect 5956 11940 5980 11942
rect 6036 11940 6060 11942
rect 6116 11940 6140 11942
rect 6196 11940 6202 11942
rect 5894 11931 6202 11940
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 8974 5764 9522
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5828 8634 5856 11018
rect 5894 10908 6202 10917
rect 5894 10906 5900 10908
rect 5956 10906 5980 10908
rect 6036 10906 6060 10908
rect 6116 10906 6140 10908
rect 6196 10906 6202 10908
rect 5956 10854 5958 10906
rect 6138 10854 6140 10906
rect 5894 10852 5900 10854
rect 5956 10852 5980 10854
rect 6036 10852 6060 10854
rect 6116 10852 6140 10854
rect 6196 10852 6202 10854
rect 5894 10843 6202 10852
rect 5894 9820 6202 9829
rect 5894 9818 5900 9820
rect 5956 9818 5980 9820
rect 6036 9818 6060 9820
rect 6116 9818 6140 9820
rect 6196 9818 6202 9820
rect 5956 9766 5958 9818
rect 6138 9766 6140 9818
rect 5894 9764 5900 9766
rect 5956 9764 5980 9766
rect 6036 9764 6060 9766
rect 6116 9764 6140 9766
rect 6196 9764 6202 9766
rect 5894 9755 6202 9764
rect 5894 8732 6202 8741
rect 5894 8730 5900 8732
rect 5956 8730 5980 8732
rect 6036 8730 6060 8732
rect 6116 8730 6140 8732
rect 6196 8730 6202 8732
rect 5956 8678 5958 8730
rect 6138 8678 6140 8730
rect 5894 8676 5900 8678
rect 5956 8676 5980 8678
rect 6036 8676 6060 8678
rect 6116 8676 6140 8678
rect 6196 8676 6202 8678
rect 5894 8667 6202 8676
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5736 7886 5764 8434
rect 5828 7886 5856 8570
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7886 6224 8366
rect 6472 8090 6500 13194
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6564 11762 6592 12174
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6564 10674 6592 11698
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 9586 6592 10610
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 6184 7880 6236 7886
rect 6236 7840 6316 7868
rect 6184 7822 6236 7828
rect 5894 7644 6202 7653
rect 5894 7642 5900 7644
rect 5956 7642 5980 7644
rect 6036 7642 6060 7644
rect 6116 7642 6140 7644
rect 6196 7642 6202 7644
rect 5956 7590 5958 7642
rect 6138 7590 6140 7642
rect 5894 7588 5900 7590
rect 5956 7588 5980 7590
rect 6036 7588 6060 7590
rect 6116 7588 6140 7590
rect 6196 7588 6202 7590
rect 5894 7579 6202 7588
rect 6288 7410 6316 7840
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5920 6866 5948 7346
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5894 6556 6202 6565
rect 5894 6554 5900 6556
rect 5956 6554 5980 6556
rect 6036 6554 6060 6556
rect 6116 6554 6140 6556
rect 6196 6554 6202 6556
rect 5956 6502 5958 6554
rect 6138 6502 6140 6554
rect 5894 6500 5900 6502
rect 5956 6500 5980 6502
rect 6036 6500 6060 6502
rect 6116 6500 6140 6502
rect 6196 6500 6202 6502
rect 5894 6491 6202 6500
rect 6288 6390 6316 7346
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6472 6458 6500 6870
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5828 5216 5856 6258
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 5894 5468 6202 5477
rect 5894 5466 5900 5468
rect 5956 5466 5980 5468
rect 6036 5466 6060 5468
rect 6116 5466 6140 5468
rect 6196 5466 6202 5468
rect 5956 5414 5958 5466
rect 6138 5414 6140 5466
rect 5894 5412 5900 5414
rect 5956 5412 5980 5414
rect 6036 5412 6060 5414
rect 6116 5412 6140 5414
rect 6196 5412 6202 5414
rect 5894 5403 6202 5412
rect 6288 5370 6316 5646
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6656 5302 6684 11222
rect 6840 8634 6868 11698
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6748 7750 6776 8434
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5574 6868 6258
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6000 5228 6052 5234
rect 5828 5188 6000 5216
rect 6000 5170 6052 5176
rect 6012 4690 6040 5170
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6288 4622 6316 4694
rect 6656 4622 6684 5102
rect 7116 4758 7144 6190
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7300 5370 7328 5578
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7392 4690 7420 5646
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 5894 4380 6202 4389
rect 5894 4378 5900 4380
rect 5956 4378 5980 4380
rect 6036 4378 6060 4380
rect 6116 4378 6140 4380
rect 6196 4378 6202 4380
rect 5956 4326 5958 4378
rect 6138 4326 6140 4378
rect 5894 4324 5900 4326
rect 5956 4324 5980 4326
rect 6036 4324 6060 4326
rect 6116 4324 6140 4326
rect 6196 4324 6202 4326
rect 5894 4315 6202 4324
rect 5894 3292 6202 3301
rect 5894 3290 5900 3292
rect 5956 3290 5980 3292
rect 6036 3290 6060 3292
rect 6116 3290 6140 3292
rect 6196 3290 6202 3292
rect 5956 3238 5958 3290
rect 6138 3238 6140 3290
rect 5894 3236 5900 3238
rect 5956 3236 5980 3238
rect 6036 3236 6060 3238
rect 6116 3236 6140 3238
rect 6196 3236 6202 3238
rect 5894 3227 6202 3236
rect 3422 2748 3730 2757
rect 3422 2746 3428 2748
rect 3484 2746 3508 2748
rect 3564 2746 3588 2748
rect 3644 2746 3668 2748
rect 3724 2746 3730 2748
rect 3484 2694 3486 2746
rect 3666 2694 3668 2746
rect 3422 2692 3428 2694
rect 3484 2692 3508 2694
rect 3564 2692 3588 2694
rect 3644 2692 3668 2694
rect 3724 2692 3730 2694
rect 3422 2683 3730 2692
rect 5552 2746 5672 2774
rect 5552 2446 5580 2746
rect 7484 2446 7512 13126
rect 7576 8634 7604 14282
rect 7944 13938 7972 14350
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7944 12850 7972 13874
rect 8367 13628 8675 13637
rect 8367 13626 8373 13628
rect 8429 13626 8453 13628
rect 8509 13626 8533 13628
rect 8589 13626 8613 13628
rect 8669 13626 8675 13628
rect 8429 13574 8431 13626
rect 8611 13574 8613 13626
rect 8367 13572 8373 13574
rect 8429 13572 8453 13574
rect 8509 13572 8533 13574
rect 8589 13572 8613 13574
rect 8669 13572 8675 13574
rect 8367 13563 8675 13572
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12238 7972 12786
rect 8367 12540 8675 12549
rect 8367 12538 8373 12540
rect 8429 12538 8453 12540
rect 8509 12538 8533 12540
rect 8589 12538 8613 12540
rect 8669 12538 8675 12540
rect 8429 12486 8431 12538
rect 8611 12486 8613 12538
rect 8367 12484 8373 12486
rect 8429 12484 8453 12486
rect 8509 12484 8533 12486
rect 8589 12484 8613 12486
rect 8669 12484 8675 12486
rect 8367 12475 8675 12484
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7760 9178 7788 9998
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 7954 7696 8434
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7478 7696 7890
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7576 6186 7604 6666
rect 7668 6390 7696 6734
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7760 6322 7788 6598
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 5234 7604 6122
rect 7564 5228 7616 5234
rect 7616 5188 7696 5216
rect 7564 5170 7616 5176
rect 7668 4622 7696 5188
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7852 2774 7880 11494
rect 8367 11452 8675 11461
rect 8367 11450 8373 11452
rect 8429 11450 8453 11452
rect 8509 11450 8533 11452
rect 8589 11450 8613 11452
rect 8669 11450 8675 11452
rect 8429 11398 8431 11450
rect 8611 11398 8613 11450
rect 8367 11396 8373 11398
rect 8429 11396 8453 11398
rect 8509 11396 8533 11398
rect 8589 11396 8613 11398
rect 8669 11396 8675 11398
rect 8367 11387 8675 11396
rect 8367 10364 8675 10373
rect 8367 10362 8373 10364
rect 8429 10362 8453 10364
rect 8509 10362 8533 10364
rect 8589 10362 8613 10364
rect 8669 10362 8675 10364
rect 8429 10310 8431 10362
rect 8611 10310 8613 10362
rect 8367 10308 8373 10310
rect 8429 10308 8453 10310
rect 8509 10308 8533 10310
rect 8589 10308 8613 10310
rect 8669 10308 8675 10310
rect 8367 10299 8675 10308
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7944 6798 7972 9862
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 8090 8064 9522
rect 8367 9276 8675 9285
rect 8367 9274 8373 9276
rect 8429 9274 8453 9276
rect 8509 9274 8533 9276
rect 8589 9274 8613 9276
rect 8669 9274 8675 9276
rect 8429 9222 8431 9274
rect 8611 9222 8613 9274
rect 8367 9220 8373 9222
rect 8429 9220 8453 9222
rect 8509 9220 8533 9222
rect 8589 9220 8613 9222
rect 8669 9220 8675 9222
rect 8367 9211 8675 9220
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8128 8498 8156 8842
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8128 7886 8156 8434
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8036 6254 8064 6666
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5166 8064 6190
rect 8128 5846 8156 7822
rect 8220 6322 8248 8366
rect 8367 8188 8675 8197
rect 8367 8186 8373 8188
rect 8429 8186 8453 8188
rect 8509 8186 8533 8188
rect 8589 8186 8613 8188
rect 8669 8186 8675 8188
rect 8429 8134 8431 8186
rect 8611 8134 8613 8186
rect 8367 8132 8373 8134
rect 8429 8132 8453 8134
rect 8509 8132 8533 8134
rect 8589 8132 8613 8134
rect 8669 8132 8675 8134
rect 8367 8123 8675 8132
rect 8367 7100 8675 7109
rect 8367 7098 8373 7100
rect 8429 7098 8453 7100
rect 8509 7098 8533 7100
rect 8589 7098 8613 7100
rect 8669 7098 8675 7100
rect 8429 7046 8431 7098
rect 8611 7046 8613 7098
rect 8367 7044 8373 7046
rect 8429 7044 8453 7046
rect 8509 7044 8533 7046
rect 8589 7044 8613 7046
rect 8669 7044 8675 7046
rect 8367 7035 8675 7044
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8220 5692 8248 6054
rect 8367 6012 8675 6021
rect 8367 6010 8373 6012
rect 8429 6010 8453 6012
rect 8509 6010 8533 6012
rect 8589 6010 8613 6012
rect 8669 6010 8675 6012
rect 8429 5958 8431 6010
rect 8611 5958 8613 6010
rect 8367 5956 8373 5958
rect 8429 5956 8453 5958
rect 8509 5956 8533 5958
rect 8589 5956 8613 5958
rect 8669 5956 8675 5958
rect 8367 5947 8675 5956
rect 8300 5704 8352 5710
rect 8220 5664 8300 5692
rect 8300 5646 8352 5652
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7944 4622 7972 5034
rect 8367 4924 8675 4933
rect 8367 4922 8373 4924
rect 8429 4922 8453 4924
rect 8509 4922 8533 4924
rect 8589 4922 8613 4924
rect 8669 4922 8675 4924
rect 8429 4870 8431 4922
rect 8611 4870 8613 4922
rect 8367 4868 8373 4870
rect 8429 4868 8453 4870
rect 8509 4868 8533 4870
rect 8589 4868 8613 4870
rect 8669 4868 8675 4870
rect 8367 4859 8675 4868
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8367 3836 8675 3845
rect 8367 3834 8373 3836
rect 8429 3834 8453 3836
rect 8509 3834 8533 3836
rect 8589 3834 8613 3836
rect 8669 3834 8675 3836
rect 8429 3782 8431 3834
rect 8611 3782 8613 3834
rect 8367 3780 8373 3782
rect 8429 3780 8453 3782
rect 8509 3780 8533 3782
rect 8589 3780 8613 3782
rect 8669 3780 8675 3782
rect 8367 3771 8675 3780
rect 7852 2746 7972 2774
rect 7944 2582 7972 2746
rect 8367 2748 8675 2757
rect 8367 2746 8373 2748
rect 8429 2746 8453 2748
rect 8509 2746 8533 2748
rect 8589 2746 8613 2748
rect 8669 2746 8675 2748
rect 8429 2694 8431 2746
rect 8611 2694 8613 2746
rect 8367 2692 8373 2694
rect 8429 2692 8453 2694
rect 8509 2692 8533 2694
rect 8589 2692 8613 2694
rect 8669 2692 8675 2694
rect 8367 2683 8675 2692
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 8772 2514 8800 14214
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8864 8566 8892 12718
rect 9140 12434 9168 16050
rect 9232 15026 9260 16594
rect 10520 16590 10548 16623
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 14482 9260 14962
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9324 12434 9352 16458
rect 10612 16250 10640 16730
rect 11716 16658 11744 17070
rect 13312 16892 13620 16901
rect 13312 16890 13318 16892
rect 13374 16890 13398 16892
rect 13454 16890 13478 16892
rect 13534 16890 13558 16892
rect 13614 16890 13620 16892
rect 13374 16838 13376 16890
rect 13556 16838 13558 16890
rect 13312 16836 13318 16838
rect 13374 16836 13398 16838
rect 13454 16836 13478 16838
rect 13534 16836 13558 16838
rect 13614 16836 13620 16838
rect 13312 16827 13620 16836
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 10839 16348 11147 16357
rect 10839 16346 10845 16348
rect 10901 16346 10925 16348
rect 10981 16346 11005 16348
rect 11061 16346 11085 16348
rect 11141 16346 11147 16348
rect 10901 16294 10903 16346
rect 11083 16294 11085 16346
rect 10839 16292 10845 16294
rect 10901 16292 10925 16294
rect 10981 16292 11005 16294
rect 11061 16292 11085 16294
rect 11141 16292 11147 16294
rect 10839 16283 11147 16292
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 11716 16114 11744 16594
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9140 12406 9260 12434
rect 9324 12406 9444 12434
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8090 9076 8230
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6458 8984 6666
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8864 5710 8892 6326
rect 9140 6322 9168 8774
rect 9232 6458 9260 12406
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9324 7886 9352 8434
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9416 7342 9444 12406
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9508 6390 9536 15846
rect 11716 15706 11744 16050
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9600 15162 9628 15370
rect 10839 15260 11147 15269
rect 10839 15258 10845 15260
rect 10901 15258 10925 15260
rect 10981 15258 11005 15260
rect 11061 15258 11085 15260
rect 11141 15258 11147 15260
rect 10901 15206 10903 15258
rect 11083 15206 11085 15258
rect 10839 15204 10845 15206
rect 10901 15204 10925 15206
rect 10981 15204 11005 15206
rect 11061 15204 11085 15206
rect 11141 15204 11147 15206
rect 10839 15195 11147 15204
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9600 9994 9628 15098
rect 11716 15026 11744 15642
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 7886 9628 8298
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9508 6118 9536 6326
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5166 9444 5646
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 9692 2446 9720 12038
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9784 9042 9812 9522
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9876 8566 9904 14350
rect 10839 14172 11147 14181
rect 10839 14170 10845 14172
rect 10901 14170 10925 14172
rect 10981 14170 11005 14172
rect 11061 14170 11085 14172
rect 11141 14170 11147 14172
rect 10901 14118 10903 14170
rect 11083 14118 11085 14170
rect 10839 14116 10845 14118
rect 10901 14116 10925 14118
rect 10981 14116 11005 14118
rect 11061 14116 11085 14118
rect 11141 14116 11147 14118
rect 10839 14107 11147 14116
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 6322 9812 7686
rect 9968 6662 9996 10542
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7274 10088 8230
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 5710 9996 6190
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10060 5710 10088 6122
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10152 4826 10180 13874
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 10839 13084 11147 13093
rect 10839 13082 10845 13084
rect 10901 13082 10925 13084
rect 10981 13082 11005 13084
rect 11061 13082 11085 13084
rect 11141 13082 11147 13084
rect 10901 13030 10903 13082
rect 11083 13030 11085 13082
rect 10839 13028 10845 13030
rect 10901 13028 10925 13030
rect 10981 13028 11005 13030
rect 11061 13028 11085 13030
rect 11141 13028 11147 13030
rect 10839 13019 11147 13028
rect 11716 12850 11744 13806
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7478 10272 7686
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10336 7410 10364 8502
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10428 7546 10456 8434
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10428 6798 10456 7482
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10230 6352 10286 6361
rect 10230 6287 10232 6296
rect 10284 6287 10286 6296
rect 10232 6258 10284 6264
rect 10428 5710 10456 6734
rect 10612 5914 10640 12106
rect 10839 11996 11147 12005
rect 10839 11994 10845 11996
rect 10901 11994 10925 11996
rect 10981 11994 11005 11996
rect 11061 11994 11085 11996
rect 11141 11994 11147 11996
rect 10901 11942 10903 11994
rect 11083 11942 11085 11994
rect 10839 11940 10845 11942
rect 10901 11940 10925 11942
rect 10981 11940 11005 11942
rect 11061 11940 11085 11942
rect 11141 11940 11147 11942
rect 10839 11931 11147 11940
rect 10839 10908 11147 10917
rect 10839 10906 10845 10908
rect 10901 10906 10925 10908
rect 10981 10906 11005 10908
rect 11061 10906 11085 10908
rect 11141 10906 11147 10908
rect 10901 10854 10903 10906
rect 11083 10854 11085 10906
rect 10839 10852 10845 10854
rect 10901 10852 10925 10854
rect 10981 10852 11005 10854
rect 11061 10852 11085 10854
rect 11141 10852 11147 10854
rect 10839 10843 11147 10852
rect 10839 9820 11147 9829
rect 10839 9818 10845 9820
rect 10901 9818 10925 9820
rect 10981 9818 11005 9820
rect 11061 9818 11085 9820
rect 11141 9818 11147 9820
rect 10901 9766 10903 9818
rect 11083 9766 11085 9818
rect 10839 9764 10845 9766
rect 10901 9764 10925 9766
rect 10981 9764 11005 9766
rect 11061 9764 11085 9766
rect 11141 9764 11147 9766
rect 10839 9755 11147 9764
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8634 10732 8842
rect 10839 8732 11147 8741
rect 10839 8730 10845 8732
rect 10901 8730 10925 8732
rect 10981 8730 11005 8732
rect 11061 8730 11085 8732
rect 11141 8730 11147 8732
rect 10901 8678 10903 8730
rect 11083 8678 11085 8730
rect 10839 8676 10845 8678
rect 10901 8676 10925 8678
rect 10981 8676 11005 8678
rect 11061 8676 11085 8678
rect 11141 8676 11147 8678
rect 10839 8667 11147 8676
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10888 8498 10916 8570
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11164 8090 11192 8434
rect 11256 8362 11284 12582
rect 11716 12238 11744 12786
rect 11900 12442 11928 16186
rect 13312 15804 13620 15813
rect 13312 15802 13318 15804
rect 13374 15802 13398 15804
rect 13454 15802 13478 15804
rect 13534 15802 13558 15804
rect 13614 15802 13620 15804
rect 13374 15750 13376 15802
rect 13556 15750 13558 15802
rect 13312 15748 13318 15750
rect 13374 15748 13398 15750
rect 13454 15748 13478 15750
rect 13534 15748 13558 15750
rect 13614 15748 13620 15750
rect 13312 15739 13620 15748
rect 13648 15434 13676 16662
rect 13740 15978 13768 17138
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13312 14716 13620 14725
rect 13312 14714 13318 14716
rect 13374 14714 13398 14716
rect 13454 14714 13478 14716
rect 13534 14714 13558 14716
rect 13614 14714 13620 14716
rect 13374 14662 13376 14714
rect 13556 14662 13558 14714
rect 13312 14660 13318 14662
rect 13374 14660 13398 14662
rect 13454 14660 13478 14662
rect 13534 14660 13558 14662
rect 13614 14660 13620 14662
rect 13312 14651 13620 14660
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 13870 12204 14350
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 13312 13628 13620 13637
rect 13312 13626 13318 13628
rect 13374 13626 13398 13628
rect 13454 13626 13478 13628
rect 13534 13626 13558 13628
rect 13614 13626 13620 13628
rect 13374 13574 13376 13626
rect 13556 13574 13558 13626
rect 13312 13572 13318 13574
rect 13374 13572 13398 13574
rect 13454 13572 13478 13574
rect 13534 13572 13558 13574
rect 13614 13572 13620 13574
rect 13312 13563 13620 13572
rect 13312 12540 13620 12549
rect 13312 12538 13318 12540
rect 13374 12538 13398 12540
rect 13454 12538 13478 12540
rect 13534 12538 13558 12540
rect 13614 12538 13620 12540
rect 13374 12486 13376 12538
rect 13556 12486 13558 12538
rect 13312 12484 13318 12486
rect 13374 12484 13398 12486
rect 13454 12484 13478 12486
rect 13534 12484 13558 12486
rect 13614 12484 13620 12486
rect 13312 12475 13620 12484
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11218 11652 12038
rect 11716 11762 11744 12174
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 12268 10674 12296 11698
rect 13312 11452 13620 11461
rect 13312 11450 13318 11452
rect 13374 11450 13398 11452
rect 13454 11450 13478 11452
rect 13534 11450 13558 11452
rect 13614 11450 13620 11452
rect 13374 11398 13376 11450
rect 13556 11398 13558 11450
rect 13312 11396 13318 11398
rect 13374 11396 13398 11398
rect 13454 11396 13478 11398
rect 13534 11396 13558 11398
rect 13614 11396 13620 11398
rect 13312 11387 13620 11396
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 8906 11652 10406
rect 12268 10130 12296 10610
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12268 9586 12296 10066
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11256 7818 11284 8298
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 10839 7644 11147 7653
rect 10839 7642 10845 7644
rect 10901 7642 10925 7644
rect 10981 7642 11005 7644
rect 11061 7642 11085 7644
rect 11141 7642 11147 7644
rect 10901 7590 10903 7642
rect 11083 7590 11085 7642
rect 10839 7588 10845 7590
rect 10901 7588 10925 7590
rect 10981 7588 11005 7590
rect 11061 7588 11085 7590
rect 11141 7588 11147 7590
rect 10839 7579 11147 7588
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6254 10732 6598
rect 10839 6556 11147 6565
rect 10839 6554 10845 6556
rect 10901 6554 10925 6556
rect 10981 6554 11005 6556
rect 11061 6554 11085 6556
rect 11141 6554 11147 6556
rect 10901 6502 10903 6554
rect 11083 6502 11085 6554
rect 10839 6500 10845 6502
rect 10901 6500 10925 6502
rect 10981 6500 11005 6502
rect 11061 6500 11085 6502
rect 11141 6500 11147 6502
rect 10839 6491 11147 6500
rect 11256 6322 11284 6666
rect 11348 6458 11376 8366
rect 11624 7206 11652 8842
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11716 7886 11744 8502
rect 11900 8430 11928 9318
rect 11888 8424 11940 8430
rect 11808 8372 11888 8378
rect 11808 8366 11940 8372
rect 11808 8350 11928 8366
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10704 5794 10732 6190
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5846 10824 6054
rect 10612 5766 10732 5794
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10612 4622 10640 5766
rect 10839 5468 11147 5477
rect 10839 5466 10845 5468
rect 10901 5466 10925 5468
rect 10981 5466 11005 5468
rect 11061 5466 11085 5468
rect 11141 5466 11147 5468
rect 10901 5414 10903 5466
rect 11083 5414 11085 5466
rect 10839 5412 10845 5414
rect 10901 5412 10925 5414
rect 10981 5412 11005 5414
rect 11061 5412 11085 5414
rect 11141 5412 11147 5414
rect 10839 5403 11147 5412
rect 11256 5234 11284 6258
rect 11348 6118 11376 6394
rect 11624 6322 11652 7142
rect 11716 6934 11744 7822
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11808 6798 11836 8350
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11900 7818 11928 8230
rect 11992 8022 12020 9522
rect 12268 8974 12296 9522
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12084 8362 12112 8502
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 12084 7274 12112 8298
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 7478 12296 7686
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12268 6934 12296 7414
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12452 6798 12480 8434
rect 12544 7478 12572 11154
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13312 10364 13620 10373
rect 13312 10362 13318 10364
rect 13374 10362 13398 10364
rect 13454 10362 13478 10364
rect 13534 10362 13558 10364
rect 13614 10362 13620 10364
rect 13374 10310 13376 10362
rect 13556 10310 13558 10362
rect 13312 10308 13318 10310
rect 13374 10308 13398 10310
rect 13454 10308 13478 10310
rect 13534 10308 13558 10310
rect 13614 10308 13620 10310
rect 13312 10299 13620 10308
rect 13740 9654 13768 10474
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 8090 12756 8230
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 11796 6792 11848 6798
rect 12440 6792 12492 6798
rect 11796 6734 11848 6740
rect 11992 6718 12204 6746
rect 12440 6734 12492 6740
rect 11992 6662 12020 6718
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12084 6474 12112 6598
rect 11992 6458 12112 6474
rect 11980 6452 12112 6458
rect 12032 6446 12112 6452
rect 11980 6394 12032 6400
rect 12176 6338 12204 6718
rect 12544 6662 12572 7414
rect 12728 6866 12756 7822
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11980 6316 12032 6322
rect 12176 6310 12296 6338
rect 11980 6258 12032 6264
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11808 6066 11836 6258
rect 11348 5642 11376 6054
rect 11808 6038 11928 6066
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10612 4078 10640 4558
rect 11256 4554 11284 5170
rect 11900 4622 11928 6038
rect 11992 5370 12020 6258
rect 12268 6254 12296 6310
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11992 4758 12020 5306
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 12084 4622 12112 6054
rect 12820 4826 12848 8842
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12912 5914 12940 6938
rect 13004 6730 13032 9318
rect 13312 9276 13620 9285
rect 13312 9274 13318 9276
rect 13374 9274 13398 9276
rect 13454 9274 13478 9276
rect 13534 9274 13558 9276
rect 13614 9274 13620 9276
rect 13374 9222 13376 9274
rect 13556 9222 13558 9274
rect 13312 9220 13318 9222
rect 13374 9220 13398 9222
rect 13454 9220 13478 9222
rect 13534 9220 13558 9222
rect 13614 9220 13620 9222
rect 13312 9211 13620 9220
rect 13832 9178 13860 12242
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13312 8188 13620 8197
rect 13312 8186 13318 8188
rect 13374 8186 13398 8188
rect 13454 8186 13478 8188
rect 13534 8186 13558 8188
rect 13614 8186 13620 8188
rect 13374 8134 13376 8186
rect 13556 8134 13558 8186
rect 13312 8132 13318 8134
rect 13374 8132 13398 8134
rect 13454 8132 13478 8134
rect 13534 8132 13558 8134
rect 13614 8132 13620 8134
rect 13312 8123 13620 8132
rect 13832 7410 13860 9114
rect 13924 8294 13952 9930
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7886 13952 8230
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13312 7100 13620 7109
rect 13312 7098 13318 7100
rect 13374 7098 13398 7100
rect 13454 7098 13478 7100
rect 13534 7098 13558 7100
rect 13614 7098 13620 7100
rect 13374 7046 13376 7098
rect 13556 7046 13558 7098
rect 13312 7044 13318 7046
rect 13374 7044 13398 7046
rect 13454 7044 13478 7046
rect 13534 7044 13558 7046
rect 13614 7044 13620 7046
rect 13312 7035 13620 7044
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13004 5302 13032 6054
rect 13096 5778 13124 6190
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13188 5692 13216 6394
rect 13312 6012 13620 6021
rect 13312 6010 13318 6012
rect 13374 6010 13398 6012
rect 13454 6010 13478 6012
rect 13534 6010 13558 6012
rect 13614 6010 13620 6012
rect 13374 5958 13376 6010
rect 13556 5958 13558 6010
rect 13312 5956 13318 5958
rect 13374 5956 13398 5958
rect 13454 5956 13478 5958
rect 13534 5956 13558 5958
rect 13614 5956 13620 5958
rect 13312 5947 13620 5956
rect 13648 5914 13676 7142
rect 13740 6934 13768 7278
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 6458 13768 6598
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13832 6186 13860 7346
rect 13924 6798 13952 7822
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6254 13952 6734
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13268 5704 13320 5710
rect 13188 5664 13268 5692
rect 13268 5646 13320 5652
rect 13280 5370 13308 5646
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13268 5364 13320 5370
rect 13188 5324 13268 5352
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13004 4758 13032 5238
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 10839 4380 11147 4389
rect 10839 4378 10845 4380
rect 10901 4378 10925 4380
rect 10981 4378 11005 4380
rect 11061 4378 11085 4380
rect 11141 4378 11147 4380
rect 10901 4326 10903 4378
rect 11083 4326 11085 4378
rect 10839 4324 10845 4326
rect 10901 4324 10925 4326
rect 10981 4324 11005 4326
rect 11061 4324 11085 4326
rect 11141 4324 11147 4326
rect 10839 4315 11147 4324
rect 11900 4214 11928 4558
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 12084 4146 12112 4558
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12176 4214 12204 4490
rect 13004 4282 13032 4558
rect 13188 4554 13216 5324
rect 13268 5306 13320 5312
rect 13312 4924 13620 4933
rect 13312 4922 13318 4924
rect 13374 4922 13398 4924
rect 13454 4922 13478 4924
rect 13534 4922 13558 4924
rect 13614 4922 13620 4924
rect 13374 4870 13376 4922
rect 13556 4870 13558 4922
rect 13312 4868 13318 4870
rect 13374 4868 13398 4870
rect 13454 4868 13478 4870
rect 13534 4868 13558 4870
rect 13614 4868 13620 4870
rect 13312 4859 13620 4868
rect 13648 4826 13676 5578
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14016 4826 14044 5170
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 13188 4146 13216 4490
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 13312 3836 13620 3845
rect 13312 3834 13318 3836
rect 13374 3834 13398 3836
rect 13454 3834 13478 3836
rect 13534 3834 13558 3836
rect 13614 3834 13620 3836
rect 13374 3782 13376 3834
rect 13556 3782 13558 3834
rect 13312 3780 13318 3782
rect 13374 3780 13398 3782
rect 13454 3780 13478 3782
rect 13534 3780 13558 3782
rect 13614 3780 13620 3782
rect 13312 3771 13620 3780
rect 10839 3292 11147 3301
rect 10839 3290 10845 3292
rect 10901 3290 10925 3292
rect 10981 3290 11005 3292
rect 11061 3290 11085 3292
rect 11141 3290 11147 3292
rect 10901 3238 10903 3290
rect 11083 3238 11085 3290
rect 10839 3236 10845 3238
rect 10901 3236 10925 3238
rect 10981 3236 11005 3238
rect 11061 3236 11085 3238
rect 11141 3236 11147 3238
rect 10839 3227 11147 3236
rect 13312 2748 13620 2757
rect 13312 2746 13318 2748
rect 13374 2746 13398 2748
rect 13454 2746 13478 2748
rect 13534 2746 13558 2748
rect 13614 2746 13620 2748
rect 13374 2694 13376 2746
rect 13556 2694 13558 2746
rect 13312 2692 13318 2694
rect 13374 2692 13398 2694
rect 13454 2692 13478 2694
rect 13534 2692 13558 2694
rect 13614 2692 13620 2694
rect 13312 2683 13620 2692
rect 14108 2446 14136 9522
rect 14200 8090 14228 17682
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14292 16114 14320 16934
rect 14738 16552 14794 16561
rect 14738 16487 14740 16496
rect 14792 16487 14794 16496
rect 14740 16458 14792 16464
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14292 13802 14320 16050
rect 14476 15638 14504 16050
rect 14464 15632 14516 15638
rect 14464 15574 14516 15580
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 14278 14688 14418
rect 14844 14396 14872 18022
rect 14936 17814 14964 18226
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 15028 17746 15056 18226
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 15396 17610 15424 19110
rect 15660 18692 15712 18698
rect 15660 18634 15712 18640
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15580 17746 15608 18226
rect 15672 18170 15700 18634
rect 15784 18524 16092 18533
rect 15784 18522 15790 18524
rect 15846 18522 15870 18524
rect 15926 18522 15950 18524
rect 16006 18522 16030 18524
rect 16086 18522 16092 18524
rect 15846 18470 15848 18522
rect 16028 18470 16030 18522
rect 15784 18468 15790 18470
rect 15846 18468 15870 18470
rect 15926 18468 15950 18470
rect 16006 18468 16030 18470
rect 16086 18468 16092 18470
rect 15784 18459 16092 18468
rect 16224 18222 16252 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16592 18698 16620 19178
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17236 18766 17264 19110
rect 17512 18766 17540 19110
rect 18257 19068 18565 19077
rect 18257 19066 18263 19068
rect 18319 19066 18343 19068
rect 18399 19066 18423 19068
rect 18479 19066 18503 19068
rect 18559 19066 18565 19068
rect 18319 19014 18321 19066
rect 18501 19014 18503 19066
rect 18257 19012 18263 19014
rect 18319 19012 18343 19014
rect 18399 19012 18423 19014
rect 18479 19012 18503 19014
rect 18559 19012 18565 19014
rect 18257 19003 18565 19012
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 19352 18698 19380 19246
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16212 18216 16264 18222
rect 15672 18142 15884 18170
rect 16212 18158 16264 18164
rect 15856 18086 15884 18142
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15396 17202 15424 17546
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14936 14550 14964 16526
rect 15028 15570 15056 16526
rect 15120 15994 15148 16934
rect 15580 16114 15608 17682
rect 15856 17610 15884 18022
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15784 17436 16092 17445
rect 15784 17434 15790 17436
rect 15846 17434 15870 17436
rect 15926 17434 15950 17436
rect 16006 17434 16030 17436
rect 16086 17434 16092 17436
rect 15846 17382 15848 17434
rect 16028 17382 16030 17434
rect 15784 17380 15790 17382
rect 15846 17380 15870 17382
rect 15926 17380 15950 17382
rect 16006 17380 16030 17382
rect 16086 17380 16092 17382
rect 15784 17371 16092 17380
rect 15784 16348 16092 16357
rect 15784 16346 15790 16348
rect 15846 16346 15870 16348
rect 15926 16346 15950 16348
rect 16006 16346 16030 16348
rect 16086 16346 16092 16348
rect 15846 16294 15848 16346
rect 16028 16294 16030 16346
rect 15784 16292 15790 16294
rect 15846 16292 15870 16294
rect 15926 16292 15950 16294
rect 16006 16292 16030 16294
rect 16086 16292 16092 16294
rect 15784 16283 16092 16292
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15200 16040 15252 16046
rect 15120 15988 15200 15994
rect 15120 15982 15252 15988
rect 15120 15966 15240 15982
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15120 15502 15148 15846
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 15016 14408 15068 14414
rect 14844 14368 14964 14396
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14660 10674 14688 14214
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14752 12170 14780 12582
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14476 8838 14504 9114
rect 14568 8838 14596 10406
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14660 8430 14688 10610
rect 14752 9586 14780 11834
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14752 8634 14780 9046
rect 14844 8974 14872 14214
rect 14936 13938 14964 14368
rect 15120 14396 15148 15438
rect 15304 14414 15332 15506
rect 15784 15260 16092 15269
rect 15784 15258 15790 15260
rect 15846 15258 15870 15260
rect 15926 15258 15950 15260
rect 16006 15258 16030 15260
rect 16086 15258 16092 15260
rect 15846 15206 15848 15258
rect 16028 15206 16030 15258
rect 15784 15204 15790 15206
rect 15846 15204 15870 15206
rect 15926 15204 15950 15206
rect 16006 15204 16030 15206
rect 16086 15204 16092 15206
rect 15784 15195 16092 15204
rect 15476 14884 15528 14890
rect 15476 14826 15528 14832
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 14550 15424 14758
rect 15488 14618 15516 14826
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15068 14368 15148 14396
rect 15292 14408 15344 14414
rect 15016 14350 15068 14356
rect 15292 14350 15344 14356
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15212 13870 15240 14214
rect 15304 13938 15332 14350
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 12442 15240 13670
rect 15304 12442 15332 13738
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 11762 15148 12106
rect 15396 12102 15424 12582
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14936 10810 14964 11698
rect 15488 11642 15516 14554
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15784 14172 16092 14181
rect 15784 14170 15790 14172
rect 15846 14170 15870 14172
rect 15926 14170 15950 14172
rect 16006 14170 16030 14172
rect 16086 14170 16092 14172
rect 15846 14118 15848 14170
rect 16028 14118 16030 14170
rect 15784 14116 15790 14118
rect 15846 14116 15870 14118
rect 15926 14116 15950 14118
rect 16006 14116 16030 14118
rect 16086 14116 16092 14118
rect 15784 14107 16092 14116
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15580 11898 15608 12310
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15292 11620 15344 11626
rect 15488 11614 15608 11642
rect 15292 11562 15344 11568
rect 15120 11082 15148 11562
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 15120 10606 15148 11018
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14936 10062 14964 10406
rect 15120 10198 15148 10542
rect 15304 10266 15332 11562
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11286 15516 11494
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 14936 9178 14964 9658
rect 15028 9178 15056 9862
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 5710 14228 7890
rect 14936 7886 14964 9114
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15028 8634 15056 8774
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15120 8566 15148 9998
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9518 15240 9862
rect 15304 9518 15332 10202
rect 15396 9722 15424 10406
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9042 15332 9318
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15488 8566 15516 11222
rect 15580 10266 15608 11614
rect 15672 11558 15700 13806
rect 15784 13084 16092 13093
rect 15784 13082 15790 13084
rect 15846 13082 15870 13084
rect 15926 13082 15950 13084
rect 16006 13082 16030 13084
rect 16086 13082 16092 13084
rect 15846 13030 15848 13082
rect 16028 13030 16030 13082
rect 15784 13028 15790 13030
rect 15846 13028 15870 13030
rect 15926 13028 15950 13030
rect 16006 13028 16030 13030
rect 16086 13028 16092 13030
rect 15784 13019 16092 13028
rect 16132 12238 16160 14214
rect 16224 12374 16252 18158
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16316 16114 16344 17546
rect 16592 17542 16620 18294
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16684 17610 16712 18226
rect 16960 17678 16988 18226
rect 17052 18222 17080 18634
rect 17868 18352 17920 18358
rect 17868 18294 17920 18300
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17052 17814 17080 18158
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 16726 16620 17478
rect 16856 17060 16908 17066
rect 16856 17002 16908 17008
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16592 16046 16620 16458
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16776 15978 16804 16526
rect 16868 16454 16896 17002
rect 16960 16590 16988 17614
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16868 16114 16896 16390
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16684 14414 16712 15370
rect 16868 15042 16896 16050
rect 16960 15570 16988 16050
rect 17052 15722 17080 17750
rect 17880 17610 17908 18294
rect 19352 18086 19380 18634
rect 20729 18524 21037 18533
rect 20729 18522 20735 18524
rect 20791 18522 20815 18524
rect 20871 18522 20895 18524
rect 20951 18522 20975 18524
rect 21031 18522 21037 18524
rect 20791 18470 20793 18522
rect 20973 18470 20975 18522
rect 20729 18468 20735 18470
rect 20791 18468 20815 18470
rect 20871 18468 20895 18470
rect 20951 18468 20975 18470
rect 21031 18468 21037 18470
rect 20729 18459 21037 18468
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 18257 17980 18565 17989
rect 18257 17978 18263 17980
rect 18319 17978 18343 17980
rect 18399 17978 18423 17980
rect 18479 17978 18503 17980
rect 18559 17978 18565 17980
rect 18319 17926 18321 17978
rect 18501 17926 18503 17978
rect 18257 17924 18263 17926
rect 18319 17924 18343 17926
rect 18399 17924 18423 17926
rect 18479 17924 18503 17926
rect 18559 17924 18565 17926
rect 18257 17915 18565 17924
rect 19352 17610 19380 18022
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17420 15994 17448 16458
rect 17512 16046 17540 17070
rect 18257 16892 18565 16901
rect 18257 16890 18263 16892
rect 18319 16890 18343 16892
rect 18399 16890 18423 16892
rect 18479 16890 18503 16892
rect 18559 16890 18565 16892
rect 18319 16838 18321 16890
rect 18501 16838 18503 16890
rect 18257 16836 18263 16838
rect 18319 16836 18343 16838
rect 18399 16836 18423 16838
rect 18479 16836 18503 16838
rect 18559 16836 18565 16838
rect 18257 16827 18565 16836
rect 18142 16688 18198 16697
rect 19444 16674 19472 17478
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 18142 16623 18198 16632
rect 19352 16646 19472 16674
rect 19536 16658 19564 17138
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19524 16652 19576 16658
rect 18156 16590 18184 16623
rect 19352 16590 19380 16646
rect 19524 16594 19576 16600
rect 18144 16584 18196 16590
rect 18050 16552 18106 16561
rect 18144 16526 18196 16532
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 18050 16487 18052 16496
rect 18104 16487 18106 16496
rect 18052 16458 18104 16464
rect 19536 16454 19564 16594
rect 19628 16590 19656 16934
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 17696 16114 17724 16390
rect 19536 16114 19564 16390
rect 19720 16182 19748 17138
rect 19812 16726 19840 17546
rect 20729 17436 21037 17445
rect 20729 17434 20735 17436
rect 20791 17434 20815 17436
rect 20871 17434 20895 17436
rect 20951 17434 20975 17436
rect 21031 17434 21037 17436
rect 20791 17382 20793 17434
rect 20973 17382 20975 17434
rect 20729 17380 20735 17382
rect 20791 17380 20815 17382
rect 20871 17380 20895 17382
rect 20951 17380 20975 17382
rect 21031 17380 21037 17382
rect 20729 17371 21037 17380
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19812 16250 19840 16526
rect 20729 16348 21037 16357
rect 20729 16346 20735 16348
rect 20791 16346 20815 16348
rect 20871 16346 20895 16348
rect 20951 16346 20975 16348
rect 21031 16346 21037 16348
rect 20791 16294 20793 16346
rect 20973 16294 20975 16346
rect 20729 16292 20735 16294
rect 20791 16292 20815 16294
rect 20871 16292 20895 16294
rect 20951 16292 20975 16294
rect 21031 16292 21037 16294
rect 20729 16283 21037 16292
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 17328 15966 17448 15994
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17328 15910 17356 15966
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17052 15694 17172 15722
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16776 15014 16896 15042
rect 16948 15020 17000 15026
rect 16776 14618 16804 15014
rect 16948 14962 17000 14968
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16592 14074 16620 14350
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16868 13326 16896 14894
rect 16960 14074 16988 14962
rect 17052 14414 17080 15574
rect 17144 14618 17172 15694
rect 17328 15434 17356 15846
rect 17316 15428 17368 15434
rect 17316 15370 17368 15376
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15784 11996 16092 12005
rect 15784 11994 15790 11996
rect 15846 11994 15870 11996
rect 15926 11994 15950 11996
rect 16006 11994 16030 11996
rect 16086 11994 16092 11996
rect 15846 11942 15848 11994
rect 16028 11942 16030 11994
rect 15784 11940 15790 11942
rect 15846 11940 15870 11942
rect 15926 11940 15950 11942
rect 16006 11940 16030 11942
rect 16086 11940 16092 11942
rect 15784 11931 16092 11940
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15784 10908 16092 10917
rect 15784 10906 15790 10908
rect 15846 10906 15870 10908
rect 15926 10906 15950 10908
rect 16006 10906 16030 10908
rect 16086 10906 16092 10908
rect 15846 10854 15848 10906
rect 16028 10854 16030 10906
rect 15784 10852 15790 10854
rect 15846 10852 15870 10854
rect 15926 10852 15950 10854
rect 16006 10852 16030 10854
rect 16086 10852 16092 10854
rect 15784 10843 16092 10852
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15580 8922 15608 10202
rect 15784 9820 16092 9829
rect 15784 9818 15790 9820
rect 15846 9818 15870 9820
rect 15926 9818 15950 9820
rect 16006 9818 16030 9820
rect 16086 9818 16092 9820
rect 15846 9766 15848 9818
rect 16028 9766 16030 9818
rect 15784 9764 15790 9766
rect 15846 9764 15870 9766
rect 15926 9764 15950 9766
rect 16006 9764 16030 9766
rect 16086 9764 16092 9766
rect 15784 9755 16092 9764
rect 15580 8894 15700 8922
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15028 7818 15056 8434
rect 15580 7954 15608 8774
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15028 7410 15056 7754
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6798 14320 7142
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14476 6089 14504 7278
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 14462 6080 14518 6089
rect 14462 6015 14518 6024
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5234 14228 5646
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14476 4486 14504 6015
rect 15028 5234 15056 6666
rect 15120 5778 15148 7822
rect 15580 7478 15608 7890
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15672 7410 15700 8894
rect 15784 8732 16092 8741
rect 15784 8730 15790 8732
rect 15846 8730 15870 8732
rect 15926 8730 15950 8732
rect 16006 8730 16030 8732
rect 16086 8730 16092 8732
rect 15846 8678 15848 8730
rect 16028 8678 16030 8730
rect 15784 8676 15790 8678
rect 15846 8676 15870 8678
rect 15926 8676 15950 8678
rect 16006 8676 16030 8678
rect 16086 8676 16092 8678
rect 15784 8667 16092 8676
rect 16132 8514 16160 12174
rect 16224 11150 16252 12310
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16132 8486 16252 8514
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 15784 7644 16092 7653
rect 15784 7642 15790 7644
rect 15846 7642 15870 7644
rect 15926 7642 15950 7644
rect 16006 7642 16030 7644
rect 16086 7642 16092 7644
rect 15846 7590 15848 7642
rect 16028 7590 16030 7642
rect 15784 7588 15790 7590
rect 15846 7588 15870 7590
rect 15926 7588 15950 7590
rect 16006 7588 16030 7590
rect 16086 7588 16092 7590
rect 15784 7579 16092 7588
rect 16132 7410 16160 8298
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 15672 6662 15700 7346
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15784 6556 16092 6565
rect 15784 6554 15790 6556
rect 15846 6554 15870 6556
rect 15926 6554 15950 6556
rect 16006 6554 16030 6556
rect 16086 6554 16092 6556
rect 15846 6502 15848 6554
rect 16028 6502 16030 6554
rect 15784 6500 15790 6502
rect 15846 6500 15870 6502
rect 15926 6500 15950 6502
rect 16006 6500 16030 6502
rect 16086 6500 16092 6502
rect 15784 6491 16092 6500
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 5846 15332 6190
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 16132 5778 16160 7346
rect 16224 6934 16252 8486
rect 16592 7954 16620 12106
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16684 11354 16712 11562
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16304 6384 16356 6390
rect 16408 6361 16436 6734
rect 16304 6326 16356 6332
rect 16394 6352 16450 6361
rect 16316 6186 16344 6326
rect 16394 6287 16450 6296
rect 16488 6316 16540 6322
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15028 4690 15056 5170
rect 15580 4758 15608 5170
rect 15672 5166 15700 5510
rect 15784 5468 16092 5477
rect 15784 5466 15790 5468
rect 15846 5466 15870 5468
rect 15926 5466 15950 5468
rect 16006 5466 16030 5468
rect 16086 5466 16092 5468
rect 15846 5414 15848 5466
rect 16028 5414 16030 5466
rect 15784 5412 15790 5414
rect 15846 5412 15870 5414
rect 15926 5412 15950 5414
rect 16006 5412 16030 5414
rect 16086 5412 16092 5414
rect 15784 5403 16092 5412
rect 16132 5302 16160 5510
rect 16408 5302 16436 6287
rect 16488 6258 16540 6264
rect 16500 5710 16528 6258
rect 16684 6186 16712 11086
rect 16868 10198 16896 13262
rect 17052 11286 17080 14350
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17144 13530 17172 13942
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17236 12918 17264 13670
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17236 11506 17264 12106
rect 17328 11626 17356 14214
rect 17512 12434 17540 15982
rect 17604 15706 17632 16050
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17696 15638 17724 16050
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 18257 15804 18565 15813
rect 18257 15802 18263 15804
rect 18319 15802 18343 15804
rect 18399 15802 18423 15804
rect 18479 15802 18503 15804
rect 18559 15802 18565 15804
rect 18319 15750 18321 15802
rect 18501 15750 18503 15802
rect 18257 15748 18263 15750
rect 18319 15748 18343 15750
rect 18399 15748 18423 15750
rect 18479 15748 18503 15750
rect 18559 15748 18565 15750
rect 18257 15739 18565 15748
rect 19444 15706 19472 15982
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17880 15570 17908 15642
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17776 14408 17828 14414
rect 17880 14396 17908 15506
rect 19536 15434 19564 16050
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19536 15026 19564 15370
rect 20729 15260 21037 15269
rect 20729 15258 20735 15260
rect 20791 15258 20815 15260
rect 20871 15258 20895 15260
rect 20951 15258 20975 15260
rect 21031 15258 21037 15260
rect 20791 15206 20793 15258
rect 20973 15206 20975 15258
rect 20729 15204 20735 15206
rect 20791 15204 20815 15206
rect 20871 15204 20895 15206
rect 20951 15204 20975 15206
rect 21031 15204 21037 15206
rect 20729 15195 21037 15204
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 18257 14716 18565 14725
rect 18257 14714 18263 14716
rect 18319 14714 18343 14716
rect 18399 14714 18423 14716
rect 18479 14714 18503 14716
rect 18559 14714 18565 14716
rect 18319 14662 18321 14714
rect 18501 14662 18503 14714
rect 18257 14660 18263 14662
rect 18319 14660 18343 14662
rect 18399 14660 18423 14662
rect 18479 14660 18503 14662
rect 18559 14660 18565 14662
rect 18257 14651 18565 14660
rect 19536 14618 19564 14962
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 17828 14368 17908 14396
rect 17776 14350 17828 14356
rect 17788 13802 17816 14350
rect 18432 14006 18460 14486
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18616 14006 18644 14350
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17788 13190 17816 13738
rect 18257 13628 18565 13637
rect 18257 13626 18263 13628
rect 18319 13626 18343 13628
rect 18399 13626 18423 13628
rect 18479 13626 18503 13628
rect 18559 13626 18565 13628
rect 18319 13574 18321 13626
rect 18501 13574 18503 13626
rect 18257 13572 18263 13574
rect 18319 13572 18343 13574
rect 18399 13572 18423 13574
rect 18479 13572 18503 13574
rect 18559 13572 18565 13574
rect 18257 13563 18565 13572
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17512 12406 17632 12434
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17236 11478 17356 11506
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 17052 9110 17080 11222
rect 17328 11218 17356 11478
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8498 16804 8774
rect 17052 8634 17080 8842
rect 17144 8634 17172 10678
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17236 9722 17264 9862
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17328 9586 17356 11154
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17420 9568 17448 9862
rect 17500 9580 17552 9586
rect 17420 9540 17500 9568
rect 17236 9178 17264 9522
rect 17420 9178 17448 9540
rect 17500 9522 17552 9528
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17052 8514 17080 8570
rect 17236 8514 17264 9114
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17328 8548 17356 9046
rect 17408 8560 17460 8566
rect 17328 8520 17408 8548
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16960 8486 17080 8514
rect 17144 8498 17264 8514
rect 17408 8502 17460 8508
rect 17132 8492 17264 8498
rect 16776 7342 16804 8434
rect 16960 8294 16988 8486
rect 17184 8486 17264 8492
rect 17132 8434 17184 8440
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16960 8090 16988 8230
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16868 7410 16896 7686
rect 16960 7546 16988 7686
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17052 7410 17080 8298
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15672 4554 15700 5102
rect 16132 4690 16160 5238
rect 17144 5098 17172 7482
rect 17328 7478 17356 7890
rect 17420 7886 17448 8502
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17328 6798 17356 7414
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6798 17540 7142
rect 17604 6798 17632 12406
rect 17788 12102 17816 12854
rect 17972 12714 18000 13262
rect 18616 12850 18644 13942
rect 18708 13734 18736 14418
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17972 12442 18000 12650
rect 18257 12540 18565 12549
rect 18257 12538 18263 12540
rect 18319 12538 18343 12540
rect 18399 12538 18423 12540
rect 18479 12538 18503 12540
rect 18559 12538 18565 12540
rect 18319 12486 18321 12538
rect 18501 12486 18503 12538
rect 18257 12484 18263 12486
rect 18319 12484 18343 12486
rect 18399 12484 18423 12486
rect 18479 12484 18503 12486
rect 18559 12484 18565 12486
rect 18257 12475 18565 12484
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 7410 17724 11494
rect 17788 11218 17816 12038
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17788 10742 17816 11154
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17788 7954 17816 10678
rect 17972 10470 18000 12174
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 9654 18000 10406
rect 18064 10062 18092 12310
rect 18616 11898 18644 12786
rect 18708 12782 18736 13670
rect 19168 12850 19196 14486
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19352 13530 19380 14282
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 13938 19564 14214
rect 19720 13938 19748 14758
rect 20729 14172 21037 14181
rect 20729 14170 20735 14172
rect 20791 14170 20815 14172
rect 20871 14170 20895 14172
rect 20951 14170 20975 14172
rect 21031 14170 21037 14172
rect 20791 14118 20793 14170
rect 20973 14118 20975 14170
rect 20729 14116 20735 14118
rect 20791 14116 20815 14118
rect 20871 14116 20895 14118
rect 20951 14116 20975 14118
rect 21031 14116 21037 14118
rect 20729 14107 21037 14116
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19260 12850 19288 13126
rect 19628 12986 19656 13466
rect 19720 13190 19748 13738
rect 19996 13462 20024 13942
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18696 12776 18748 12782
rect 18748 12724 18828 12730
rect 18696 12718 18828 12724
rect 18708 12702 18828 12718
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12442 18736 12582
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18800 11762 18828 12702
rect 19352 12374 19380 12854
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19628 11898 19656 12718
rect 19720 12442 19748 13126
rect 20729 13084 21037 13093
rect 20729 13082 20735 13084
rect 20791 13082 20815 13084
rect 20871 13082 20895 13084
rect 20951 13082 20975 13084
rect 21031 13082 21037 13084
rect 20791 13030 20793 13082
rect 20973 13030 20975 13082
rect 20729 13028 20735 13030
rect 20791 13028 20815 13030
rect 20871 13028 20895 13030
rect 20951 13028 20975 13030
rect 21031 13028 21037 13030
rect 20729 13019 21037 13028
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19996 12442 20024 12650
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19720 12170 19748 12378
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11898 19840 12038
rect 20729 11996 21037 12005
rect 20729 11994 20735 11996
rect 20791 11994 20815 11996
rect 20871 11994 20895 11996
rect 20951 11994 20975 11996
rect 21031 11994 21037 11996
rect 20791 11942 20793 11994
rect 20973 11942 20975 11994
rect 20729 11940 20735 11942
rect 20791 11940 20815 11942
rect 20871 11940 20895 11942
rect 20951 11940 20975 11942
rect 21031 11940 21037 11942
rect 20729 11931 21037 11940
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18257 11452 18565 11461
rect 18257 11450 18263 11452
rect 18319 11450 18343 11452
rect 18399 11450 18423 11452
rect 18479 11450 18503 11452
rect 18559 11450 18565 11452
rect 18319 11398 18321 11450
rect 18501 11398 18503 11450
rect 18257 11396 18263 11398
rect 18319 11396 18343 11398
rect 18399 11396 18423 11398
rect 18479 11396 18503 11398
rect 18559 11396 18565 11398
rect 18257 11387 18565 11396
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18524 11234 18552 11290
rect 18616 11234 18644 11698
rect 18524 11206 18644 11234
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18156 10674 18184 11086
rect 18524 11082 18552 11206
rect 18800 11150 18828 11698
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10810 18552 11018
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18616 10742 18644 10950
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 19444 10674 19472 11630
rect 19628 11354 19656 11834
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 18156 10266 18184 10610
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18257 10364 18565 10373
rect 18257 10362 18263 10364
rect 18319 10362 18343 10364
rect 18399 10362 18423 10364
rect 18479 10362 18503 10364
rect 18559 10362 18565 10364
rect 18319 10310 18321 10362
rect 18501 10310 18503 10362
rect 18257 10308 18263 10310
rect 18319 10308 18343 10310
rect 18399 10308 18423 10310
rect 18479 10308 18503 10310
rect 18559 10308 18565 10310
rect 18257 10299 18565 10308
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 18156 9586 18184 10066
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18257 9276 18565 9285
rect 18257 9274 18263 9276
rect 18319 9274 18343 9276
rect 18399 9274 18423 9276
rect 18479 9274 18503 9276
rect 18559 9274 18565 9276
rect 18319 9222 18321 9274
rect 18501 9222 18503 9274
rect 18257 9220 18263 9222
rect 18319 9220 18343 9222
rect 18399 9220 18423 9222
rect 18479 9220 18503 9222
rect 18559 9220 18565 9222
rect 18257 9211 18565 9220
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17328 6390 17356 6734
rect 17512 6458 17540 6734
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 5778 17264 6258
rect 17604 6118 17632 6734
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17604 5710 17632 6054
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17788 5574 17816 7890
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17880 7274 17908 7414
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17868 6112 17920 6118
rect 17866 6080 17868 6089
rect 17972 6100 18000 8434
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18156 7342 18184 8366
rect 18257 8188 18565 8197
rect 18257 8186 18263 8188
rect 18319 8186 18343 8188
rect 18399 8186 18423 8188
rect 18479 8186 18503 8188
rect 18559 8186 18565 8188
rect 18319 8134 18321 8186
rect 18501 8134 18503 8186
rect 18257 8132 18263 8134
rect 18319 8132 18343 8134
rect 18399 8132 18423 8134
rect 18479 8132 18503 8134
rect 18559 8132 18565 8134
rect 18257 8123 18565 8132
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18064 6458 18092 6734
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18156 6322 18184 7278
rect 18257 7100 18565 7109
rect 18257 7098 18263 7100
rect 18319 7098 18343 7100
rect 18399 7098 18423 7100
rect 18479 7098 18503 7100
rect 18559 7098 18565 7100
rect 18319 7046 18321 7098
rect 18501 7046 18503 7098
rect 18257 7044 18263 7046
rect 18319 7044 18343 7046
rect 18399 7044 18423 7046
rect 18479 7044 18503 7046
rect 18559 7044 18565 7046
rect 18257 7035 18565 7044
rect 18616 6662 18644 10542
rect 19168 9926 19196 10542
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18892 7886 18920 9522
rect 19168 9466 19196 9862
rect 19260 9586 19288 10406
rect 19444 10130 19472 10610
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19444 9654 19472 9862
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19168 9438 19288 9466
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19168 8498 19196 8978
rect 19260 8974 19288 9438
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19260 8430 19288 8910
rect 19628 8634 19656 9522
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 18708 7410 18736 7822
rect 19260 7410 19288 7822
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 17920 6080 18000 6100
rect 17922 6072 18000 6080
rect 17866 6015 17922 6024
rect 18257 6012 18565 6021
rect 18257 6010 18263 6012
rect 18319 6010 18343 6012
rect 18399 6010 18423 6012
rect 18479 6010 18503 6012
rect 18559 6010 18565 6012
rect 18319 5958 18321 6010
rect 18501 5958 18503 6010
rect 18257 5956 18263 5958
rect 18319 5956 18343 5958
rect 18399 5956 18423 5958
rect 18479 5956 18503 5958
rect 18559 5956 18565 5958
rect 18257 5947 18565 5956
rect 18616 5846 18644 6258
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 18257 4924 18565 4933
rect 18257 4922 18263 4924
rect 18319 4922 18343 4924
rect 18399 4922 18423 4924
rect 18479 4922 18503 4924
rect 18559 4922 18565 4924
rect 18319 4870 18321 4922
rect 18501 4870 18503 4922
rect 18257 4868 18263 4870
rect 18319 4868 18343 4870
rect 18399 4868 18423 4870
rect 18479 4868 18503 4870
rect 18559 4868 18565 4870
rect 18257 4859 18565 4868
rect 19260 4758 19288 7346
rect 19352 6458 19380 7754
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19628 7546 19656 7686
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19720 7206 19748 9998
rect 19812 9450 19840 11562
rect 20729 10908 21037 10917
rect 20729 10906 20735 10908
rect 20791 10906 20815 10908
rect 20871 10906 20895 10908
rect 20951 10906 20975 10908
rect 21031 10906 21037 10908
rect 20791 10854 20793 10906
rect 20973 10854 20975 10906
rect 20729 10852 20735 10854
rect 20791 10852 20815 10854
rect 20871 10852 20895 10854
rect 20951 10852 20975 10854
rect 21031 10852 21037 10854
rect 20729 10843 21037 10852
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 19904 10062 19932 10678
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 20729 9820 21037 9829
rect 20729 9818 20735 9820
rect 20791 9818 20815 9820
rect 20871 9818 20895 9820
rect 20951 9818 20975 9820
rect 21031 9818 21037 9820
rect 20791 9766 20793 9818
rect 20973 9766 20975 9818
rect 20729 9764 20735 9766
rect 20791 9764 20815 9766
rect 20871 9764 20895 9766
rect 20951 9764 20975 9766
rect 21031 9764 21037 9766
rect 20729 9755 21037 9764
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19904 9178 19932 9522
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 20729 8732 21037 8741
rect 20729 8730 20735 8732
rect 20791 8730 20815 8732
rect 20871 8730 20895 8732
rect 20951 8730 20975 8732
rect 21031 8730 21037 8732
rect 20791 8678 20793 8730
rect 20973 8678 20975 8730
rect 20729 8676 20735 8678
rect 20791 8676 20815 8678
rect 20871 8676 20895 8678
rect 20951 8676 20975 8678
rect 21031 8676 21037 8678
rect 20729 8667 21037 8676
rect 20729 7644 21037 7653
rect 20729 7642 20735 7644
rect 20791 7642 20815 7644
rect 20871 7642 20895 7644
rect 20951 7642 20975 7644
rect 21031 7642 21037 7644
rect 20791 7590 20793 7642
rect 20973 7590 20975 7642
rect 20729 7588 20735 7590
rect 20791 7588 20815 7590
rect 20871 7588 20895 7590
rect 20951 7588 20975 7590
rect 21031 7588 21037 7590
rect 20729 7579 21037 7588
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 20729 6556 21037 6565
rect 20729 6554 20735 6556
rect 20791 6554 20815 6556
rect 20871 6554 20895 6556
rect 20951 6554 20975 6556
rect 21031 6554 21037 6556
rect 20791 6502 20793 6554
rect 20973 6502 20975 6554
rect 20729 6500 20735 6502
rect 20791 6500 20815 6502
rect 20871 6500 20895 6502
rect 20951 6500 20975 6502
rect 21031 6500 21037 6502
rect 20729 6491 21037 6500
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 15784 4380 16092 4389
rect 15784 4378 15790 4380
rect 15846 4378 15870 4380
rect 15926 4378 15950 4380
rect 16006 4378 16030 4380
rect 16086 4378 16092 4380
rect 15846 4326 15848 4378
rect 16028 4326 16030 4378
rect 15784 4324 15790 4326
rect 15846 4324 15870 4326
rect 15926 4324 15950 4326
rect 16006 4324 16030 4326
rect 16086 4324 16092 4326
rect 15784 4315 16092 4324
rect 18257 3836 18565 3845
rect 18257 3834 18263 3836
rect 18319 3834 18343 3836
rect 18399 3834 18423 3836
rect 18479 3834 18503 3836
rect 18559 3834 18565 3836
rect 18319 3782 18321 3834
rect 18501 3782 18503 3834
rect 18257 3780 18263 3782
rect 18319 3780 18343 3782
rect 18399 3780 18423 3782
rect 18479 3780 18503 3782
rect 18559 3780 18565 3782
rect 18257 3771 18565 3780
rect 15784 3292 16092 3301
rect 15784 3290 15790 3292
rect 15846 3290 15870 3292
rect 15926 3290 15950 3292
rect 16006 3290 16030 3292
rect 16086 3290 16092 3292
rect 15846 3238 15848 3290
rect 16028 3238 16030 3290
rect 15784 3236 15790 3238
rect 15846 3236 15870 3238
rect 15926 3236 15950 3238
rect 16006 3236 16030 3238
rect 16086 3236 16092 3238
rect 15784 3227 16092 3236
rect 18257 2748 18565 2757
rect 18257 2746 18263 2748
rect 18319 2746 18343 2748
rect 18399 2746 18423 2748
rect 18479 2746 18503 2748
rect 18559 2746 18565 2748
rect 18319 2694 18321 2746
rect 18501 2694 18503 2746
rect 18257 2692 18263 2694
rect 18319 2692 18343 2694
rect 18399 2692 18423 2694
rect 18479 2692 18503 2694
rect 18559 2692 18565 2694
rect 18257 2683 18565 2692
rect 19904 2446 19932 6190
rect 20729 5468 21037 5477
rect 20729 5466 20735 5468
rect 20791 5466 20815 5468
rect 20871 5466 20895 5468
rect 20951 5466 20975 5468
rect 21031 5466 21037 5468
rect 20791 5414 20793 5466
rect 20973 5414 20975 5466
rect 20729 5412 20735 5414
rect 20791 5412 20815 5414
rect 20871 5412 20895 5414
rect 20951 5412 20975 5414
rect 21031 5412 21037 5414
rect 20729 5403 21037 5412
rect 20729 4380 21037 4389
rect 20729 4378 20735 4380
rect 20791 4378 20815 4380
rect 20871 4378 20895 4380
rect 20951 4378 20975 4380
rect 21031 4378 21037 4380
rect 20791 4326 20793 4378
rect 20973 4326 20975 4378
rect 20729 4324 20735 4326
rect 20791 4324 20815 4326
rect 20871 4324 20895 4326
rect 20951 4324 20975 4326
rect 21031 4324 21037 4326
rect 20729 4315 21037 4324
rect 20729 3292 21037 3301
rect 20729 3290 20735 3292
rect 20791 3290 20815 3292
rect 20871 3290 20895 3292
rect 20951 3290 20975 3292
rect 21031 3290 21037 3292
rect 20791 3238 20793 3290
rect 20973 3238 20975 3290
rect 20729 3236 20735 3238
rect 20791 3236 20815 3238
rect 20871 3236 20895 3238
rect 20951 3236 20975 3238
rect 21031 3236 21037 3238
rect 20729 3227 21037 3236
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 1596 800 1624 2314
rect 4264 800 4292 2314
rect 5894 2204 6202 2213
rect 5894 2202 5900 2204
rect 5956 2202 5980 2204
rect 6036 2202 6060 2204
rect 6116 2202 6140 2204
rect 6196 2202 6202 2204
rect 5956 2150 5958 2202
rect 6138 2150 6140 2202
rect 5894 2148 5900 2150
rect 5956 2148 5980 2150
rect 6036 2148 6060 2150
rect 6116 2148 6140 2150
rect 6196 2148 6202 2150
rect 5894 2139 6202 2148
rect 6932 800 6960 2314
rect 9600 800 9628 2314
rect 10839 2204 11147 2213
rect 10839 2202 10845 2204
rect 10901 2202 10925 2204
rect 10981 2202 11005 2204
rect 11061 2202 11085 2204
rect 11141 2202 11147 2204
rect 10901 2150 10903 2202
rect 11083 2150 11085 2202
rect 10839 2148 10845 2150
rect 10901 2148 10925 2150
rect 10981 2148 11005 2150
rect 11061 2148 11085 2150
rect 11141 2148 11147 2150
rect 10839 2139 11147 2148
rect 12268 800 12296 2314
rect 14936 800 14964 2314
rect 15784 2204 16092 2213
rect 15784 2202 15790 2204
rect 15846 2202 15870 2204
rect 15926 2202 15950 2204
rect 16006 2202 16030 2204
rect 16086 2202 16092 2204
rect 15846 2150 15848 2202
rect 16028 2150 16030 2202
rect 15784 2148 15790 2150
rect 15846 2148 15870 2150
rect 15926 2148 15950 2150
rect 16006 2148 16030 2150
rect 16086 2148 16092 2150
rect 15784 2139 16092 2148
rect 17604 800 17632 2314
rect 20272 800 20300 2314
rect 20729 2204 21037 2213
rect 20729 2202 20735 2204
rect 20791 2202 20815 2204
rect 20871 2202 20895 2204
rect 20951 2202 20975 2204
rect 21031 2202 21037 2204
rect 20791 2150 20793 2202
rect 20973 2150 20975 2202
rect 20729 2148 20735 2150
rect 20791 2148 20815 2150
rect 20871 2148 20895 2150
rect 20951 2148 20975 2150
rect 21031 2148 21037 2150
rect 20729 2139 21037 2148
rect 1582 0 1638 800
rect 4250 0 4306 800
rect 6918 0 6974 800
rect 9586 0 9642 800
rect 12254 0 12310 800
rect 14922 0 14978 800
rect 17590 0 17646 800
rect 20258 0 20314 800
<< via2 >>
rect 3428 19066 3484 19068
rect 3508 19066 3564 19068
rect 3588 19066 3644 19068
rect 3668 19066 3724 19068
rect 3428 19014 3474 19066
rect 3474 19014 3484 19066
rect 3508 19014 3538 19066
rect 3538 19014 3550 19066
rect 3550 19014 3564 19066
rect 3588 19014 3602 19066
rect 3602 19014 3614 19066
rect 3614 19014 3644 19066
rect 3668 19014 3678 19066
rect 3678 19014 3724 19066
rect 3428 19012 3484 19014
rect 3508 19012 3564 19014
rect 3588 19012 3644 19014
rect 3668 19012 3724 19014
rect 3428 17978 3484 17980
rect 3508 17978 3564 17980
rect 3588 17978 3644 17980
rect 3668 17978 3724 17980
rect 3428 17926 3474 17978
rect 3474 17926 3484 17978
rect 3508 17926 3538 17978
rect 3538 17926 3550 17978
rect 3550 17926 3564 17978
rect 3588 17926 3602 17978
rect 3602 17926 3614 17978
rect 3614 17926 3644 17978
rect 3668 17926 3678 17978
rect 3678 17926 3724 17978
rect 3428 17924 3484 17926
rect 3508 17924 3564 17926
rect 3588 17924 3644 17926
rect 3668 17924 3724 17926
rect 3428 16890 3484 16892
rect 3508 16890 3564 16892
rect 3588 16890 3644 16892
rect 3668 16890 3724 16892
rect 3428 16838 3474 16890
rect 3474 16838 3484 16890
rect 3508 16838 3538 16890
rect 3538 16838 3550 16890
rect 3550 16838 3564 16890
rect 3588 16838 3602 16890
rect 3602 16838 3614 16890
rect 3614 16838 3644 16890
rect 3668 16838 3678 16890
rect 3678 16838 3724 16890
rect 3428 16836 3484 16838
rect 3508 16836 3564 16838
rect 3588 16836 3644 16838
rect 3668 16836 3724 16838
rect 5900 19610 5956 19612
rect 5980 19610 6036 19612
rect 6060 19610 6116 19612
rect 6140 19610 6196 19612
rect 5900 19558 5946 19610
rect 5946 19558 5956 19610
rect 5980 19558 6010 19610
rect 6010 19558 6022 19610
rect 6022 19558 6036 19610
rect 6060 19558 6074 19610
rect 6074 19558 6086 19610
rect 6086 19558 6116 19610
rect 6140 19558 6150 19610
rect 6150 19558 6196 19610
rect 5900 19556 5956 19558
rect 5980 19556 6036 19558
rect 6060 19556 6116 19558
rect 6140 19556 6196 19558
rect 10845 19610 10901 19612
rect 10925 19610 10981 19612
rect 11005 19610 11061 19612
rect 11085 19610 11141 19612
rect 10845 19558 10891 19610
rect 10891 19558 10901 19610
rect 10925 19558 10955 19610
rect 10955 19558 10967 19610
rect 10967 19558 10981 19610
rect 11005 19558 11019 19610
rect 11019 19558 11031 19610
rect 11031 19558 11061 19610
rect 11085 19558 11095 19610
rect 11095 19558 11141 19610
rect 10845 19556 10901 19558
rect 10925 19556 10981 19558
rect 11005 19556 11061 19558
rect 11085 19556 11141 19558
rect 3428 15802 3484 15804
rect 3508 15802 3564 15804
rect 3588 15802 3644 15804
rect 3668 15802 3724 15804
rect 3428 15750 3474 15802
rect 3474 15750 3484 15802
rect 3508 15750 3538 15802
rect 3538 15750 3550 15802
rect 3550 15750 3564 15802
rect 3588 15750 3602 15802
rect 3602 15750 3614 15802
rect 3614 15750 3644 15802
rect 3668 15750 3678 15802
rect 3678 15750 3724 15802
rect 3428 15748 3484 15750
rect 3508 15748 3564 15750
rect 3588 15748 3644 15750
rect 3668 15748 3724 15750
rect 8373 19066 8429 19068
rect 8453 19066 8509 19068
rect 8533 19066 8589 19068
rect 8613 19066 8669 19068
rect 8373 19014 8419 19066
rect 8419 19014 8429 19066
rect 8453 19014 8483 19066
rect 8483 19014 8495 19066
rect 8495 19014 8509 19066
rect 8533 19014 8547 19066
rect 8547 19014 8559 19066
rect 8559 19014 8589 19066
rect 8613 19014 8623 19066
rect 8623 19014 8669 19066
rect 8373 19012 8429 19014
rect 8453 19012 8509 19014
rect 8533 19012 8589 19014
rect 8613 19012 8669 19014
rect 13318 19066 13374 19068
rect 13398 19066 13454 19068
rect 13478 19066 13534 19068
rect 13558 19066 13614 19068
rect 13318 19014 13364 19066
rect 13364 19014 13374 19066
rect 13398 19014 13428 19066
rect 13428 19014 13440 19066
rect 13440 19014 13454 19066
rect 13478 19014 13492 19066
rect 13492 19014 13504 19066
rect 13504 19014 13534 19066
rect 13558 19014 13568 19066
rect 13568 19014 13614 19066
rect 13318 19012 13374 19014
rect 13398 19012 13454 19014
rect 13478 19012 13534 19014
rect 13558 19012 13614 19014
rect 5900 18522 5956 18524
rect 5980 18522 6036 18524
rect 6060 18522 6116 18524
rect 6140 18522 6196 18524
rect 5900 18470 5946 18522
rect 5946 18470 5956 18522
rect 5980 18470 6010 18522
rect 6010 18470 6022 18522
rect 6022 18470 6036 18522
rect 6060 18470 6074 18522
rect 6074 18470 6086 18522
rect 6086 18470 6116 18522
rect 6140 18470 6150 18522
rect 6150 18470 6196 18522
rect 5900 18468 5956 18470
rect 5980 18468 6036 18470
rect 6060 18468 6116 18470
rect 6140 18468 6196 18470
rect 8206 18300 8208 18320
rect 8208 18300 8260 18320
rect 8260 18300 8262 18320
rect 8206 18264 8262 18300
rect 10845 18522 10901 18524
rect 10925 18522 10981 18524
rect 11005 18522 11061 18524
rect 11085 18522 11141 18524
rect 10845 18470 10891 18522
rect 10891 18470 10901 18522
rect 10925 18470 10955 18522
rect 10955 18470 10967 18522
rect 10967 18470 10981 18522
rect 11005 18470 11019 18522
rect 11019 18470 11031 18522
rect 11031 18470 11061 18522
rect 11085 18470 11095 18522
rect 11095 18470 11141 18522
rect 10845 18468 10901 18470
rect 10925 18468 10981 18470
rect 11005 18468 11061 18470
rect 11085 18468 11141 18470
rect 8373 17978 8429 17980
rect 8453 17978 8509 17980
rect 8533 17978 8589 17980
rect 8613 17978 8669 17980
rect 8373 17926 8419 17978
rect 8419 17926 8429 17978
rect 8453 17926 8483 17978
rect 8483 17926 8495 17978
rect 8495 17926 8509 17978
rect 8533 17926 8547 17978
rect 8547 17926 8559 17978
rect 8559 17926 8589 17978
rect 8613 17926 8623 17978
rect 8623 17926 8669 17978
rect 8373 17924 8429 17926
rect 8453 17924 8509 17926
rect 8533 17924 8589 17926
rect 8613 17924 8669 17926
rect 5900 17434 5956 17436
rect 5980 17434 6036 17436
rect 6060 17434 6116 17436
rect 6140 17434 6196 17436
rect 5900 17382 5946 17434
rect 5946 17382 5956 17434
rect 5980 17382 6010 17434
rect 6010 17382 6022 17434
rect 6022 17382 6036 17434
rect 6060 17382 6074 17434
rect 6074 17382 6086 17434
rect 6086 17382 6116 17434
rect 6140 17382 6150 17434
rect 6150 17382 6196 17434
rect 5900 17380 5956 17382
rect 5980 17380 6036 17382
rect 6060 17380 6116 17382
rect 6140 17380 6196 17382
rect 3428 14714 3484 14716
rect 3508 14714 3564 14716
rect 3588 14714 3644 14716
rect 3668 14714 3724 14716
rect 3428 14662 3474 14714
rect 3474 14662 3484 14714
rect 3508 14662 3538 14714
rect 3538 14662 3550 14714
rect 3550 14662 3564 14714
rect 3588 14662 3602 14714
rect 3602 14662 3614 14714
rect 3614 14662 3644 14714
rect 3668 14662 3678 14714
rect 3678 14662 3724 14714
rect 3428 14660 3484 14662
rect 3508 14660 3564 14662
rect 3588 14660 3644 14662
rect 3668 14660 3724 14662
rect 3428 13626 3484 13628
rect 3508 13626 3564 13628
rect 3588 13626 3644 13628
rect 3668 13626 3724 13628
rect 3428 13574 3474 13626
rect 3474 13574 3484 13626
rect 3508 13574 3538 13626
rect 3538 13574 3550 13626
rect 3550 13574 3564 13626
rect 3588 13574 3602 13626
rect 3602 13574 3614 13626
rect 3614 13574 3644 13626
rect 3668 13574 3678 13626
rect 3678 13574 3724 13626
rect 3428 13572 3484 13574
rect 3508 13572 3564 13574
rect 3588 13572 3644 13574
rect 3668 13572 3724 13574
rect 10845 17434 10901 17436
rect 10925 17434 10981 17436
rect 11005 17434 11061 17436
rect 11085 17434 11141 17436
rect 10845 17382 10891 17434
rect 10891 17382 10901 17434
rect 10925 17382 10955 17434
rect 10955 17382 10967 17434
rect 10967 17382 10981 17434
rect 11005 17382 11019 17434
rect 11019 17382 11031 17434
rect 11031 17382 11061 17434
rect 11085 17382 11095 17434
rect 11095 17382 11141 17434
rect 10845 17380 10901 17382
rect 10925 17380 10981 17382
rect 11005 17380 11061 17382
rect 11085 17380 11141 17382
rect 8373 16890 8429 16892
rect 8453 16890 8509 16892
rect 8533 16890 8589 16892
rect 8613 16890 8669 16892
rect 8373 16838 8419 16890
rect 8419 16838 8429 16890
rect 8453 16838 8483 16890
rect 8483 16838 8495 16890
rect 8495 16838 8509 16890
rect 8533 16838 8547 16890
rect 8547 16838 8559 16890
rect 8559 16838 8589 16890
rect 8613 16838 8623 16890
rect 8623 16838 8669 16890
rect 8373 16836 8429 16838
rect 8453 16836 8509 16838
rect 8533 16836 8589 16838
rect 8613 16836 8669 16838
rect 5900 16346 5956 16348
rect 5980 16346 6036 16348
rect 6060 16346 6116 16348
rect 6140 16346 6196 16348
rect 5900 16294 5946 16346
rect 5946 16294 5956 16346
rect 5980 16294 6010 16346
rect 6010 16294 6022 16346
rect 6022 16294 6036 16346
rect 6060 16294 6074 16346
rect 6074 16294 6086 16346
rect 6086 16294 6116 16346
rect 6140 16294 6150 16346
rect 6150 16294 6196 16346
rect 5900 16292 5956 16294
rect 5980 16292 6036 16294
rect 6060 16292 6116 16294
rect 6140 16292 6196 16294
rect 13318 17978 13374 17980
rect 13398 17978 13454 17980
rect 13478 17978 13534 17980
rect 13558 17978 13614 17980
rect 13318 17926 13364 17978
rect 13364 17926 13374 17978
rect 13398 17926 13428 17978
rect 13428 17926 13440 17978
rect 13440 17926 13454 17978
rect 13478 17926 13492 17978
rect 13492 17926 13504 17978
rect 13504 17926 13534 17978
rect 13558 17926 13568 17978
rect 13568 17926 13614 17978
rect 13318 17924 13374 17926
rect 13398 17924 13454 17926
rect 13478 17924 13534 17926
rect 13558 17924 13614 17926
rect 15790 19610 15846 19612
rect 15870 19610 15926 19612
rect 15950 19610 16006 19612
rect 16030 19610 16086 19612
rect 15790 19558 15836 19610
rect 15836 19558 15846 19610
rect 15870 19558 15900 19610
rect 15900 19558 15912 19610
rect 15912 19558 15926 19610
rect 15950 19558 15964 19610
rect 15964 19558 15976 19610
rect 15976 19558 16006 19610
rect 16030 19558 16040 19610
rect 16040 19558 16086 19610
rect 15790 19556 15846 19558
rect 15870 19556 15926 19558
rect 15950 19556 16006 19558
rect 16030 19556 16086 19558
rect 20735 19610 20791 19612
rect 20815 19610 20871 19612
rect 20895 19610 20951 19612
rect 20975 19610 21031 19612
rect 20735 19558 20781 19610
rect 20781 19558 20791 19610
rect 20815 19558 20845 19610
rect 20845 19558 20857 19610
rect 20857 19558 20871 19610
rect 20895 19558 20909 19610
rect 20909 19558 20921 19610
rect 20921 19558 20951 19610
rect 20975 19558 20985 19610
rect 20985 19558 21031 19610
rect 20735 19556 20791 19558
rect 20815 19556 20871 19558
rect 20895 19556 20951 19558
rect 20975 19556 21031 19558
rect 15198 18264 15254 18320
rect 10506 16632 10562 16688
rect 8373 15802 8429 15804
rect 8453 15802 8509 15804
rect 8533 15802 8589 15804
rect 8613 15802 8669 15804
rect 8373 15750 8419 15802
rect 8419 15750 8429 15802
rect 8453 15750 8483 15802
rect 8483 15750 8495 15802
rect 8495 15750 8509 15802
rect 8533 15750 8547 15802
rect 8547 15750 8559 15802
rect 8559 15750 8589 15802
rect 8613 15750 8623 15802
rect 8623 15750 8669 15802
rect 8373 15748 8429 15750
rect 8453 15748 8509 15750
rect 8533 15748 8589 15750
rect 8613 15748 8669 15750
rect 5900 15258 5956 15260
rect 5980 15258 6036 15260
rect 6060 15258 6116 15260
rect 6140 15258 6196 15260
rect 5900 15206 5946 15258
rect 5946 15206 5956 15258
rect 5980 15206 6010 15258
rect 6010 15206 6022 15258
rect 6022 15206 6036 15258
rect 6060 15206 6074 15258
rect 6074 15206 6086 15258
rect 6086 15206 6116 15258
rect 6140 15206 6150 15258
rect 6150 15206 6196 15258
rect 5900 15204 5956 15206
rect 5980 15204 6036 15206
rect 6060 15204 6116 15206
rect 6140 15204 6196 15206
rect 8373 14714 8429 14716
rect 8453 14714 8509 14716
rect 8533 14714 8589 14716
rect 8613 14714 8669 14716
rect 8373 14662 8419 14714
rect 8419 14662 8429 14714
rect 8453 14662 8483 14714
rect 8483 14662 8495 14714
rect 8495 14662 8509 14714
rect 8533 14662 8547 14714
rect 8547 14662 8559 14714
rect 8559 14662 8589 14714
rect 8613 14662 8623 14714
rect 8623 14662 8669 14714
rect 8373 14660 8429 14662
rect 8453 14660 8509 14662
rect 8533 14660 8589 14662
rect 8613 14660 8669 14662
rect 5900 14170 5956 14172
rect 5980 14170 6036 14172
rect 6060 14170 6116 14172
rect 6140 14170 6196 14172
rect 5900 14118 5946 14170
rect 5946 14118 5956 14170
rect 5980 14118 6010 14170
rect 6010 14118 6022 14170
rect 6022 14118 6036 14170
rect 6060 14118 6074 14170
rect 6074 14118 6086 14170
rect 6086 14118 6116 14170
rect 6140 14118 6150 14170
rect 6150 14118 6196 14170
rect 5900 14116 5956 14118
rect 5980 14116 6036 14118
rect 6060 14116 6116 14118
rect 6140 14116 6196 14118
rect 5900 13082 5956 13084
rect 5980 13082 6036 13084
rect 6060 13082 6116 13084
rect 6140 13082 6196 13084
rect 5900 13030 5946 13082
rect 5946 13030 5956 13082
rect 5980 13030 6010 13082
rect 6010 13030 6022 13082
rect 6022 13030 6036 13082
rect 6060 13030 6074 13082
rect 6074 13030 6086 13082
rect 6086 13030 6116 13082
rect 6140 13030 6150 13082
rect 6150 13030 6196 13082
rect 5900 13028 5956 13030
rect 5980 13028 6036 13030
rect 6060 13028 6116 13030
rect 6140 13028 6196 13030
rect 3428 12538 3484 12540
rect 3508 12538 3564 12540
rect 3588 12538 3644 12540
rect 3668 12538 3724 12540
rect 3428 12486 3474 12538
rect 3474 12486 3484 12538
rect 3508 12486 3538 12538
rect 3538 12486 3550 12538
rect 3550 12486 3564 12538
rect 3588 12486 3602 12538
rect 3602 12486 3614 12538
rect 3614 12486 3644 12538
rect 3668 12486 3678 12538
rect 3678 12486 3724 12538
rect 3428 12484 3484 12486
rect 3508 12484 3564 12486
rect 3588 12484 3644 12486
rect 3668 12484 3724 12486
rect 3428 11450 3484 11452
rect 3508 11450 3564 11452
rect 3588 11450 3644 11452
rect 3668 11450 3724 11452
rect 3428 11398 3474 11450
rect 3474 11398 3484 11450
rect 3508 11398 3538 11450
rect 3538 11398 3550 11450
rect 3550 11398 3564 11450
rect 3588 11398 3602 11450
rect 3602 11398 3614 11450
rect 3614 11398 3644 11450
rect 3668 11398 3678 11450
rect 3678 11398 3724 11450
rect 3428 11396 3484 11398
rect 3508 11396 3564 11398
rect 3588 11396 3644 11398
rect 3668 11396 3724 11398
rect 3428 10362 3484 10364
rect 3508 10362 3564 10364
rect 3588 10362 3644 10364
rect 3668 10362 3724 10364
rect 3428 10310 3474 10362
rect 3474 10310 3484 10362
rect 3508 10310 3538 10362
rect 3538 10310 3550 10362
rect 3550 10310 3564 10362
rect 3588 10310 3602 10362
rect 3602 10310 3614 10362
rect 3614 10310 3644 10362
rect 3668 10310 3678 10362
rect 3678 10310 3724 10362
rect 3428 10308 3484 10310
rect 3508 10308 3564 10310
rect 3588 10308 3644 10310
rect 3668 10308 3724 10310
rect 3428 9274 3484 9276
rect 3508 9274 3564 9276
rect 3588 9274 3644 9276
rect 3668 9274 3724 9276
rect 3428 9222 3474 9274
rect 3474 9222 3484 9274
rect 3508 9222 3538 9274
rect 3538 9222 3550 9274
rect 3550 9222 3564 9274
rect 3588 9222 3602 9274
rect 3602 9222 3614 9274
rect 3614 9222 3644 9274
rect 3668 9222 3678 9274
rect 3678 9222 3724 9274
rect 3428 9220 3484 9222
rect 3508 9220 3564 9222
rect 3588 9220 3644 9222
rect 3668 9220 3724 9222
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3588 8186 3644 8188
rect 3668 8186 3724 8188
rect 3428 8134 3474 8186
rect 3474 8134 3484 8186
rect 3508 8134 3538 8186
rect 3538 8134 3550 8186
rect 3550 8134 3564 8186
rect 3588 8134 3602 8186
rect 3602 8134 3614 8186
rect 3614 8134 3644 8186
rect 3668 8134 3678 8186
rect 3678 8134 3724 8186
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 3588 8132 3644 8134
rect 3668 8132 3724 8134
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3588 7098 3644 7100
rect 3668 7098 3724 7100
rect 3428 7046 3474 7098
rect 3474 7046 3484 7098
rect 3508 7046 3538 7098
rect 3538 7046 3550 7098
rect 3550 7046 3564 7098
rect 3588 7046 3602 7098
rect 3602 7046 3614 7098
rect 3614 7046 3644 7098
rect 3668 7046 3678 7098
rect 3678 7046 3724 7098
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 3588 7044 3644 7046
rect 3668 7044 3724 7046
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3588 6010 3644 6012
rect 3668 6010 3724 6012
rect 3428 5958 3474 6010
rect 3474 5958 3484 6010
rect 3508 5958 3538 6010
rect 3538 5958 3550 6010
rect 3550 5958 3564 6010
rect 3588 5958 3602 6010
rect 3602 5958 3614 6010
rect 3614 5958 3644 6010
rect 3668 5958 3678 6010
rect 3678 5958 3724 6010
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 3588 5956 3644 5958
rect 3668 5956 3724 5958
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3588 4922 3644 4924
rect 3668 4922 3724 4924
rect 3428 4870 3474 4922
rect 3474 4870 3484 4922
rect 3508 4870 3538 4922
rect 3538 4870 3550 4922
rect 3550 4870 3564 4922
rect 3588 4870 3602 4922
rect 3602 4870 3614 4922
rect 3614 4870 3644 4922
rect 3668 4870 3678 4922
rect 3678 4870 3724 4922
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 3588 4868 3644 4870
rect 3668 4868 3724 4870
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3588 3834 3644 3836
rect 3668 3834 3724 3836
rect 3428 3782 3474 3834
rect 3474 3782 3484 3834
rect 3508 3782 3538 3834
rect 3538 3782 3550 3834
rect 3550 3782 3564 3834
rect 3588 3782 3602 3834
rect 3602 3782 3614 3834
rect 3614 3782 3644 3834
rect 3668 3782 3678 3834
rect 3678 3782 3724 3834
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 3588 3780 3644 3782
rect 3668 3780 3724 3782
rect 5900 11994 5956 11996
rect 5980 11994 6036 11996
rect 6060 11994 6116 11996
rect 6140 11994 6196 11996
rect 5900 11942 5946 11994
rect 5946 11942 5956 11994
rect 5980 11942 6010 11994
rect 6010 11942 6022 11994
rect 6022 11942 6036 11994
rect 6060 11942 6074 11994
rect 6074 11942 6086 11994
rect 6086 11942 6116 11994
rect 6140 11942 6150 11994
rect 6150 11942 6196 11994
rect 5900 11940 5956 11942
rect 5980 11940 6036 11942
rect 6060 11940 6116 11942
rect 6140 11940 6196 11942
rect 5900 10906 5956 10908
rect 5980 10906 6036 10908
rect 6060 10906 6116 10908
rect 6140 10906 6196 10908
rect 5900 10854 5946 10906
rect 5946 10854 5956 10906
rect 5980 10854 6010 10906
rect 6010 10854 6022 10906
rect 6022 10854 6036 10906
rect 6060 10854 6074 10906
rect 6074 10854 6086 10906
rect 6086 10854 6116 10906
rect 6140 10854 6150 10906
rect 6150 10854 6196 10906
rect 5900 10852 5956 10854
rect 5980 10852 6036 10854
rect 6060 10852 6116 10854
rect 6140 10852 6196 10854
rect 5900 9818 5956 9820
rect 5980 9818 6036 9820
rect 6060 9818 6116 9820
rect 6140 9818 6196 9820
rect 5900 9766 5946 9818
rect 5946 9766 5956 9818
rect 5980 9766 6010 9818
rect 6010 9766 6022 9818
rect 6022 9766 6036 9818
rect 6060 9766 6074 9818
rect 6074 9766 6086 9818
rect 6086 9766 6116 9818
rect 6140 9766 6150 9818
rect 6150 9766 6196 9818
rect 5900 9764 5956 9766
rect 5980 9764 6036 9766
rect 6060 9764 6116 9766
rect 6140 9764 6196 9766
rect 5900 8730 5956 8732
rect 5980 8730 6036 8732
rect 6060 8730 6116 8732
rect 6140 8730 6196 8732
rect 5900 8678 5946 8730
rect 5946 8678 5956 8730
rect 5980 8678 6010 8730
rect 6010 8678 6022 8730
rect 6022 8678 6036 8730
rect 6060 8678 6074 8730
rect 6074 8678 6086 8730
rect 6086 8678 6116 8730
rect 6140 8678 6150 8730
rect 6150 8678 6196 8730
rect 5900 8676 5956 8678
rect 5980 8676 6036 8678
rect 6060 8676 6116 8678
rect 6140 8676 6196 8678
rect 5900 7642 5956 7644
rect 5980 7642 6036 7644
rect 6060 7642 6116 7644
rect 6140 7642 6196 7644
rect 5900 7590 5946 7642
rect 5946 7590 5956 7642
rect 5980 7590 6010 7642
rect 6010 7590 6022 7642
rect 6022 7590 6036 7642
rect 6060 7590 6074 7642
rect 6074 7590 6086 7642
rect 6086 7590 6116 7642
rect 6140 7590 6150 7642
rect 6150 7590 6196 7642
rect 5900 7588 5956 7590
rect 5980 7588 6036 7590
rect 6060 7588 6116 7590
rect 6140 7588 6196 7590
rect 5900 6554 5956 6556
rect 5980 6554 6036 6556
rect 6060 6554 6116 6556
rect 6140 6554 6196 6556
rect 5900 6502 5946 6554
rect 5946 6502 5956 6554
rect 5980 6502 6010 6554
rect 6010 6502 6022 6554
rect 6022 6502 6036 6554
rect 6060 6502 6074 6554
rect 6074 6502 6086 6554
rect 6086 6502 6116 6554
rect 6140 6502 6150 6554
rect 6150 6502 6196 6554
rect 5900 6500 5956 6502
rect 5980 6500 6036 6502
rect 6060 6500 6116 6502
rect 6140 6500 6196 6502
rect 5900 5466 5956 5468
rect 5980 5466 6036 5468
rect 6060 5466 6116 5468
rect 6140 5466 6196 5468
rect 5900 5414 5946 5466
rect 5946 5414 5956 5466
rect 5980 5414 6010 5466
rect 6010 5414 6022 5466
rect 6022 5414 6036 5466
rect 6060 5414 6074 5466
rect 6074 5414 6086 5466
rect 6086 5414 6116 5466
rect 6140 5414 6150 5466
rect 6150 5414 6196 5466
rect 5900 5412 5956 5414
rect 5980 5412 6036 5414
rect 6060 5412 6116 5414
rect 6140 5412 6196 5414
rect 5900 4378 5956 4380
rect 5980 4378 6036 4380
rect 6060 4378 6116 4380
rect 6140 4378 6196 4380
rect 5900 4326 5946 4378
rect 5946 4326 5956 4378
rect 5980 4326 6010 4378
rect 6010 4326 6022 4378
rect 6022 4326 6036 4378
rect 6060 4326 6074 4378
rect 6074 4326 6086 4378
rect 6086 4326 6116 4378
rect 6140 4326 6150 4378
rect 6150 4326 6196 4378
rect 5900 4324 5956 4326
rect 5980 4324 6036 4326
rect 6060 4324 6116 4326
rect 6140 4324 6196 4326
rect 5900 3290 5956 3292
rect 5980 3290 6036 3292
rect 6060 3290 6116 3292
rect 6140 3290 6196 3292
rect 5900 3238 5946 3290
rect 5946 3238 5956 3290
rect 5980 3238 6010 3290
rect 6010 3238 6022 3290
rect 6022 3238 6036 3290
rect 6060 3238 6074 3290
rect 6074 3238 6086 3290
rect 6086 3238 6116 3290
rect 6140 3238 6150 3290
rect 6150 3238 6196 3290
rect 5900 3236 5956 3238
rect 5980 3236 6036 3238
rect 6060 3236 6116 3238
rect 6140 3236 6196 3238
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3588 2746 3644 2748
rect 3668 2746 3724 2748
rect 3428 2694 3474 2746
rect 3474 2694 3484 2746
rect 3508 2694 3538 2746
rect 3538 2694 3550 2746
rect 3550 2694 3564 2746
rect 3588 2694 3602 2746
rect 3602 2694 3614 2746
rect 3614 2694 3644 2746
rect 3668 2694 3678 2746
rect 3678 2694 3724 2746
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 3588 2692 3644 2694
rect 3668 2692 3724 2694
rect 8373 13626 8429 13628
rect 8453 13626 8509 13628
rect 8533 13626 8589 13628
rect 8613 13626 8669 13628
rect 8373 13574 8419 13626
rect 8419 13574 8429 13626
rect 8453 13574 8483 13626
rect 8483 13574 8495 13626
rect 8495 13574 8509 13626
rect 8533 13574 8547 13626
rect 8547 13574 8559 13626
rect 8559 13574 8589 13626
rect 8613 13574 8623 13626
rect 8623 13574 8669 13626
rect 8373 13572 8429 13574
rect 8453 13572 8509 13574
rect 8533 13572 8589 13574
rect 8613 13572 8669 13574
rect 8373 12538 8429 12540
rect 8453 12538 8509 12540
rect 8533 12538 8589 12540
rect 8613 12538 8669 12540
rect 8373 12486 8419 12538
rect 8419 12486 8429 12538
rect 8453 12486 8483 12538
rect 8483 12486 8495 12538
rect 8495 12486 8509 12538
rect 8533 12486 8547 12538
rect 8547 12486 8559 12538
rect 8559 12486 8589 12538
rect 8613 12486 8623 12538
rect 8623 12486 8669 12538
rect 8373 12484 8429 12486
rect 8453 12484 8509 12486
rect 8533 12484 8589 12486
rect 8613 12484 8669 12486
rect 8373 11450 8429 11452
rect 8453 11450 8509 11452
rect 8533 11450 8589 11452
rect 8613 11450 8669 11452
rect 8373 11398 8419 11450
rect 8419 11398 8429 11450
rect 8453 11398 8483 11450
rect 8483 11398 8495 11450
rect 8495 11398 8509 11450
rect 8533 11398 8547 11450
rect 8547 11398 8559 11450
rect 8559 11398 8589 11450
rect 8613 11398 8623 11450
rect 8623 11398 8669 11450
rect 8373 11396 8429 11398
rect 8453 11396 8509 11398
rect 8533 11396 8589 11398
rect 8613 11396 8669 11398
rect 8373 10362 8429 10364
rect 8453 10362 8509 10364
rect 8533 10362 8589 10364
rect 8613 10362 8669 10364
rect 8373 10310 8419 10362
rect 8419 10310 8429 10362
rect 8453 10310 8483 10362
rect 8483 10310 8495 10362
rect 8495 10310 8509 10362
rect 8533 10310 8547 10362
rect 8547 10310 8559 10362
rect 8559 10310 8589 10362
rect 8613 10310 8623 10362
rect 8623 10310 8669 10362
rect 8373 10308 8429 10310
rect 8453 10308 8509 10310
rect 8533 10308 8589 10310
rect 8613 10308 8669 10310
rect 8373 9274 8429 9276
rect 8453 9274 8509 9276
rect 8533 9274 8589 9276
rect 8613 9274 8669 9276
rect 8373 9222 8419 9274
rect 8419 9222 8429 9274
rect 8453 9222 8483 9274
rect 8483 9222 8495 9274
rect 8495 9222 8509 9274
rect 8533 9222 8547 9274
rect 8547 9222 8559 9274
rect 8559 9222 8589 9274
rect 8613 9222 8623 9274
rect 8623 9222 8669 9274
rect 8373 9220 8429 9222
rect 8453 9220 8509 9222
rect 8533 9220 8589 9222
rect 8613 9220 8669 9222
rect 8373 8186 8429 8188
rect 8453 8186 8509 8188
rect 8533 8186 8589 8188
rect 8613 8186 8669 8188
rect 8373 8134 8419 8186
rect 8419 8134 8429 8186
rect 8453 8134 8483 8186
rect 8483 8134 8495 8186
rect 8495 8134 8509 8186
rect 8533 8134 8547 8186
rect 8547 8134 8559 8186
rect 8559 8134 8589 8186
rect 8613 8134 8623 8186
rect 8623 8134 8669 8186
rect 8373 8132 8429 8134
rect 8453 8132 8509 8134
rect 8533 8132 8589 8134
rect 8613 8132 8669 8134
rect 8373 7098 8429 7100
rect 8453 7098 8509 7100
rect 8533 7098 8589 7100
rect 8613 7098 8669 7100
rect 8373 7046 8419 7098
rect 8419 7046 8429 7098
rect 8453 7046 8483 7098
rect 8483 7046 8495 7098
rect 8495 7046 8509 7098
rect 8533 7046 8547 7098
rect 8547 7046 8559 7098
rect 8559 7046 8589 7098
rect 8613 7046 8623 7098
rect 8623 7046 8669 7098
rect 8373 7044 8429 7046
rect 8453 7044 8509 7046
rect 8533 7044 8589 7046
rect 8613 7044 8669 7046
rect 8373 6010 8429 6012
rect 8453 6010 8509 6012
rect 8533 6010 8589 6012
rect 8613 6010 8669 6012
rect 8373 5958 8419 6010
rect 8419 5958 8429 6010
rect 8453 5958 8483 6010
rect 8483 5958 8495 6010
rect 8495 5958 8509 6010
rect 8533 5958 8547 6010
rect 8547 5958 8559 6010
rect 8559 5958 8589 6010
rect 8613 5958 8623 6010
rect 8623 5958 8669 6010
rect 8373 5956 8429 5958
rect 8453 5956 8509 5958
rect 8533 5956 8589 5958
rect 8613 5956 8669 5958
rect 8373 4922 8429 4924
rect 8453 4922 8509 4924
rect 8533 4922 8589 4924
rect 8613 4922 8669 4924
rect 8373 4870 8419 4922
rect 8419 4870 8429 4922
rect 8453 4870 8483 4922
rect 8483 4870 8495 4922
rect 8495 4870 8509 4922
rect 8533 4870 8547 4922
rect 8547 4870 8559 4922
rect 8559 4870 8589 4922
rect 8613 4870 8623 4922
rect 8623 4870 8669 4922
rect 8373 4868 8429 4870
rect 8453 4868 8509 4870
rect 8533 4868 8589 4870
rect 8613 4868 8669 4870
rect 8373 3834 8429 3836
rect 8453 3834 8509 3836
rect 8533 3834 8589 3836
rect 8613 3834 8669 3836
rect 8373 3782 8419 3834
rect 8419 3782 8429 3834
rect 8453 3782 8483 3834
rect 8483 3782 8495 3834
rect 8495 3782 8509 3834
rect 8533 3782 8547 3834
rect 8547 3782 8559 3834
rect 8559 3782 8589 3834
rect 8613 3782 8623 3834
rect 8623 3782 8669 3834
rect 8373 3780 8429 3782
rect 8453 3780 8509 3782
rect 8533 3780 8589 3782
rect 8613 3780 8669 3782
rect 8373 2746 8429 2748
rect 8453 2746 8509 2748
rect 8533 2746 8589 2748
rect 8613 2746 8669 2748
rect 8373 2694 8419 2746
rect 8419 2694 8429 2746
rect 8453 2694 8483 2746
rect 8483 2694 8495 2746
rect 8495 2694 8509 2746
rect 8533 2694 8547 2746
rect 8547 2694 8559 2746
rect 8559 2694 8589 2746
rect 8613 2694 8623 2746
rect 8623 2694 8669 2746
rect 8373 2692 8429 2694
rect 8453 2692 8509 2694
rect 8533 2692 8589 2694
rect 8613 2692 8669 2694
rect 13318 16890 13374 16892
rect 13398 16890 13454 16892
rect 13478 16890 13534 16892
rect 13558 16890 13614 16892
rect 13318 16838 13364 16890
rect 13364 16838 13374 16890
rect 13398 16838 13428 16890
rect 13428 16838 13440 16890
rect 13440 16838 13454 16890
rect 13478 16838 13492 16890
rect 13492 16838 13504 16890
rect 13504 16838 13534 16890
rect 13558 16838 13568 16890
rect 13568 16838 13614 16890
rect 13318 16836 13374 16838
rect 13398 16836 13454 16838
rect 13478 16836 13534 16838
rect 13558 16836 13614 16838
rect 10845 16346 10901 16348
rect 10925 16346 10981 16348
rect 11005 16346 11061 16348
rect 11085 16346 11141 16348
rect 10845 16294 10891 16346
rect 10891 16294 10901 16346
rect 10925 16294 10955 16346
rect 10955 16294 10967 16346
rect 10967 16294 10981 16346
rect 11005 16294 11019 16346
rect 11019 16294 11031 16346
rect 11031 16294 11061 16346
rect 11085 16294 11095 16346
rect 11095 16294 11141 16346
rect 10845 16292 10901 16294
rect 10925 16292 10981 16294
rect 11005 16292 11061 16294
rect 11085 16292 11141 16294
rect 10845 15258 10901 15260
rect 10925 15258 10981 15260
rect 11005 15258 11061 15260
rect 11085 15258 11141 15260
rect 10845 15206 10891 15258
rect 10891 15206 10901 15258
rect 10925 15206 10955 15258
rect 10955 15206 10967 15258
rect 10967 15206 10981 15258
rect 11005 15206 11019 15258
rect 11019 15206 11031 15258
rect 11031 15206 11061 15258
rect 11085 15206 11095 15258
rect 11095 15206 11141 15258
rect 10845 15204 10901 15206
rect 10925 15204 10981 15206
rect 11005 15204 11061 15206
rect 11085 15204 11141 15206
rect 10845 14170 10901 14172
rect 10925 14170 10981 14172
rect 11005 14170 11061 14172
rect 11085 14170 11141 14172
rect 10845 14118 10891 14170
rect 10891 14118 10901 14170
rect 10925 14118 10955 14170
rect 10955 14118 10967 14170
rect 10967 14118 10981 14170
rect 11005 14118 11019 14170
rect 11019 14118 11031 14170
rect 11031 14118 11061 14170
rect 11085 14118 11095 14170
rect 11095 14118 11141 14170
rect 10845 14116 10901 14118
rect 10925 14116 10981 14118
rect 11005 14116 11061 14118
rect 11085 14116 11141 14118
rect 10845 13082 10901 13084
rect 10925 13082 10981 13084
rect 11005 13082 11061 13084
rect 11085 13082 11141 13084
rect 10845 13030 10891 13082
rect 10891 13030 10901 13082
rect 10925 13030 10955 13082
rect 10955 13030 10967 13082
rect 10967 13030 10981 13082
rect 11005 13030 11019 13082
rect 11019 13030 11031 13082
rect 11031 13030 11061 13082
rect 11085 13030 11095 13082
rect 11095 13030 11141 13082
rect 10845 13028 10901 13030
rect 10925 13028 10981 13030
rect 11005 13028 11061 13030
rect 11085 13028 11141 13030
rect 10230 6316 10286 6352
rect 10230 6296 10232 6316
rect 10232 6296 10284 6316
rect 10284 6296 10286 6316
rect 10845 11994 10901 11996
rect 10925 11994 10981 11996
rect 11005 11994 11061 11996
rect 11085 11994 11141 11996
rect 10845 11942 10891 11994
rect 10891 11942 10901 11994
rect 10925 11942 10955 11994
rect 10955 11942 10967 11994
rect 10967 11942 10981 11994
rect 11005 11942 11019 11994
rect 11019 11942 11031 11994
rect 11031 11942 11061 11994
rect 11085 11942 11095 11994
rect 11095 11942 11141 11994
rect 10845 11940 10901 11942
rect 10925 11940 10981 11942
rect 11005 11940 11061 11942
rect 11085 11940 11141 11942
rect 10845 10906 10901 10908
rect 10925 10906 10981 10908
rect 11005 10906 11061 10908
rect 11085 10906 11141 10908
rect 10845 10854 10891 10906
rect 10891 10854 10901 10906
rect 10925 10854 10955 10906
rect 10955 10854 10967 10906
rect 10967 10854 10981 10906
rect 11005 10854 11019 10906
rect 11019 10854 11031 10906
rect 11031 10854 11061 10906
rect 11085 10854 11095 10906
rect 11095 10854 11141 10906
rect 10845 10852 10901 10854
rect 10925 10852 10981 10854
rect 11005 10852 11061 10854
rect 11085 10852 11141 10854
rect 10845 9818 10901 9820
rect 10925 9818 10981 9820
rect 11005 9818 11061 9820
rect 11085 9818 11141 9820
rect 10845 9766 10891 9818
rect 10891 9766 10901 9818
rect 10925 9766 10955 9818
rect 10955 9766 10967 9818
rect 10967 9766 10981 9818
rect 11005 9766 11019 9818
rect 11019 9766 11031 9818
rect 11031 9766 11061 9818
rect 11085 9766 11095 9818
rect 11095 9766 11141 9818
rect 10845 9764 10901 9766
rect 10925 9764 10981 9766
rect 11005 9764 11061 9766
rect 11085 9764 11141 9766
rect 10845 8730 10901 8732
rect 10925 8730 10981 8732
rect 11005 8730 11061 8732
rect 11085 8730 11141 8732
rect 10845 8678 10891 8730
rect 10891 8678 10901 8730
rect 10925 8678 10955 8730
rect 10955 8678 10967 8730
rect 10967 8678 10981 8730
rect 11005 8678 11019 8730
rect 11019 8678 11031 8730
rect 11031 8678 11061 8730
rect 11085 8678 11095 8730
rect 11095 8678 11141 8730
rect 10845 8676 10901 8678
rect 10925 8676 10981 8678
rect 11005 8676 11061 8678
rect 11085 8676 11141 8678
rect 13318 15802 13374 15804
rect 13398 15802 13454 15804
rect 13478 15802 13534 15804
rect 13558 15802 13614 15804
rect 13318 15750 13364 15802
rect 13364 15750 13374 15802
rect 13398 15750 13428 15802
rect 13428 15750 13440 15802
rect 13440 15750 13454 15802
rect 13478 15750 13492 15802
rect 13492 15750 13504 15802
rect 13504 15750 13534 15802
rect 13558 15750 13568 15802
rect 13568 15750 13614 15802
rect 13318 15748 13374 15750
rect 13398 15748 13454 15750
rect 13478 15748 13534 15750
rect 13558 15748 13614 15750
rect 13318 14714 13374 14716
rect 13398 14714 13454 14716
rect 13478 14714 13534 14716
rect 13558 14714 13614 14716
rect 13318 14662 13364 14714
rect 13364 14662 13374 14714
rect 13398 14662 13428 14714
rect 13428 14662 13440 14714
rect 13440 14662 13454 14714
rect 13478 14662 13492 14714
rect 13492 14662 13504 14714
rect 13504 14662 13534 14714
rect 13558 14662 13568 14714
rect 13568 14662 13614 14714
rect 13318 14660 13374 14662
rect 13398 14660 13454 14662
rect 13478 14660 13534 14662
rect 13558 14660 13614 14662
rect 13318 13626 13374 13628
rect 13398 13626 13454 13628
rect 13478 13626 13534 13628
rect 13558 13626 13614 13628
rect 13318 13574 13364 13626
rect 13364 13574 13374 13626
rect 13398 13574 13428 13626
rect 13428 13574 13440 13626
rect 13440 13574 13454 13626
rect 13478 13574 13492 13626
rect 13492 13574 13504 13626
rect 13504 13574 13534 13626
rect 13558 13574 13568 13626
rect 13568 13574 13614 13626
rect 13318 13572 13374 13574
rect 13398 13572 13454 13574
rect 13478 13572 13534 13574
rect 13558 13572 13614 13574
rect 13318 12538 13374 12540
rect 13398 12538 13454 12540
rect 13478 12538 13534 12540
rect 13558 12538 13614 12540
rect 13318 12486 13364 12538
rect 13364 12486 13374 12538
rect 13398 12486 13428 12538
rect 13428 12486 13440 12538
rect 13440 12486 13454 12538
rect 13478 12486 13492 12538
rect 13492 12486 13504 12538
rect 13504 12486 13534 12538
rect 13558 12486 13568 12538
rect 13568 12486 13614 12538
rect 13318 12484 13374 12486
rect 13398 12484 13454 12486
rect 13478 12484 13534 12486
rect 13558 12484 13614 12486
rect 13318 11450 13374 11452
rect 13398 11450 13454 11452
rect 13478 11450 13534 11452
rect 13558 11450 13614 11452
rect 13318 11398 13364 11450
rect 13364 11398 13374 11450
rect 13398 11398 13428 11450
rect 13428 11398 13440 11450
rect 13440 11398 13454 11450
rect 13478 11398 13492 11450
rect 13492 11398 13504 11450
rect 13504 11398 13534 11450
rect 13558 11398 13568 11450
rect 13568 11398 13614 11450
rect 13318 11396 13374 11398
rect 13398 11396 13454 11398
rect 13478 11396 13534 11398
rect 13558 11396 13614 11398
rect 10845 7642 10901 7644
rect 10925 7642 10981 7644
rect 11005 7642 11061 7644
rect 11085 7642 11141 7644
rect 10845 7590 10891 7642
rect 10891 7590 10901 7642
rect 10925 7590 10955 7642
rect 10955 7590 10967 7642
rect 10967 7590 10981 7642
rect 11005 7590 11019 7642
rect 11019 7590 11031 7642
rect 11031 7590 11061 7642
rect 11085 7590 11095 7642
rect 11095 7590 11141 7642
rect 10845 7588 10901 7590
rect 10925 7588 10981 7590
rect 11005 7588 11061 7590
rect 11085 7588 11141 7590
rect 10845 6554 10901 6556
rect 10925 6554 10981 6556
rect 11005 6554 11061 6556
rect 11085 6554 11141 6556
rect 10845 6502 10891 6554
rect 10891 6502 10901 6554
rect 10925 6502 10955 6554
rect 10955 6502 10967 6554
rect 10967 6502 10981 6554
rect 11005 6502 11019 6554
rect 11019 6502 11031 6554
rect 11031 6502 11061 6554
rect 11085 6502 11095 6554
rect 11095 6502 11141 6554
rect 10845 6500 10901 6502
rect 10925 6500 10981 6502
rect 11005 6500 11061 6502
rect 11085 6500 11141 6502
rect 10845 5466 10901 5468
rect 10925 5466 10981 5468
rect 11005 5466 11061 5468
rect 11085 5466 11141 5468
rect 10845 5414 10891 5466
rect 10891 5414 10901 5466
rect 10925 5414 10955 5466
rect 10955 5414 10967 5466
rect 10967 5414 10981 5466
rect 11005 5414 11019 5466
rect 11019 5414 11031 5466
rect 11031 5414 11061 5466
rect 11085 5414 11095 5466
rect 11095 5414 11141 5466
rect 10845 5412 10901 5414
rect 10925 5412 10981 5414
rect 11005 5412 11061 5414
rect 11085 5412 11141 5414
rect 13318 10362 13374 10364
rect 13398 10362 13454 10364
rect 13478 10362 13534 10364
rect 13558 10362 13614 10364
rect 13318 10310 13364 10362
rect 13364 10310 13374 10362
rect 13398 10310 13428 10362
rect 13428 10310 13440 10362
rect 13440 10310 13454 10362
rect 13478 10310 13492 10362
rect 13492 10310 13504 10362
rect 13504 10310 13534 10362
rect 13558 10310 13568 10362
rect 13568 10310 13614 10362
rect 13318 10308 13374 10310
rect 13398 10308 13454 10310
rect 13478 10308 13534 10310
rect 13558 10308 13614 10310
rect 13318 9274 13374 9276
rect 13398 9274 13454 9276
rect 13478 9274 13534 9276
rect 13558 9274 13614 9276
rect 13318 9222 13364 9274
rect 13364 9222 13374 9274
rect 13398 9222 13428 9274
rect 13428 9222 13440 9274
rect 13440 9222 13454 9274
rect 13478 9222 13492 9274
rect 13492 9222 13504 9274
rect 13504 9222 13534 9274
rect 13558 9222 13568 9274
rect 13568 9222 13614 9274
rect 13318 9220 13374 9222
rect 13398 9220 13454 9222
rect 13478 9220 13534 9222
rect 13558 9220 13614 9222
rect 13318 8186 13374 8188
rect 13398 8186 13454 8188
rect 13478 8186 13534 8188
rect 13558 8186 13614 8188
rect 13318 8134 13364 8186
rect 13364 8134 13374 8186
rect 13398 8134 13428 8186
rect 13428 8134 13440 8186
rect 13440 8134 13454 8186
rect 13478 8134 13492 8186
rect 13492 8134 13504 8186
rect 13504 8134 13534 8186
rect 13558 8134 13568 8186
rect 13568 8134 13614 8186
rect 13318 8132 13374 8134
rect 13398 8132 13454 8134
rect 13478 8132 13534 8134
rect 13558 8132 13614 8134
rect 13318 7098 13374 7100
rect 13398 7098 13454 7100
rect 13478 7098 13534 7100
rect 13558 7098 13614 7100
rect 13318 7046 13364 7098
rect 13364 7046 13374 7098
rect 13398 7046 13428 7098
rect 13428 7046 13440 7098
rect 13440 7046 13454 7098
rect 13478 7046 13492 7098
rect 13492 7046 13504 7098
rect 13504 7046 13534 7098
rect 13558 7046 13568 7098
rect 13568 7046 13614 7098
rect 13318 7044 13374 7046
rect 13398 7044 13454 7046
rect 13478 7044 13534 7046
rect 13558 7044 13614 7046
rect 13318 6010 13374 6012
rect 13398 6010 13454 6012
rect 13478 6010 13534 6012
rect 13558 6010 13614 6012
rect 13318 5958 13364 6010
rect 13364 5958 13374 6010
rect 13398 5958 13428 6010
rect 13428 5958 13440 6010
rect 13440 5958 13454 6010
rect 13478 5958 13492 6010
rect 13492 5958 13504 6010
rect 13504 5958 13534 6010
rect 13558 5958 13568 6010
rect 13568 5958 13614 6010
rect 13318 5956 13374 5958
rect 13398 5956 13454 5958
rect 13478 5956 13534 5958
rect 13558 5956 13614 5958
rect 10845 4378 10901 4380
rect 10925 4378 10981 4380
rect 11005 4378 11061 4380
rect 11085 4378 11141 4380
rect 10845 4326 10891 4378
rect 10891 4326 10901 4378
rect 10925 4326 10955 4378
rect 10955 4326 10967 4378
rect 10967 4326 10981 4378
rect 11005 4326 11019 4378
rect 11019 4326 11031 4378
rect 11031 4326 11061 4378
rect 11085 4326 11095 4378
rect 11095 4326 11141 4378
rect 10845 4324 10901 4326
rect 10925 4324 10981 4326
rect 11005 4324 11061 4326
rect 11085 4324 11141 4326
rect 13318 4922 13374 4924
rect 13398 4922 13454 4924
rect 13478 4922 13534 4924
rect 13558 4922 13614 4924
rect 13318 4870 13364 4922
rect 13364 4870 13374 4922
rect 13398 4870 13428 4922
rect 13428 4870 13440 4922
rect 13440 4870 13454 4922
rect 13478 4870 13492 4922
rect 13492 4870 13504 4922
rect 13504 4870 13534 4922
rect 13558 4870 13568 4922
rect 13568 4870 13614 4922
rect 13318 4868 13374 4870
rect 13398 4868 13454 4870
rect 13478 4868 13534 4870
rect 13558 4868 13614 4870
rect 13318 3834 13374 3836
rect 13398 3834 13454 3836
rect 13478 3834 13534 3836
rect 13558 3834 13614 3836
rect 13318 3782 13364 3834
rect 13364 3782 13374 3834
rect 13398 3782 13428 3834
rect 13428 3782 13440 3834
rect 13440 3782 13454 3834
rect 13478 3782 13492 3834
rect 13492 3782 13504 3834
rect 13504 3782 13534 3834
rect 13558 3782 13568 3834
rect 13568 3782 13614 3834
rect 13318 3780 13374 3782
rect 13398 3780 13454 3782
rect 13478 3780 13534 3782
rect 13558 3780 13614 3782
rect 10845 3290 10901 3292
rect 10925 3290 10981 3292
rect 11005 3290 11061 3292
rect 11085 3290 11141 3292
rect 10845 3238 10891 3290
rect 10891 3238 10901 3290
rect 10925 3238 10955 3290
rect 10955 3238 10967 3290
rect 10967 3238 10981 3290
rect 11005 3238 11019 3290
rect 11019 3238 11031 3290
rect 11031 3238 11061 3290
rect 11085 3238 11095 3290
rect 11095 3238 11141 3290
rect 10845 3236 10901 3238
rect 10925 3236 10981 3238
rect 11005 3236 11061 3238
rect 11085 3236 11141 3238
rect 13318 2746 13374 2748
rect 13398 2746 13454 2748
rect 13478 2746 13534 2748
rect 13558 2746 13614 2748
rect 13318 2694 13364 2746
rect 13364 2694 13374 2746
rect 13398 2694 13428 2746
rect 13428 2694 13440 2746
rect 13440 2694 13454 2746
rect 13478 2694 13492 2746
rect 13492 2694 13504 2746
rect 13504 2694 13534 2746
rect 13558 2694 13568 2746
rect 13568 2694 13614 2746
rect 13318 2692 13374 2694
rect 13398 2692 13454 2694
rect 13478 2692 13534 2694
rect 13558 2692 13614 2694
rect 14738 16516 14794 16552
rect 14738 16496 14740 16516
rect 14740 16496 14792 16516
rect 14792 16496 14794 16516
rect 15790 18522 15846 18524
rect 15870 18522 15926 18524
rect 15950 18522 16006 18524
rect 16030 18522 16086 18524
rect 15790 18470 15836 18522
rect 15836 18470 15846 18522
rect 15870 18470 15900 18522
rect 15900 18470 15912 18522
rect 15912 18470 15926 18522
rect 15950 18470 15964 18522
rect 15964 18470 15976 18522
rect 15976 18470 16006 18522
rect 16030 18470 16040 18522
rect 16040 18470 16086 18522
rect 15790 18468 15846 18470
rect 15870 18468 15926 18470
rect 15950 18468 16006 18470
rect 16030 18468 16086 18470
rect 18263 19066 18319 19068
rect 18343 19066 18399 19068
rect 18423 19066 18479 19068
rect 18503 19066 18559 19068
rect 18263 19014 18309 19066
rect 18309 19014 18319 19066
rect 18343 19014 18373 19066
rect 18373 19014 18385 19066
rect 18385 19014 18399 19066
rect 18423 19014 18437 19066
rect 18437 19014 18449 19066
rect 18449 19014 18479 19066
rect 18503 19014 18513 19066
rect 18513 19014 18559 19066
rect 18263 19012 18319 19014
rect 18343 19012 18399 19014
rect 18423 19012 18479 19014
rect 18503 19012 18559 19014
rect 15790 17434 15846 17436
rect 15870 17434 15926 17436
rect 15950 17434 16006 17436
rect 16030 17434 16086 17436
rect 15790 17382 15836 17434
rect 15836 17382 15846 17434
rect 15870 17382 15900 17434
rect 15900 17382 15912 17434
rect 15912 17382 15926 17434
rect 15950 17382 15964 17434
rect 15964 17382 15976 17434
rect 15976 17382 16006 17434
rect 16030 17382 16040 17434
rect 16040 17382 16086 17434
rect 15790 17380 15846 17382
rect 15870 17380 15926 17382
rect 15950 17380 16006 17382
rect 16030 17380 16086 17382
rect 15790 16346 15846 16348
rect 15870 16346 15926 16348
rect 15950 16346 16006 16348
rect 16030 16346 16086 16348
rect 15790 16294 15836 16346
rect 15836 16294 15846 16346
rect 15870 16294 15900 16346
rect 15900 16294 15912 16346
rect 15912 16294 15926 16346
rect 15950 16294 15964 16346
rect 15964 16294 15976 16346
rect 15976 16294 16006 16346
rect 16030 16294 16040 16346
rect 16040 16294 16086 16346
rect 15790 16292 15846 16294
rect 15870 16292 15926 16294
rect 15950 16292 16006 16294
rect 16030 16292 16086 16294
rect 15790 15258 15846 15260
rect 15870 15258 15926 15260
rect 15950 15258 16006 15260
rect 16030 15258 16086 15260
rect 15790 15206 15836 15258
rect 15836 15206 15846 15258
rect 15870 15206 15900 15258
rect 15900 15206 15912 15258
rect 15912 15206 15926 15258
rect 15950 15206 15964 15258
rect 15964 15206 15976 15258
rect 15976 15206 16006 15258
rect 16030 15206 16040 15258
rect 16040 15206 16086 15258
rect 15790 15204 15846 15206
rect 15870 15204 15926 15206
rect 15950 15204 16006 15206
rect 16030 15204 16086 15206
rect 15790 14170 15846 14172
rect 15870 14170 15926 14172
rect 15950 14170 16006 14172
rect 16030 14170 16086 14172
rect 15790 14118 15836 14170
rect 15836 14118 15846 14170
rect 15870 14118 15900 14170
rect 15900 14118 15912 14170
rect 15912 14118 15926 14170
rect 15950 14118 15964 14170
rect 15964 14118 15976 14170
rect 15976 14118 16006 14170
rect 16030 14118 16040 14170
rect 16040 14118 16086 14170
rect 15790 14116 15846 14118
rect 15870 14116 15926 14118
rect 15950 14116 16006 14118
rect 16030 14116 16086 14118
rect 15790 13082 15846 13084
rect 15870 13082 15926 13084
rect 15950 13082 16006 13084
rect 16030 13082 16086 13084
rect 15790 13030 15836 13082
rect 15836 13030 15846 13082
rect 15870 13030 15900 13082
rect 15900 13030 15912 13082
rect 15912 13030 15926 13082
rect 15950 13030 15964 13082
rect 15964 13030 15976 13082
rect 15976 13030 16006 13082
rect 16030 13030 16040 13082
rect 16040 13030 16086 13082
rect 15790 13028 15846 13030
rect 15870 13028 15926 13030
rect 15950 13028 16006 13030
rect 16030 13028 16086 13030
rect 20735 18522 20791 18524
rect 20815 18522 20871 18524
rect 20895 18522 20951 18524
rect 20975 18522 21031 18524
rect 20735 18470 20781 18522
rect 20781 18470 20791 18522
rect 20815 18470 20845 18522
rect 20845 18470 20857 18522
rect 20857 18470 20871 18522
rect 20895 18470 20909 18522
rect 20909 18470 20921 18522
rect 20921 18470 20951 18522
rect 20975 18470 20985 18522
rect 20985 18470 21031 18522
rect 20735 18468 20791 18470
rect 20815 18468 20871 18470
rect 20895 18468 20951 18470
rect 20975 18468 21031 18470
rect 18263 17978 18319 17980
rect 18343 17978 18399 17980
rect 18423 17978 18479 17980
rect 18503 17978 18559 17980
rect 18263 17926 18309 17978
rect 18309 17926 18319 17978
rect 18343 17926 18373 17978
rect 18373 17926 18385 17978
rect 18385 17926 18399 17978
rect 18423 17926 18437 17978
rect 18437 17926 18449 17978
rect 18449 17926 18479 17978
rect 18503 17926 18513 17978
rect 18513 17926 18559 17978
rect 18263 17924 18319 17926
rect 18343 17924 18399 17926
rect 18423 17924 18479 17926
rect 18503 17924 18559 17926
rect 18263 16890 18319 16892
rect 18343 16890 18399 16892
rect 18423 16890 18479 16892
rect 18503 16890 18559 16892
rect 18263 16838 18309 16890
rect 18309 16838 18319 16890
rect 18343 16838 18373 16890
rect 18373 16838 18385 16890
rect 18385 16838 18399 16890
rect 18423 16838 18437 16890
rect 18437 16838 18449 16890
rect 18449 16838 18479 16890
rect 18503 16838 18513 16890
rect 18513 16838 18559 16890
rect 18263 16836 18319 16838
rect 18343 16836 18399 16838
rect 18423 16836 18479 16838
rect 18503 16836 18559 16838
rect 18142 16632 18198 16688
rect 18050 16516 18106 16552
rect 18050 16496 18052 16516
rect 18052 16496 18104 16516
rect 18104 16496 18106 16516
rect 20735 17434 20791 17436
rect 20815 17434 20871 17436
rect 20895 17434 20951 17436
rect 20975 17434 21031 17436
rect 20735 17382 20781 17434
rect 20781 17382 20791 17434
rect 20815 17382 20845 17434
rect 20845 17382 20857 17434
rect 20857 17382 20871 17434
rect 20895 17382 20909 17434
rect 20909 17382 20921 17434
rect 20921 17382 20951 17434
rect 20975 17382 20985 17434
rect 20985 17382 21031 17434
rect 20735 17380 20791 17382
rect 20815 17380 20871 17382
rect 20895 17380 20951 17382
rect 20975 17380 21031 17382
rect 20735 16346 20791 16348
rect 20815 16346 20871 16348
rect 20895 16346 20951 16348
rect 20975 16346 21031 16348
rect 20735 16294 20781 16346
rect 20781 16294 20791 16346
rect 20815 16294 20845 16346
rect 20845 16294 20857 16346
rect 20857 16294 20871 16346
rect 20895 16294 20909 16346
rect 20909 16294 20921 16346
rect 20921 16294 20951 16346
rect 20975 16294 20985 16346
rect 20985 16294 21031 16346
rect 20735 16292 20791 16294
rect 20815 16292 20871 16294
rect 20895 16292 20951 16294
rect 20975 16292 21031 16294
rect 15790 11994 15846 11996
rect 15870 11994 15926 11996
rect 15950 11994 16006 11996
rect 16030 11994 16086 11996
rect 15790 11942 15836 11994
rect 15836 11942 15846 11994
rect 15870 11942 15900 11994
rect 15900 11942 15912 11994
rect 15912 11942 15926 11994
rect 15950 11942 15964 11994
rect 15964 11942 15976 11994
rect 15976 11942 16006 11994
rect 16030 11942 16040 11994
rect 16040 11942 16086 11994
rect 15790 11940 15846 11942
rect 15870 11940 15926 11942
rect 15950 11940 16006 11942
rect 16030 11940 16086 11942
rect 15790 10906 15846 10908
rect 15870 10906 15926 10908
rect 15950 10906 16006 10908
rect 16030 10906 16086 10908
rect 15790 10854 15836 10906
rect 15836 10854 15846 10906
rect 15870 10854 15900 10906
rect 15900 10854 15912 10906
rect 15912 10854 15926 10906
rect 15950 10854 15964 10906
rect 15964 10854 15976 10906
rect 15976 10854 16006 10906
rect 16030 10854 16040 10906
rect 16040 10854 16086 10906
rect 15790 10852 15846 10854
rect 15870 10852 15926 10854
rect 15950 10852 16006 10854
rect 16030 10852 16086 10854
rect 15790 9818 15846 9820
rect 15870 9818 15926 9820
rect 15950 9818 16006 9820
rect 16030 9818 16086 9820
rect 15790 9766 15836 9818
rect 15836 9766 15846 9818
rect 15870 9766 15900 9818
rect 15900 9766 15912 9818
rect 15912 9766 15926 9818
rect 15950 9766 15964 9818
rect 15964 9766 15976 9818
rect 15976 9766 16006 9818
rect 16030 9766 16040 9818
rect 16040 9766 16086 9818
rect 15790 9764 15846 9766
rect 15870 9764 15926 9766
rect 15950 9764 16006 9766
rect 16030 9764 16086 9766
rect 14462 6024 14518 6080
rect 15790 8730 15846 8732
rect 15870 8730 15926 8732
rect 15950 8730 16006 8732
rect 16030 8730 16086 8732
rect 15790 8678 15836 8730
rect 15836 8678 15846 8730
rect 15870 8678 15900 8730
rect 15900 8678 15912 8730
rect 15912 8678 15926 8730
rect 15950 8678 15964 8730
rect 15964 8678 15976 8730
rect 15976 8678 16006 8730
rect 16030 8678 16040 8730
rect 16040 8678 16086 8730
rect 15790 8676 15846 8678
rect 15870 8676 15926 8678
rect 15950 8676 16006 8678
rect 16030 8676 16086 8678
rect 15790 7642 15846 7644
rect 15870 7642 15926 7644
rect 15950 7642 16006 7644
rect 16030 7642 16086 7644
rect 15790 7590 15836 7642
rect 15836 7590 15846 7642
rect 15870 7590 15900 7642
rect 15900 7590 15912 7642
rect 15912 7590 15926 7642
rect 15950 7590 15964 7642
rect 15964 7590 15976 7642
rect 15976 7590 16006 7642
rect 16030 7590 16040 7642
rect 16040 7590 16086 7642
rect 15790 7588 15846 7590
rect 15870 7588 15926 7590
rect 15950 7588 16006 7590
rect 16030 7588 16086 7590
rect 15790 6554 15846 6556
rect 15870 6554 15926 6556
rect 15950 6554 16006 6556
rect 16030 6554 16086 6556
rect 15790 6502 15836 6554
rect 15836 6502 15846 6554
rect 15870 6502 15900 6554
rect 15900 6502 15912 6554
rect 15912 6502 15926 6554
rect 15950 6502 15964 6554
rect 15964 6502 15976 6554
rect 15976 6502 16006 6554
rect 16030 6502 16040 6554
rect 16040 6502 16086 6554
rect 15790 6500 15846 6502
rect 15870 6500 15926 6502
rect 15950 6500 16006 6502
rect 16030 6500 16086 6502
rect 16394 6296 16450 6352
rect 15790 5466 15846 5468
rect 15870 5466 15926 5468
rect 15950 5466 16006 5468
rect 16030 5466 16086 5468
rect 15790 5414 15836 5466
rect 15836 5414 15846 5466
rect 15870 5414 15900 5466
rect 15900 5414 15912 5466
rect 15912 5414 15926 5466
rect 15950 5414 15964 5466
rect 15964 5414 15976 5466
rect 15976 5414 16006 5466
rect 16030 5414 16040 5466
rect 16040 5414 16086 5466
rect 15790 5412 15846 5414
rect 15870 5412 15926 5414
rect 15950 5412 16006 5414
rect 16030 5412 16086 5414
rect 18263 15802 18319 15804
rect 18343 15802 18399 15804
rect 18423 15802 18479 15804
rect 18503 15802 18559 15804
rect 18263 15750 18309 15802
rect 18309 15750 18319 15802
rect 18343 15750 18373 15802
rect 18373 15750 18385 15802
rect 18385 15750 18399 15802
rect 18423 15750 18437 15802
rect 18437 15750 18449 15802
rect 18449 15750 18479 15802
rect 18503 15750 18513 15802
rect 18513 15750 18559 15802
rect 18263 15748 18319 15750
rect 18343 15748 18399 15750
rect 18423 15748 18479 15750
rect 18503 15748 18559 15750
rect 20735 15258 20791 15260
rect 20815 15258 20871 15260
rect 20895 15258 20951 15260
rect 20975 15258 21031 15260
rect 20735 15206 20781 15258
rect 20781 15206 20791 15258
rect 20815 15206 20845 15258
rect 20845 15206 20857 15258
rect 20857 15206 20871 15258
rect 20895 15206 20909 15258
rect 20909 15206 20921 15258
rect 20921 15206 20951 15258
rect 20975 15206 20985 15258
rect 20985 15206 21031 15258
rect 20735 15204 20791 15206
rect 20815 15204 20871 15206
rect 20895 15204 20951 15206
rect 20975 15204 21031 15206
rect 18263 14714 18319 14716
rect 18343 14714 18399 14716
rect 18423 14714 18479 14716
rect 18503 14714 18559 14716
rect 18263 14662 18309 14714
rect 18309 14662 18319 14714
rect 18343 14662 18373 14714
rect 18373 14662 18385 14714
rect 18385 14662 18399 14714
rect 18423 14662 18437 14714
rect 18437 14662 18449 14714
rect 18449 14662 18479 14714
rect 18503 14662 18513 14714
rect 18513 14662 18559 14714
rect 18263 14660 18319 14662
rect 18343 14660 18399 14662
rect 18423 14660 18479 14662
rect 18503 14660 18559 14662
rect 18263 13626 18319 13628
rect 18343 13626 18399 13628
rect 18423 13626 18479 13628
rect 18503 13626 18559 13628
rect 18263 13574 18309 13626
rect 18309 13574 18319 13626
rect 18343 13574 18373 13626
rect 18373 13574 18385 13626
rect 18385 13574 18399 13626
rect 18423 13574 18437 13626
rect 18437 13574 18449 13626
rect 18449 13574 18479 13626
rect 18503 13574 18513 13626
rect 18513 13574 18559 13626
rect 18263 13572 18319 13574
rect 18343 13572 18399 13574
rect 18423 13572 18479 13574
rect 18503 13572 18559 13574
rect 18263 12538 18319 12540
rect 18343 12538 18399 12540
rect 18423 12538 18479 12540
rect 18503 12538 18559 12540
rect 18263 12486 18309 12538
rect 18309 12486 18319 12538
rect 18343 12486 18373 12538
rect 18373 12486 18385 12538
rect 18385 12486 18399 12538
rect 18423 12486 18437 12538
rect 18437 12486 18449 12538
rect 18449 12486 18479 12538
rect 18503 12486 18513 12538
rect 18513 12486 18559 12538
rect 18263 12484 18319 12486
rect 18343 12484 18399 12486
rect 18423 12484 18479 12486
rect 18503 12484 18559 12486
rect 20735 14170 20791 14172
rect 20815 14170 20871 14172
rect 20895 14170 20951 14172
rect 20975 14170 21031 14172
rect 20735 14118 20781 14170
rect 20781 14118 20791 14170
rect 20815 14118 20845 14170
rect 20845 14118 20857 14170
rect 20857 14118 20871 14170
rect 20895 14118 20909 14170
rect 20909 14118 20921 14170
rect 20921 14118 20951 14170
rect 20975 14118 20985 14170
rect 20985 14118 21031 14170
rect 20735 14116 20791 14118
rect 20815 14116 20871 14118
rect 20895 14116 20951 14118
rect 20975 14116 21031 14118
rect 20735 13082 20791 13084
rect 20815 13082 20871 13084
rect 20895 13082 20951 13084
rect 20975 13082 21031 13084
rect 20735 13030 20781 13082
rect 20781 13030 20791 13082
rect 20815 13030 20845 13082
rect 20845 13030 20857 13082
rect 20857 13030 20871 13082
rect 20895 13030 20909 13082
rect 20909 13030 20921 13082
rect 20921 13030 20951 13082
rect 20975 13030 20985 13082
rect 20985 13030 21031 13082
rect 20735 13028 20791 13030
rect 20815 13028 20871 13030
rect 20895 13028 20951 13030
rect 20975 13028 21031 13030
rect 20735 11994 20791 11996
rect 20815 11994 20871 11996
rect 20895 11994 20951 11996
rect 20975 11994 21031 11996
rect 20735 11942 20781 11994
rect 20781 11942 20791 11994
rect 20815 11942 20845 11994
rect 20845 11942 20857 11994
rect 20857 11942 20871 11994
rect 20895 11942 20909 11994
rect 20909 11942 20921 11994
rect 20921 11942 20951 11994
rect 20975 11942 20985 11994
rect 20985 11942 21031 11994
rect 20735 11940 20791 11942
rect 20815 11940 20871 11942
rect 20895 11940 20951 11942
rect 20975 11940 21031 11942
rect 18263 11450 18319 11452
rect 18343 11450 18399 11452
rect 18423 11450 18479 11452
rect 18503 11450 18559 11452
rect 18263 11398 18309 11450
rect 18309 11398 18319 11450
rect 18343 11398 18373 11450
rect 18373 11398 18385 11450
rect 18385 11398 18399 11450
rect 18423 11398 18437 11450
rect 18437 11398 18449 11450
rect 18449 11398 18479 11450
rect 18503 11398 18513 11450
rect 18513 11398 18559 11450
rect 18263 11396 18319 11398
rect 18343 11396 18399 11398
rect 18423 11396 18479 11398
rect 18503 11396 18559 11398
rect 18263 10362 18319 10364
rect 18343 10362 18399 10364
rect 18423 10362 18479 10364
rect 18503 10362 18559 10364
rect 18263 10310 18309 10362
rect 18309 10310 18319 10362
rect 18343 10310 18373 10362
rect 18373 10310 18385 10362
rect 18385 10310 18399 10362
rect 18423 10310 18437 10362
rect 18437 10310 18449 10362
rect 18449 10310 18479 10362
rect 18503 10310 18513 10362
rect 18513 10310 18559 10362
rect 18263 10308 18319 10310
rect 18343 10308 18399 10310
rect 18423 10308 18479 10310
rect 18503 10308 18559 10310
rect 18263 9274 18319 9276
rect 18343 9274 18399 9276
rect 18423 9274 18479 9276
rect 18503 9274 18559 9276
rect 18263 9222 18309 9274
rect 18309 9222 18319 9274
rect 18343 9222 18373 9274
rect 18373 9222 18385 9274
rect 18385 9222 18399 9274
rect 18423 9222 18437 9274
rect 18437 9222 18449 9274
rect 18449 9222 18479 9274
rect 18503 9222 18513 9274
rect 18513 9222 18559 9274
rect 18263 9220 18319 9222
rect 18343 9220 18399 9222
rect 18423 9220 18479 9222
rect 18503 9220 18559 9222
rect 18263 8186 18319 8188
rect 18343 8186 18399 8188
rect 18423 8186 18479 8188
rect 18503 8186 18559 8188
rect 18263 8134 18309 8186
rect 18309 8134 18319 8186
rect 18343 8134 18373 8186
rect 18373 8134 18385 8186
rect 18385 8134 18399 8186
rect 18423 8134 18437 8186
rect 18437 8134 18449 8186
rect 18449 8134 18479 8186
rect 18503 8134 18513 8186
rect 18513 8134 18559 8186
rect 18263 8132 18319 8134
rect 18343 8132 18399 8134
rect 18423 8132 18479 8134
rect 18503 8132 18559 8134
rect 18263 7098 18319 7100
rect 18343 7098 18399 7100
rect 18423 7098 18479 7100
rect 18503 7098 18559 7100
rect 18263 7046 18309 7098
rect 18309 7046 18319 7098
rect 18343 7046 18373 7098
rect 18373 7046 18385 7098
rect 18385 7046 18399 7098
rect 18423 7046 18437 7098
rect 18437 7046 18449 7098
rect 18449 7046 18479 7098
rect 18503 7046 18513 7098
rect 18513 7046 18559 7098
rect 18263 7044 18319 7046
rect 18343 7044 18399 7046
rect 18423 7044 18479 7046
rect 18503 7044 18559 7046
rect 17866 6060 17868 6080
rect 17868 6060 17920 6080
rect 17920 6060 17922 6080
rect 17866 6024 17922 6060
rect 18263 6010 18319 6012
rect 18343 6010 18399 6012
rect 18423 6010 18479 6012
rect 18503 6010 18559 6012
rect 18263 5958 18309 6010
rect 18309 5958 18319 6010
rect 18343 5958 18373 6010
rect 18373 5958 18385 6010
rect 18385 5958 18399 6010
rect 18423 5958 18437 6010
rect 18437 5958 18449 6010
rect 18449 5958 18479 6010
rect 18503 5958 18513 6010
rect 18513 5958 18559 6010
rect 18263 5956 18319 5958
rect 18343 5956 18399 5958
rect 18423 5956 18479 5958
rect 18503 5956 18559 5958
rect 18263 4922 18319 4924
rect 18343 4922 18399 4924
rect 18423 4922 18479 4924
rect 18503 4922 18559 4924
rect 18263 4870 18309 4922
rect 18309 4870 18319 4922
rect 18343 4870 18373 4922
rect 18373 4870 18385 4922
rect 18385 4870 18399 4922
rect 18423 4870 18437 4922
rect 18437 4870 18449 4922
rect 18449 4870 18479 4922
rect 18503 4870 18513 4922
rect 18513 4870 18559 4922
rect 18263 4868 18319 4870
rect 18343 4868 18399 4870
rect 18423 4868 18479 4870
rect 18503 4868 18559 4870
rect 20735 10906 20791 10908
rect 20815 10906 20871 10908
rect 20895 10906 20951 10908
rect 20975 10906 21031 10908
rect 20735 10854 20781 10906
rect 20781 10854 20791 10906
rect 20815 10854 20845 10906
rect 20845 10854 20857 10906
rect 20857 10854 20871 10906
rect 20895 10854 20909 10906
rect 20909 10854 20921 10906
rect 20921 10854 20951 10906
rect 20975 10854 20985 10906
rect 20985 10854 21031 10906
rect 20735 10852 20791 10854
rect 20815 10852 20871 10854
rect 20895 10852 20951 10854
rect 20975 10852 21031 10854
rect 20735 9818 20791 9820
rect 20815 9818 20871 9820
rect 20895 9818 20951 9820
rect 20975 9818 21031 9820
rect 20735 9766 20781 9818
rect 20781 9766 20791 9818
rect 20815 9766 20845 9818
rect 20845 9766 20857 9818
rect 20857 9766 20871 9818
rect 20895 9766 20909 9818
rect 20909 9766 20921 9818
rect 20921 9766 20951 9818
rect 20975 9766 20985 9818
rect 20985 9766 21031 9818
rect 20735 9764 20791 9766
rect 20815 9764 20871 9766
rect 20895 9764 20951 9766
rect 20975 9764 21031 9766
rect 20735 8730 20791 8732
rect 20815 8730 20871 8732
rect 20895 8730 20951 8732
rect 20975 8730 21031 8732
rect 20735 8678 20781 8730
rect 20781 8678 20791 8730
rect 20815 8678 20845 8730
rect 20845 8678 20857 8730
rect 20857 8678 20871 8730
rect 20895 8678 20909 8730
rect 20909 8678 20921 8730
rect 20921 8678 20951 8730
rect 20975 8678 20985 8730
rect 20985 8678 21031 8730
rect 20735 8676 20791 8678
rect 20815 8676 20871 8678
rect 20895 8676 20951 8678
rect 20975 8676 21031 8678
rect 20735 7642 20791 7644
rect 20815 7642 20871 7644
rect 20895 7642 20951 7644
rect 20975 7642 21031 7644
rect 20735 7590 20781 7642
rect 20781 7590 20791 7642
rect 20815 7590 20845 7642
rect 20845 7590 20857 7642
rect 20857 7590 20871 7642
rect 20895 7590 20909 7642
rect 20909 7590 20921 7642
rect 20921 7590 20951 7642
rect 20975 7590 20985 7642
rect 20985 7590 21031 7642
rect 20735 7588 20791 7590
rect 20815 7588 20871 7590
rect 20895 7588 20951 7590
rect 20975 7588 21031 7590
rect 20735 6554 20791 6556
rect 20815 6554 20871 6556
rect 20895 6554 20951 6556
rect 20975 6554 21031 6556
rect 20735 6502 20781 6554
rect 20781 6502 20791 6554
rect 20815 6502 20845 6554
rect 20845 6502 20857 6554
rect 20857 6502 20871 6554
rect 20895 6502 20909 6554
rect 20909 6502 20921 6554
rect 20921 6502 20951 6554
rect 20975 6502 20985 6554
rect 20985 6502 21031 6554
rect 20735 6500 20791 6502
rect 20815 6500 20871 6502
rect 20895 6500 20951 6502
rect 20975 6500 21031 6502
rect 15790 4378 15846 4380
rect 15870 4378 15926 4380
rect 15950 4378 16006 4380
rect 16030 4378 16086 4380
rect 15790 4326 15836 4378
rect 15836 4326 15846 4378
rect 15870 4326 15900 4378
rect 15900 4326 15912 4378
rect 15912 4326 15926 4378
rect 15950 4326 15964 4378
rect 15964 4326 15976 4378
rect 15976 4326 16006 4378
rect 16030 4326 16040 4378
rect 16040 4326 16086 4378
rect 15790 4324 15846 4326
rect 15870 4324 15926 4326
rect 15950 4324 16006 4326
rect 16030 4324 16086 4326
rect 18263 3834 18319 3836
rect 18343 3834 18399 3836
rect 18423 3834 18479 3836
rect 18503 3834 18559 3836
rect 18263 3782 18309 3834
rect 18309 3782 18319 3834
rect 18343 3782 18373 3834
rect 18373 3782 18385 3834
rect 18385 3782 18399 3834
rect 18423 3782 18437 3834
rect 18437 3782 18449 3834
rect 18449 3782 18479 3834
rect 18503 3782 18513 3834
rect 18513 3782 18559 3834
rect 18263 3780 18319 3782
rect 18343 3780 18399 3782
rect 18423 3780 18479 3782
rect 18503 3780 18559 3782
rect 15790 3290 15846 3292
rect 15870 3290 15926 3292
rect 15950 3290 16006 3292
rect 16030 3290 16086 3292
rect 15790 3238 15836 3290
rect 15836 3238 15846 3290
rect 15870 3238 15900 3290
rect 15900 3238 15912 3290
rect 15912 3238 15926 3290
rect 15950 3238 15964 3290
rect 15964 3238 15976 3290
rect 15976 3238 16006 3290
rect 16030 3238 16040 3290
rect 16040 3238 16086 3290
rect 15790 3236 15846 3238
rect 15870 3236 15926 3238
rect 15950 3236 16006 3238
rect 16030 3236 16086 3238
rect 18263 2746 18319 2748
rect 18343 2746 18399 2748
rect 18423 2746 18479 2748
rect 18503 2746 18559 2748
rect 18263 2694 18309 2746
rect 18309 2694 18319 2746
rect 18343 2694 18373 2746
rect 18373 2694 18385 2746
rect 18385 2694 18399 2746
rect 18423 2694 18437 2746
rect 18437 2694 18449 2746
rect 18449 2694 18479 2746
rect 18503 2694 18513 2746
rect 18513 2694 18559 2746
rect 18263 2692 18319 2694
rect 18343 2692 18399 2694
rect 18423 2692 18479 2694
rect 18503 2692 18559 2694
rect 20735 5466 20791 5468
rect 20815 5466 20871 5468
rect 20895 5466 20951 5468
rect 20975 5466 21031 5468
rect 20735 5414 20781 5466
rect 20781 5414 20791 5466
rect 20815 5414 20845 5466
rect 20845 5414 20857 5466
rect 20857 5414 20871 5466
rect 20895 5414 20909 5466
rect 20909 5414 20921 5466
rect 20921 5414 20951 5466
rect 20975 5414 20985 5466
rect 20985 5414 21031 5466
rect 20735 5412 20791 5414
rect 20815 5412 20871 5414
rect 20895 5412 20951 5414
rect 20975 5412 21031 5414
rect 20735 4378 20791 4380
rect 20815 4378 20871 4380
rect 20895 4378 20951 4380
rect 20975 4378 21031 4380
rect 20735 4326 20781 4378
rect 20781 4326 20791 4378
rect 20815 4326 20845 4378
rect 20845 4326 20857 4378
rect 20857 4326 20871 4378
rect 20895 4326 20909 4378
rect 20909 4326 20921 4378
rect 20921 4326 20951 4378
rect 20975 4326 20985 4378
rect 20985 4326 21031 4378
rect 20735 4324 20791 4326
rect 20815 4324 20871 4326
rect 20895 4324 20951 4326
rect 20975 4324 21031 4326
rect 20735 3290 20791 3292
rect 20815 3290 20871 3292
rect 20895 3290 20951 3292
rect 20975 3290 21031 3292
rect 20735 3238 20781 3290
rect 20781 3238 20791 3290
rect 20815 3238 20845 3290
rect 20845 3238 20857 3290
rect 20857 3238 20871 3290
rect 20895 3238 20909 3290
rect 20909 3238 20921 3290
rect 20921 3238 20951 3290
rect 20975 3238 20985 3290
rect 20985 3238 21031 3290
rect 20735 3236 20791 3238
rect 20815 3236 20871 3238
rect 20895 3236 20951 3238
rect 20975 3236 21031 3238
rect 5900 2202 5956 2204
rect 5980 2202 6036 2204
rect 6060 2202 6116 2204
rect 6140 2202 6196 2204
rect 5900 2150 5946 2202
rect 5946 2150 5956 2202
rect 5980 2150 6010 2202
rect 6010 2150 6022 2202
rect 6022 2150 6036 2202
rect 6060 2150 6074 2202
rect 6074 2150 6086 2202
rect 6086 2150 6116 2202
rect 6140 2150 6150 2202
rect 6150 2150 6196 2202
rect 5900 2148 5956 2150
rect 5980 2148 6036 2150
rect 6060 2148 6116 2150
rect 6140 2148 6196 2150
rect 10845 2202 10901 2204
rect 10925 2202 10981 2204
rect 11005 2202 11061 2204
rect 11085 2202 11141 2204
rect 10845 2150 10891 2202
rect 10891 2150 10901 2202
rect 10925 2150 10955 2202
rect 10955 2150 10967 2202
rect 10967 2150 10981 2202
rect 11005 2150 11019 2202
rect 11019 2150 11031 2202
rect 11031 2150 11061 2202
rect 11085 2150 11095 2202
rect 11095 2150 11141 2202
rect 10845 2148 10901 2150
rect 10925 2148 10981 2150
rect 11005 2148 11061 2150
rect 11085 2148 11141 2150
rect 15790 2202 15846 2204
rect 15870 2202 15926 2204
rect 15950 2202 16006 2204
rect 16030 2202 16086 2204
rect 15790 2150 15836 2202
rect 15836 2150 15846 2202
rect 15870 2150 15900 2202
rect 15900 2150 15912 2202
rect 15912 2150 15926 2202
rect 15950 2150 15964 2202
rect 15964 2150 15976 2202
rect 15976 2150 16006 2202
rect 16030 2150 16040 2202
rect 16040 2150 16086 2202
rect 15790 2148 15846 2150
rect 15870 2148 15926 2150
rect 15950 2148 16006 2150
rect 16030 2148 16086 2150
rect 20735 2202 20791 2204
rect 20815 2202 20871 2204
rect 20895 2202 20951 2204
rect 20975 2202 21031 2204
rect 20735 2150 20781 2202
rect 20781 2150 20791 2202
rect 20815 2150 20845 2202
rect 20845 2150 20857 2202
rect 20857 2150 20871 2202
rect 20895 2150 20909 2202
rect 20909 2150 20921 2202
rect 20921 2150 20951 2202
rect 20975 2150 20985 2202
rect 20985 2150 21031 2202
rect 20735 2148 20791 2150
rect 20815 2148 20871 2150
rect 20895 2148 20951 2150
rect 20975 2148 21031 2150
<< metal3 >>
rect 5890 19616 6206 19617
rect 5890 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6206 19616
rect 5890 19551 6206 19552
rect 10835 19616 11151 19617
rect 10835 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11151 19616
rect 10835 19551 11151 19552
rect 15780 19616 16096 19617
rect 15780 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16096 19616
rect 15780 19551 16096 19552
rect 20725 19616 21041 19617
rect 20725 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21041 19616
rect 20725 19551 21041 19552
rect 3418 19072 3734 19073
rect 3418 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3734 19072
rect 3418 19007 3734 19008
rect 8363 19072 8679 19073
rect 8363 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8679 19072
rect 8363 19007 8679 19008
rect 13308 19072 13624 19073
rect 13308 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13624 19072
rect 13308 19007 13624 19008
rect 18253 19072 18569 19073
rect 18253 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18569 19072
rect 18253 19007 18569 19008
rect 5890 18528 6206 18529
rect 5890 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6206 18528
rect 5890 18463 6206 18464
rect 10835 18528 11151 18529
rect 10835 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11151 18528
rect 10835 18463 11151 18464
rect 15780 18528 16096 18529
rect 15780 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16096 18528
rect 15780 18463 16096 18464
rect 20725 18528 21041 18529
rect 20725 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21041 18528
rect 20725 18463 21041 18464
rect 8201 18322 8267 18325
rect 15193 18322 15259 18325
rect 8201 18320 15259 18322
rect 8201 18264 8206 18320
rect 8262 18264 15198 18320
rect 15254 18264 15259 18320
rect 8201 18262 15259 18264
rect 8201 18259 8267 18262
rect 15193 18259 15259 18262
rect 3418 17984 3734 17985
rect 3418 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3734 17984
rect 3418 17919 3734 17920
rect 8363 17984 8679 17985
rect 8363 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8679 17984
rect 8363 17919 8679 17920
rect 13308 17984 13624 17985
rect 13308 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13624 17984
rect 13308 17919 13624 17920
rect 18253 17984 18569 17985
rect 18253 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18569 17984
rect 18253 17919 18569 17920
rect 5890 17440 6206 17441
rect 5890 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6206 17440
rect 5890 17375 6206 17376
rect 10835 17440 11151 17441
rect 10835 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11151 17440
rect 10835 17375 11151 17376
rect 15780 17440 16096 17441
rect 15780 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16096 17440
rect 15780 17375 16096 17376
rect 20725 17440 21041 17441
rect 20725 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21041 17440
rect 20725 17375 21041 17376
rect 3418 16896 3734 16897
rect 3418 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3734 16896
rect 3418 16831 3734 16832
rect 8363 16896 8679 16897
rect 8363 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8679 16896
rect 8363 16831 8679 16832
rect 13308 16896 13624 16897
rect 13308 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13624 16896
rect 13308 16831 13624 16832
rect 18253 16896 18569 16897
rect 18253 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18569 16896
rect 18253 16831 18569 16832
rect 10501 16690 10567 16693
rect 18137 16690 18203 16693
rect 10501 16688 18203 16690
rect 10501 16632 10506 16688
rect 10562 16632 18142 16688
rect 18198 16632 18203 16688
rect 10501 16630 18203 16632
rect 10501 16627 10567 16630
rect 18137 16627 18203 16630
rect 14733 16554 14799 16557
rect 18045 16554 18111 16557
rect 14733 16552 18111 16554
rect 14733 16496 14738 16552
rect 14794 16496 18050 16552
rect 18106 16496 18111 16552
rect 14733 16494 18111 16496
rect 14733 16491 14799 16494
rect 18045 16491 18111 16494
rect 5890 16352 6206 16353
rect 5890 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6206 16352
rect 5890 16287 6206 16288
rect 10835 16352 11151 16353
rect 10835 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11151 16352
rect 10835 16287 11151 16288
rect 15780 16352 16096 16353
rect 15780 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16096 16352
rect 15780 16287 16096 16288
rect 20725 16352 21041 16353
rect 20725 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21041 16352
rect 20725 16287 21041 16288
rect 3418 15808 3734 15809
rect 3418 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3734 15808
rect 3418 15743 3734 15744
rect 8363 15808 8679 15809
rect 8363 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8679 15808
rect 8363 15743 8679 15744
rect 13308 15808 13624 15809
rect 13308 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13624 15808
rect 13308 15743 13624 15744
rect 18253 15808 18569 15809
rect 18253 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18569 15808
rect 18253 15743 18569 15744
rect 5890 15264 6206 15265
rect 5890 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6206 15264
rect 5890 15199 6206 15200
rect 10835 15264 11151 15265
rect 10835 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11151 15264
rect 10835 15199 11151 15200
rect 15780 15264 16096 15265
rect 15780 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16096 15264
rect 15780 15199 16096 15200
rect 20725 15264 21041 15265
rect 20725 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21041 15264
rect 20725 15199 21041 15200
rect 3418 14720 3734 14721
rect 3418 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3734 14720
rect 3418 14655 3734 14656
rect 8363 14720 8679 14721
rect 8363 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8679 14720
rect 8363 14655 8679 14656
rect 13308 14720 13624 14721
rect 13308 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13624 14720
rect 13308 14655 13624 14656
rect 18253 14720 18569 14721
rect 18253 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18569 14720
rect 18253 14655 18569 14656
rect 5890 14176 6206 14177
rect 5890 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6206 14176
rect 5890 14111 6206 14112
rect 10835 14176 11151 14177
rect 10835 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11151 14176
rect 10835 14111 11151 14112
rect 15780 14176 16096 14177
rect 15780 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16096 14176
rect 15780 14111 16096 14112
rect 20725 14176 21041 14177
rect 20725 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21041 14176
rect 20725 14111 21041 14112
rect 3418 13632 3734 13633
rect 3418 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3734 13632
rect 3418 13567 3734 13568
rect 8363 13632 8679 13633
rect 8363 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8679 13632
rect 8363 13567 8679 13568
rect 13308 13632 13624 13633
rect 13308 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13624 13632
rect 13308 13567 13624 13568
rect 18253 13632 18569 13633
rect 18253 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18569 13632
rect 18253 13567 18569 13568
rect 5890 13088 6206 13089
rect 5890 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6206 13088
rect 5890 13023 6206 13024
rect 10835 13088 11151 13089
rect 10835 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11151 13088
rect 10835 13023 11151 13024
rect 15780 13088 16096 13089
rect 15780 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16096 13088
rect 15780 13023 16096 13024
rect 20725 13088 21041 13089
rect 20725 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21041 13088
rect 20725 13023 21041 13024
rect 3418 12544 3734 12545
rect 3418 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3734 12544
rect 3418 12479 3734 12480
rect 8363 12544 8679 12545
rect 8363 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8679 12544
rect 8363 12479 8679 12480
rect 13308 12544 13624 12545
rect 13308 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13624 12544
rect 13308 12479 13624 12480
rect 18253 12544 18569 12545
rect 18253 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18569 12544
rect 18253 12479 18569 12480
rect 5890 12000 6206 12001
rect 5890 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6206 12000
rect 5890 11935 6206 11936
rect 10835 12000 11151 12001
rect 10835 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11151 12000
rect 10835 11935 11151 11936
rect 15780 12000 16096 12001
rect 15780 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16096 12000
rect 15780 11935 16096 11936
rect 20725 12000 21041 12001
rect 20725 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21041 12000
rect 20725 11935 21041 11936
rect 3418 11456 3734 11457
rect 3418 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3734 11456
rect 3418 11391 3734 11392
rect 8363 11456 8679 11457
rect 8363 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8679 11456
rect 8363 11391 8679 11392
rect 13308 11456 13624 11457
rect 13308 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13624 11456
rect 13308 11391 13624 11392
rect 18253 11456 18569 11457
rect 18253 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18569 11456
rect 18253 11391 18569 11392
rect 5890 10912 6206 10913
rect 5890 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6206 10912
rect 5890 10847 6206 10848
rect 10835 10912 11151 10913
rect 10835 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11151 10912
rect 10835 10847 11151 10848
rect 15780 10912 16096 10913
rect 15780 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16096 10912
rect 15780 10847 16096 10848
rect 20725 10912 21041 10913
rect 20725 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21041 10912
rect 20725 10847 21041 10848
rect 3418 10368 3734 10369
rect 3418 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3734 10368
rect 3418 10303 3734 10304
rect 8363 10368 8679 10369
rect 8363 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8679 10368
rect 8363 10303 8679 10304
rect 13308 10368 13624 10369
rect 13308 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13624 10368
rect 13308 10303 13624 10304
rect 18253 10368 18569 10369
rect 18253 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18569 10368
rect 18253 10303 18569 10304
rect 5890 9824 6206 9825
rect 5890 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6206 9824
rect 5890 9759 6206 9760
rect 10835 9824 11151 9825
rect 10835 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11151 9824
rect 10835 9759 11151 9760
rect 15780 9824 16096 9825
rect 15780 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16096 9824
rect 15780 9759 16096 9760
rect 20725 9824 21041 9825
rect 20725 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21041 9824
rect 20725 9759 21041 9760
rect 3418 9280 3734 9281
rect 3418 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3734 9280
rect 3418 9215 3734 9216
rect 8363 9280 8679 9281
rect 8363 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8679 9280
rect 8363 9215 8679 9216
rect 13308 9280 13624 9281
rect 13308 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13624 9280
rect 13308 9215 13624 9216
rect 18253 9280 18569 9281
rect 18253 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18569 9280
rect 18253 9215 18569 9216
rect 5890 8736 6206 8737
rect 5890 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6206 8736
rect 5890 8671 6206 8672
rect 10835 8736 11151 8737
rect 10835 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11151 8736
rect 10835 8671 11151 8672
rect 15780 8736 16096 8737
rect 15780 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16096 8736
rect 15780 8671 16096 8672
rect 20725 8736 21041 8737
rect 20725 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21041 8736
rect 20725 8671 21041 8672
rect 3418 8192 3734 8193
rect 3418 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3734 8192
rect 3418 8127 3734 8128
rect 8363 8192 8679 8193
rect 8363 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8679 8192
rect 8363 8127 8679 8128
rect 13308 8192 13624 8193
rect 13308 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13624 8192
rect 13308 8127 13624 8128
rect 18253 8192 18569 8193
rect 18253 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18569 8192
rect 18253 8127 18569 8128
rect 5890 7648 6206 7649
rect 5890 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6206 7648
rect 5890 7583 6206 7584
rect 10835 7648 11151 7649
rect 10835 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11151 7648
rect 10835 7583 11151 7584
rect 15780 7648 16096 7649
rect 15780 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16096 7648
rect 15780 7583 16096 7584
rect 20725 7648 21041 7649
rect 20725 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21041 7648
rect 20725 7583 21041 7584
rect 3418 7104 3734 7105
rect 3418 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3734 7104
rect 3418 7039 3734 7040
rect 8363 7104 8679 7105
rect 8363 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8679 7104
rect 8363 7039 8679 7040
rect 13308 7104 13624 7105
rect 13308 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13624 7104
rect 13308 7039 13624 7040
rect 18253 7104 18569 7105
rect 18253 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18569 7104
rect 18253 7039 18569 7040
rect 5890 6560 6206 6561
rect 5890 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6206 6560
rect 5890 6495 6206 6496
rect 10835 6560 11151 6561
rect 10835 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11151 6560
rect 10835 6495 11151 6496
rect 15780 6560 16096 6561
rect 15780 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16096 6560
rect 15780 6495 16096 6496
rect 20725 6560 21041 6561
rect 20725 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21041 6560
rect 20725 6495 21041 6496
rect 10225 6354 10291 6357
rect 16389 6354 16455 6357
rect 10225 6352 16455 6354
rect 10225 6296 10230 6352
rect 10286 6296 16394 6352
rect 16450 6296 16455 6352
rect 10225 6294 16455 6296
rect 10225 6291 10291 6294
rect 16389 6291 16455 6294
rect 14457 6082 14523 6085
rect 17861 6082 17927 6085
rect 14457 6080 17927 6082
rect 14457 6024 14462 6080
rect 14518 6024 17866 6080
rect 17922 6024 17927 6080
rect 14457 6022 17927 6024
rect 14457 6019 14523 6022
rect 17861 6019 17927 6022
rect 3418 6016 3734 6017
rect 3418 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3734 6016
rect 3418 5951 3734 5952
rect 8363 6016 8679 6017
rect 8363 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8679 6016
rect 8363 5951 8679 5952
rect 13308 6016 13624 6017
rect 13308 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13624 6016
rect 13308 5951 13624 5952
rect 18253 6016 18569 6017
rect 18253 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18569 6016
rect 18253 5951 18569 5952
rect 5890 5472 6206 5473
rect 5890 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6206 5472
rect 5890 5407 6206 5408
rect 10835 5472 11151 5473
rect 10835 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11151 5472
rect 10835 5407 11151 5408
rect 15780 5472 16096 5473
rect 15780 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16096 5472
rect 15780 5407 16096 5408
rect 20725 5472 21041 5473
rect 20725 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21041 5472
rect 20725 5407 21041 5408
rect 3418 4928 3734 4929
rect 3418 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3734 4928
rect 3418 4863 3734 4864
rect 8363 4928 8679 4929
rect 8363 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8679 4928
rect 8363 4863 8679 4864
rect 13308 4928 13624 4929
rect 13308 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13624 4928
rect 13308 4863 13624 4864
rect 18253 4928 18569 4929
rect 18253 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18569 4928
rect 18253 4863 18569 4864
rect 5890 4384 6206 4385
rect 5890 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6206 4384
rect 5890 4319 6206 4320
rect 10835 4384 11151 4385
rect 10835 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11151 4384
rect 10835 4319 11151 4320
rect 15780 4384 16096 4385
rect 15780 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16096 4384
rect 15780 4319 16096 4320
rect 20725 4384 21041 4385
rect 20725 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21041 4384
rect 20725 4319 21041 4320
rect 3418 3840 3734 3841
rect 3418 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3734 3840
rect 3418 3775 3734 3776
rect 8363 3840 8679 3841
rect 8363 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8679 3840
rect 8363 3775 8679 3776
rect 13308 3840 13624 3841
rect 13308 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13624 3840
rect 13308 3775 13624 3776
rect 18253 3840 18569 3841
rect 18253 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18569 3840
rect 18253 3775 18569 3776
rect 5890 3296 6206 3297
rect 5890 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6206 3296
rect 5890 3231 6206 3232
rect 10835 3296 11151 3297
rect 10835 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11151 3296
rect 10835 3231 11151 3232
rect 15780 3296 16096 3297
rect 15780 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16096 3296
rect 15780 3231 16096 3232
rect 20725 3296 21041 3297
rect 20725 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21041 3296
rect 20725 3231 21041 3232
rect 3418 2752 3734 2753
rect 3418 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3734 2752
rect 3418 2687 3734 2688
rect 8363 2752 8679 2753
rect 8363 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8679 2752
rect 8363 2687 8679 2688
rect 13308 2752 13624 2753
rect 13308 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13624 2752
rect 13308 2687 13624 2688
rect 18253 2752 18569 2753
rect 18253 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18569 2752
rect 18253 2687 18569 2688
rect 5890 2208 6206 2209
rect 5890 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6206 2208
rect 5890 2143 6206 2144
rect 10835 2208 11151 2209
rect 10835 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11151 2208
rect 10835 2143 11151 2144
rect 15780 2208 16096 2209
rect 15780 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16096 2208
rect 15780 2143 16096 2144
rect 20725 2208 21041 2209
rect 20725 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21041 2208
rect 20725 2143 21041 2144
<< via3 >>
rect 5896 19612 5960 19616
rect 5896 19556 5900 19612
rect 5900 19556 5956 19612
rect 5956 19556 5960 19612
rect 5896 19552 5960 19556
rect 5976 19612 6040 19616
rect 5976 19556 5980 19612
rect 5980 19556 6036 19612
rect 6036 19556 6040 19612
rect 5976 19552 6040 19556
rect 6056 19612 6120 19616
rect 6056 19556 6060 19612
rect 6060 19556 6116 19612
rect 6116 19556 6120 19612
rect 6056 19552 6120 19556
rect 6136 19612 6200 19616
rect 6136 19556 6140 19612
rect 6140 19556 6196 19612
rect 6196 19556 6200 19612
rect 6136 19552 6200 19556
rect 10841 19612 10905 19616
rect 10841 19556 10845 19612
rect 10845 19556 10901 19612
rect 10901 19556 10905 19612
rect 10841 19552 10905 19556
rect 10921 19612 10985 19616
rect 10921 19556 10925 19612
rect 10925 19556 10981 19612
rect 10981 19556 10985 19612
rect 10921 19552 10985 19556
rect 11001 19612 11065 19616
rect 11001 19556 11005 19612
rect 11005 19556 11061 19612
rect 11061 19556 11065 19612
rect 11001 19552 11065 19556
rect 11081 19612 11145 19616
rect 11081 19556 11085 19612
rect 11085 19556 11141 19612
rect 11141 19556 11145 19612
rect 11081 19552 11145 19556
rect 15786 19612 15850 19616
rect 15786 19556 15790 19612
rect 15790 19556 15846 19612
rect 15846 19556 15850 19612
rect 15786 19552 15850 19556
rect 15866 19612 15930 19616
rect 15866 19556 15870 19612
rect 15870 19556 15926 19612
rect 15926 19556 15930 19612
rect 15866 19552 15930 19556
rect 15946 19612 16010 19616
rect 15946 19556 15950 19612
rect 15950 19556 16006 19612
rect 16006 19556 16010 19612
rect 15946 19552 16010 19556
rect 16026 19612 16090 19616
rect 16026 19556 16030 19612
rect 16030 19556 16086 19612
rect 16086 19556 16090 19612
rect 16026 19552 16090 19556
rect 20731 19612 20795 19616
rect 20731 19556 20735 19612
rect 20735 19556 20791 19612
rect 20791 19556 20795 19612
rect 20731 19552 20795 19556
rect 20811 19612 20875 19616
rect 20811 19556 20815 19612
rect 20815 19556 20871 19612
rect 20871 19556 20875 19612
rect 20811 19552 20875 19556
rect 20891 19612 20955 19616
rect 20891 19556 20895 19612
rect 20895 19556 20951 19612
rect 20951 19556 20955 19612
rect 20891 19552 20955 19556
rect 20971 19612 21035 19616
rect 20971 19556 20975 19612
rect 20975 19556 21031 19612
rect 21031 19556 21035 19612
rect 20971 19552 21035 19556
rect 3424 19068 3488 19072
rect 3424 19012 3428 19068
rect 3428 19012 3484 19068
rect 3484 19012 3488 19068
rect 3424 19008 3488 19012
rect 3504 19068 3568 19072
rect 3504 19012 3508 19068
rect 3508 19012 3564 19068
rect 3564 19012 3568 19068
rect 3504 19008 3568 19012
rect 3584 19068 3648 19072
rect 3584 19012 3588 19068
rect 3588 19012 3644 19068
rect 3644 19012 3648 19068
rect 3584 19008 3648 19012
rect 3664 19068 3728 19072
rect 3664 19012 3668 19068
rect 3668 19012 3724 19068
rect 3724 19012 3728 19068
rect 3664 19008 3728 19012
rect 8369 19068 8433 19072
rect 8369 19012 8373 19068
rect 8373 19012 8429 19068
rect 8429 19012 8433 19068
rect 8369 19008 8433 19012
rect 8449 19068 8513 19072
rect 8449 19012 8453 19068
rect 8453 19012 8509 19068
rect 8509 19012 8513 19068
rect 8449 19008 8513 19012
rect 8529 19068 8593 19072
rect 8529 19012 8533 19068
rect 8533 19012 8589 19068
rect 8589 19012 8593 19068
rect 8529 19008 8593 19012
rect 8609 19068 8673 19072
rect 8609 19012 8613 19068
rect 8613 19012 8669 19068
rect 8669 19012 8673 19068
rect 8609 19008 8673 19012
rect 13314 19068 13378 19072
rect 13314 19012 13318 19068
rect 13318 19012 13374 19068
rect 13374 19012 13378 19068
rect 13314 19008 13378 19012
rect 13394 19068 13458 19072
rect 13394 19012 13398 19068
rect 13398 19012 13454 19068
rect 13454 19012 13458 19068
rect 13394 19008 13458 19012
rect 13474 19068 13538 19072
rect 13474 19012 13478 19068
rect 13478 19012 13534 19068
rect 13534 19012 13538 19068
rect 13474 19008 13538 19012
rect 13554 19068 13618 19072
rect 13554 19012 13558 19068
rect 13558 19012 13614 19068
rect 13614 19012 13618 19068
rect 13554 19008 13618 19012
rect 18259 19068 18323 19072
rect 18259 19012 18263 19068
rect 18263 19012 18319 19068
rect 18319 19012 18323 19068
rect 18259 19008 18323 19012
rect 18339 19068 18403 19072
rect 18339 19012 18343 19068
rect 18343 19012 18399 19068
rect 18399 19012 18403 19068
rect 18339 19008 18403 19012
rect 18419 19068 18483 19072
rect 18419 19012 18423 19068
rect 18423 19012 18479 19068
rect 18479 19012 18483 19068
rect 18419 19008 18483 19012
rect 18499 19068 18563 19072
rect 18499 19012 18503 19068
rect 18503 19012 18559 19068
rect 18559 19012 18563 19068
rect 18499 19008 18563 19012
rect 5896 18524 5960 18528
rect 5896 18468 5900 18524
rect 5900 18468 5956 18524
rect 5956 18468 5960 18524
rect 5896 18464 5960 18468
rect 5976 18524 6040 18528
rect 5976 18468 5980 18524
rect 5980 18468 6036 18524
rect 6036 18468 6040 18524
rect 5976 18464 6040 18468
rect 6056 18524 6120 18528
rect 6056 18468 6060 18524
rect 6060 18468 6116 18524
rect 6116 18468 6120 18524
rect 6056 18464 6120 18468
rect 6136 18524 6200 18528
rect 6136 18468 6140 18524
rect 6140 18468 6196 18524
rect 6196 18468 6200 18524
rect 6136 18464 6200 18468
rect 10841 18524 10905 18528
rect 10841 18468 10845 18524
rect 10845 18468 10901 18524
rect 10901 18468 10905 18524
rect 10841 18464 10905 18468
rect 10921 18524 10985 18528
rect 10921 18468 10925 18524
rect 10925 18468 10981 18524
rect 10981 18468 10985 18524
rect 10921 18464 10985 18468
rect 11001 18524 11065 18528
rect 11001 18468 11005 18524
rect 11005 18468 11061 18524
rect 11061 18468 11065 18524
rect 11001 18464 11065 18468
rect 11081 18524 11145 18528
rect 11081 18468 11085 18524
rect 11085 18468 11141 18524
rect 11141 18468 11145 18524
rect 11081 18464 11145 18468
rect 15786 18524 15850 18528
rect 15786 18468 15790 18524
rect 15790 18468 15846 18524
rect 15846 18468 15850 18524
rect 15786 18464 15850 18468
rect 15866 18524 15930 18528
rect 15866 18468 15870 18524
rect 15870 18468 15926 18524
rect 15926 18468 15930 18524
rect 15866 18464 15930 18468
rect 15946 18524 16010 18528
rect 15946 18468 15950 18524
rect 15950 18468 16006 18524
rect 16006 18468 16010 18524
rect 15946 18464 16010 18468
rect 16026 18524 16090 18528
rect 16026 18468 16030 18524
rect 16030 18468 16086 18524
rect 16086 18468 16090 18524
rect 16026 18464 16090 18468
rect 20731 18524 20795 18528
rect 20731 18468 20735 18524
rect 20735 18468 20791 18524
rect 20791 18468 20795 18524
rect 20731 18464 20795 18468
rect 20811 18524 20875 18528
rect 20811 18468 20815 18524
rect 20815 18468 20871 18524
rect 20871 18468 20875 18524
rect 20811 18464 20875 18468
rect 20891 18524 20955 18528
rect 20891 18468 20895 18524
rect 20895 18468 20951 18524
rect 20951 18468 20955 18524
rect 20891 18464 20955 18468
rect 20971 18524 21035 18528
rect 20971 18468 20975 18524
rect 20975 18468 21031 18524
rect 21031 18468 21035 18524
rect 20971 18464 21035 18468
rect 3424 17980 3488 17984
rect 3424 17924 3428 17980
rect 3428 17924 3484 17980
rect 3484 17924 3488 17980
rect 3424 17920 3488 17924
rect 3504 17980 3568 17984
rect 3504 17924 3508 17980
rect 3508 17924 3564 17980
rect 3564 17924 3568 17980
rect 3504 17920 3568 17924
rect 3584 17980 3648 17984
rect 3584 17924 3588 17980
rect 3588 17924 3644 17980
rect 3644 17924 3648 17980
rect 3584 17920 3648 17924
rect 3664 17980 3728 17984
rect 3664 17924 3668 17980
rect 3668 17924 3724 17980
rect 3724 17924 3728 17980
rect 3664 17920 3728 17924
rect 8369 17980 8433 17984
rect 8369 17924 8373 17980
rect 8373 17924 8429 17980
rect 8429 17924 8433 17980
rect 8369 17920 8433 17924
rect 8449 17980 8513 17984
rect 8449 17924 8453 17980
rect 8453 17924 8509 17980
rect 8509 17924 8513 17980
rect 8449 17920 8513 17924
rect 8529 17980 8593 17984
rect 8529 17924 8533 17980
rect 8533 17924 8589 17980
rect 8589 17924 8593 17980
rect 8529 17920 8593 17924
rect 8609 17980 8673 17984
rect 8609 17924 8613 17980
rect 8613 17924 8669 17980
rect 8669 17924 8673 17980
rect 8609 17920 8673 17924
rect 13314 17980 13378 17984
rect 13314 17924 13318 17980
rect 13318 17924 13374 17980
rect 13374 17924 13378 17980
rect 13314 17920 13378 17924
rect 13394 17980 13458 17984
rect 13394 17924 13398 17980
rect 13398 17924 13454 17980
rect 13454 17924 13458 17980
rect 13394 17920 13458 17924
rect 13474 17980 13538 17984
rect 13474 17924 13478 17980
rect 13478 17924 13534 17980
rect 13534 17924 13538 17980
rect 13474 17920 13538 17924
rect 13554 17980 13618 17984
rect 13554 17924 13558 17980
rect 13558 17924 13614 17980
rect 13614 17924 13618 17980
rect 13554 17920 13618 17924
rect 18259 17980 18323 17984
rect 18259 17924 18263 17980
rect 18263 17924 18319 17980
rect 18319 17924 18323 17980
rect 18259 17920 18323 17924
rect 18339 17980 18403 17984
rect 18339 17924 18343 17980
rect 18343 17924 18399 17980
rect 18399 17924 18403 17980
rect 18339 17920 18403 17924
rect 18419 17980 18483 17984
rect 18419 17924 18423 17980
rect 18423 17924 18479 17980
rect 18479 17924 18483 17980
rect 18419 17920 18483 17924
rect 18499 17980 18563 17984
rect 18499 17924 18503 17980
rect 18503 17924 18559 17980
rect 18559 17924 18563 17980
rect 18499 17920 18563 17924
rect 5896 17436 5960 17440
rect 5896 17380 5900 17436
rect 5900 17380 5956 17436
rect 5956 17380 5960 17436
rect 5896 17376 5960 17380
rect 5976 17436 6040 17440
rect 5976 17380 5980 17436
rect 5980 17380 6036 17436
rect 6036 17380 6040 17436
rect 5976 17376 6040 17380
rect 6056 17436 6120 17440
rect 6056 17380 6060 17436
rect 6060 17380 6116 17436
rect 6116 17380 6120 17436
rect 6056 17376 6120 17380
rect 6136 17436 6200 17440
rect 6136 17380 6140 17436
rect 6140 17380 6196 17436
rect 6196 17380 6200 17436
rect 6136 17376 6200 17380
rect 10841 17436 10905 17440
rect 10841 17380 10845 17436
rect 10845 17380 10901 17436
rect 10901 17380 10905 17436
rect 10841 17376 10905 17380
rect 10921 17436 10985 17440
rect 10921 17380 10925 17436
rect 10925 17380 10981 17436
rect 10981 17380 10985 17436
rect 10921 17376 10985 17380
rect 11001 17436 11065 17440
rect 11001 17380 11005 17436
rect 11005 17380 11061 17436
rect 11061 17380 11065 17436
rect 11001 17376 11065 17380
rect 11081 17436 11145 17440
rect 11081 17380 11085 17436
rect 11085 17380 11141 17436
rect 11141 17380 11145 17436
rect 11081 17376 11145 17380
rect 15786 17436 15850 17440
rect 15786 17380 15790 17436
rect 15790 17380 15846 17436
rect 15846 17380 15850 17436
rect 15786 17376 15850 17380
rect 15866 17436 15930 17440
rect 15866 17380 15870 17436
rect 15870 17380 15926 17436
rect 15926 17380 15930 17436
rect 15866 17376 15930 17380
rect 15946 17436 16010 17440
rect 15946 17380 15950 17436
rect 15950 17380 16006 17436
rect 16006 17380 16010 17436
rect 15946 17376 16010 17380
rect 16026 17436 16090 17440
rect 16026 17380 16030 17436
rect 16030 17380 16086 17436
rect 16086 17380 16090 17436
rect 16026 17376 16090 17380
rect 20731 17436 20795 17440
rect 20731 17380 20735 17436
rect 20735 17380 20791 17436
rect 20791 17380 20795 17436
rect 20731 17376 20795 17380
rect 20811 17436 20875 17440
rect 20811 17380 20815 17436
rect 20815 17380 20871 17436
rect 20871 17380 20875 17436
rect 20811 17376 20875 17380
rect 20891 17436 20955 17440
rect 20891 17380 20895 17436
rect 20895 17380 20951 17436
rect 20951 17380 20955 17436
rect 20891 17376 20955 17380
rect 20971 17436 21035 17440
rect 20971 17380 20975 17436
rect 20975 17380 21031 17436
rect 21031 17380 21035 17436
rect 20971 17376 21035 17380
rect 3424 16892 3488 16896
rect 3424 16836 3428 16892
rect 3428 16836 3484 16892
rect 3484 16836 3488 16892
rect 3424 16832 3488 16836
rect 3504 16892 3568 16896
rect 3504 16836 3508 16892
rect 3508 16836 3564 16892
rect 3564 16836 3568 16892
rect 3504 16832 3568 16836
rect 3584 16892 3648 16896
rect 3584 16836 3588 16892
rect 3588 16836 3644 16892
rect 3644 16836 3648 16892
rect 3584 16832 3648 16836
rect 3664 16892 3728 16896
rect 3664 16836 3668 16892
rect 3668 16836 3724 16892
rect 3724 16836 3728 16892
rect 3664 16832 3728 16836
rect 8369 16892 8433 16896
rect 8369 16836 8373 16892
rect 8373 16836 8429 16892
rect 8429 16836 8433 16892
rect 8369 16832 8433 16836
rect 8449 16892 8513 16896
rect 8449 16836 8453 16892
rect 8453 16836 8509 16892
rect 8509 16836 8513 16892
rect 8449 16832 8513 16836
rect 8529 16892 8593 16896
rect 8529 16836 8533 16892
rect 8533 16836 8589 16892
rect 8589 16836 8593 16892
rect 8529 16832 8593 16836
rect 8609 16892 8673 16896
rect 8609 16836 8613 16892
rect 8613 16836 8669 16892
rect 8669 16836 8673 16892
rect 8609 16832 8673 16836
rect 13314 16892 13378 16896
rect 13314 16836 13318 16892
rect 13318 16836 13374 16892
rect 13374 16836 13378 16892
rect 13314 16832 13378 16836
rect 13394 16892 13458 16896
rect 13394 16836 13398 16892
rect 13398 16836 13454 16892
rect 13454 16836 13458 16892
rect 13394 16832 13458 16836
rect 13474 16892 13538 16896
rect 13474 16836 13478 16892
rect 13478 16836 13534 16892
rect 13534 16836 13538 16892
rect 13474 16832 13538 16836
rect 13554 16892 13618 16896
rect 13554 16836 13558 16892
rect 13558 16836 13614 16892
rect 13614 16836 13618 16892
rect 13554 16832 13618 16836
rect 18259 16892 18323 16896
rect 18259 16836 18263 16892
rect 18263 16836 18319 16892
rect 18319 16836 18323 16892
rect 18259 16832 18323 16836
rect 18339 16892 18403 16896
rect 18339 16836 18343 16892
rect 18343 16836 18399 16892
rect 18399 16836 18403 16892
rect 18339 16832 18403 16836
rect 18419 16892 18483 16896
rect 18419 16836 18423 16892
rect 18423 16836 18479 16892
rect 18479 16836 18483 16892
rect 18419 16832 18483 16836
rect 18499 16892 18563 16896
rect 18499 16836 18503 16892
rect 18503 16836 18559 16892
rect 18559 16836 18563 16892
rect 18499 16832 18563 16836
rect 5896 16348 5960 16352
rect 5896 16292 5900 16348
rect 5900 16292 5956 16348
rect 5956 16292 5960 16348
rect 5896 16288 5960 16292
rect 5976 16348 6040 16352
rect 5976 16292 5980 16348
rect 5980 16292 6036 16348
rect 6036 16292 6040 16348
rect 5976 16288 6040 16292
rect 6056 16348 6120 16352
rect 6056 16292 6060 16348
rect 6060 16292 6116 16348
rect 6116 16292 6120 16348
rect 6056 16288 6120 16292
rect 6136 16348 6200 16352
rect 6136 16292 6140 16348
rect 6140 16292 6196 16348
rect 6196 16292 6200 16348
rect 6136 16288 6200 16292
rect 10841 16348 10905 16352
rect 10841 16292 10845 16348
rect 10845 16292 10901 16348
rect 10901 16292 10905 16348
rect 10841 16288 10905 16292
rect 10921 16348 10985 16352
rect 10921 16292 10925 16348
rect 10925 16292 10981 16348
rect 10981 16292 10985 16348
rect 10921 16288 10985 16292
rect 11001 16348 11065 16352
rect 11001 16292 11005 16348
rect 11005 16292 11061 16348
rect 11061 16292 11065 16348
rect 11001 16288 11065 16292
rect 11081 16348 11145 16352
rect 11081 16292 11085 16348
rect 11085 16292 11141 16348
rect 11141 16292 11145 16348
rect 11081 16288 11145 16292
rect 15786 16348 15850 16352
rect 15786 16292 15790 16348
rect 15790 16292 15846 16348
rect 15846 16292 15850 16348
rect 15786 16288 15850 16292
rect 15866 16348 15930 16352
rect 15866 16292 15870 16348
rect 15870 16292 15926 16348
rect 15926 16292 15930 16348
rect 15866 16288 15930 16292
rect 15946 16348 16010 16352
rect 15946 16292 15950 16348
rect 15950 16292 16006 16348
rect 16006 16292 16010 16348
rect 15946 16288 16010 16292
rect 16026 16348 16090 16352
rect 16026 16292 16030 16348
rect 16030 16292 16086 16348
rect 16086 16292 16090 16348
rect 16026 16288 16090 16292
rect 20731 16348 20795 16352
rect 20731 16292 20735 16348
rect 20735 16292 20791 16348
rect 20791 16292 20795 16348
rect 20731 16288 20795 16292
rect 20811 16348 20875 16352
rect 20811 16292 20815 16348
rect 20815 16292 20871 16348
rect 20871 16292 20875 16348
rect 20811 16288 20875 16292
rect 20891 16348 20955 16352
rect 20891 16292 20895 16348
rect 20895 16292 20951 16348
rect 20951 16292 20955 16348
rect 20891 16288 20955 16292
rect 20971 16348 21035 16352
rect 20971 16292 20975 16348
rect 20975 16292 21031 16348
rect 21031 16292 21035 16348
rect 20971 16288 21035 16292
rect 3424 15804 3488 15808
rect 3424 15748 3428 15804
rect 3428 15748 3484 15804
rect 3484 15748 3488 15804
rect 3424 15744 3488 15748
rect 3504 15804 3568 15808
rect 3504 15748 3508 15804
rect 3508 15748 3564 15804
rect 3564 15748 3568 15804
rect 3504 15744 3568 15748
rect 3584 15804 3648 15808
rect 3584 15748 3588 15804
rect 3588 15748 3644 15804
rect 3644 15748 3648 15804
rect 3584 15744 3648 15748
rect 3664 15804 3728 15808
rect 3664 15748 3668 15804
rect 3668 15748 3724 15804
rect 3724 15748 3728 15804
rect 3664 15744 3728 15748
rect 8369 15804 8433 15808
rect 8369 15748 8373 15804
rect 8373 15748 8429 15804
rect 8429 15748 8433 15804
rect 8369 15744 8433 15748
rect 8449 15804 8513 15808
rect 8449 15748 8453 15804
rect 8453 15748 8509 15804
rect 8509 15748 8513 15804
rect 8449 15744 8513 15748
rect 8529 15804 8593 15808
rect 8529 15748 8533 15804
rect 8533 15748 8589 15804
rect 8589 15748 8593 15804
rect 8529 15744 8593 15748
rect 8609 15804 8673 15808
rect 8609 15748 8613 15804
rect 8613 15748 8669 15804
rect 8669 15748 8673 15804
rect 8609 15744 8673 15748
rect 13314 15804 13378 15808
rect 13314 15748 13318 15804
rect 13318 15748 13374 15804
rect 13374 15748 13378 15804
rect 13314 15744 13378 15748
rect 13394 15804 13458 15808
rect 13394 15748 13398 15804
rect 13398 15748 13454 15804
rect 13454 15748 13458 15804
rect 13394 15744 13458 15748
rect 13474 15804 13538 15808
rect 13474 15748 13478 15804
rect 13478 15748 13534 15804
rect 13534 15748 13538 15804
rect 13474 15744 13538 15748
rect 13554 15804 13618 15808
rect 13554 15748 13558 15804
rect 13558 15748 13614 15804
rect 13614 15748 13618 15804
rect 13554 15744 13618 15748
rect 18259 15804 18323 15808
rect 18259 15748 18263 15804
rect 18263 15748 18319 15804
rect 18319 15748 18323 15804
rect 18259 15744 18323 15748
rect 18339 15804 18403 15808
rect 18339 15748 18343 15804
rect 18343 15748 18399 15804
rect 18399 15748 18403 15804
rect 18339 15744 18403 15748
rect 18419 15804 18483 15808
rect 18419 15748 18423 15804
rect 18423 15748 18479 15804
rect 18479 15748 18483 15804
rect 18419 15744 18483 15748
rect 18499 15804 18563 15808
rect 18499 15748 18503 15804
rect 18503 15748 18559 15804
rect 18559 15748 18563 15804
rect 18499 15744 18563 15748
rect 5896 15260 5960 15264
rect 5896 15204 5900 15260
rect 5900 15204 5956 15260
rect 5956 15204 5960 15260
rect 5896 15200 5960 15204
rect 5976 15260 6040 15264
rect 5976 15204 5980 15260
rect 5980 15204 6036 15260
rect 6036 15204 6040 15260
rect 5976 15200 6040 15204
rect 6056 15260 6120 15264
rect 6056 15204 6060 15260
rect 6060 15204 6116 15260
rect 6116 15204 6120 15260
rect 6056 15200 6120 15204
rect 6136 15260 6200 15264
rect 6136 15204 6140 15260
rect 6140 15204 6196 15260
rect 6196 15204 6200 15260
rect 6136 15200 6200 15204
rect 10841 15260 10905 15264
rect 10841 15204 10845 15260
rect 10845 15204 10901 15260
rect 10901 15204 10905 15260
rect 10841 15200 10905 15204
rect 10921 15260 10985 15264
rect 10921 15204 10925 15260
rect 10925 15204 10981 15260
rect 10981 15204 10985 15260
rect 10921 15200 10985 15204
rect 11001 15260 11065 15264
rect 11001 15204 11005 15260
rect 11005 15204 11061 15260
rect 11061 15204 11065 15260
rect 11001 15200 11065 15204
rect 11081 15260 11145 15264
rect 11081 15204 11085 15260
rect 11085 15204 11141 15260
rect 11141 15204 11145 15260
rect 11081 15200 11145 15204
rect 15786 15260 15850 15264
rect 15786 15204 15790 15260
rect 15790 15204 15846 15260
rect 15846 15204 15850 15260
rect 15786 15200 15850 15204
rect 15866 15260 15930 15264
rect 15866 15204 15870 15260
rect 15870 15204 15926 15260
rect 15926 15204 15930 15260
rect 15866 15200 15930 15204
rect 15946 15260 16010 15264
rect 15946 15204 15950 15260
rect 15950 15204 16006 15260
rect 16006 15204 16010 15260
rect 15946 15200 16010 15204
rect 16026 15260 16090 15264
rect 16026 15204 16030 15260
rect 16030 15204 16086 15260
rect 16086 15204 16090 15260
rect 16026 15200 16090 15204
rect 20731 15260 20795 15264
rect 20731 15204 20735 15260
rect 20735 15204 20791 15260
rect 20791 15204 20795 15260
rect 20731 15200 20795 15204
rect 20811 15260 20875 15264
rect 20811 15204 20815 15260
rect 20815 15204 20871 15260
rect 20871 15204 20875 15260
rect 20811 15200 20875 15204
rect 20891 15260 20955 15264
rect 20891 15204 20895 15260
rect 20895 15204 20951 15260
rect 20951 15204 20955 15260
rect 20891 15200 20955 15204
rect 20971 15260 21035 15264
rect 20971 15204 20975 15260
rect 20975 15204 21031 15260
rect 21031 15204 21035 15260
rect 20971 15200 21035 15204
rect 3424 14716 3488 14720
rect 3424 14660 3428 14716
rect 3428 14660 3484 14716
rect 3484 14660 3488 14716
rect 3424 14656 3488 14660
rect 3504 14716 3568 14720
rect 3504 14660 3508 14716
rect 3508 14660 3564 14716
rect 3564 14660 3568 14716
rect 3504 14656 3568 14660
rect 3584 14716 3648 14720
rect 3584 14660 3588 14716
rect 3588 14660 3644 14716
rect 3644 14660 3648 14716
rect 3584 14656 3648 14660
rect 3664 14716 3728 14720
rect 3664 14660 3668 14716
rect 3668 14660 3724 14716
rect 3724 14660 3728 14716
rect 3664 14656 3728 14660
rect 8369 14716 8433 14720
rect 8369 14660 8373 14716
rect 8373 14660 8429 14716
rect 8429 14660 8433 14716
rect 8369 14656 8433 14660
rect 8449 14716 8513 14720
rect 8449 14660 8453 14716
rect 8453 14660 8509 14716
rect 8509 14660 8513 14716
rect 8449 14656 8513 14660
rect 8529 14716 8593 14720
rect 8529 14660 8533 14716
rect 8533 14660 8589 14716
rect 8589 14660 8593 14716
rect 8529 14656 8593 14660
rect 8609 14716 8673 14720
rect 8609 14660 8613 14716
rect 8613 14660 8669 14716
rect 8669 14660 8673 14716
rect 8609 14656 8673 14660
rect 13314 14716 13378 14720
rect 13314 14660 13318 14716
rect 13318 14660 13374 14716
rect 13374 14660 13378 14716
rect 13314 14656 13378 14660
rect 13394 14716 13458 14720
rect 13394 14660 13398 14716
rect 13398 14660 13454 14716
rect 13454 14660 13458 14716
rect 13394 14656 13458 14660
rect 13474 14716 13538 14720
rect 13474 14660 13478 14716
rect 13478 14660 13534 14716
rect 13534 14660 13538 14716
rect 13474 14656 13538 14660
rect 13554 14716 13618 14720
rect 13554 14660 13558 14716
rect 13558 14660 13614 14716
rect 13614 14660 13618 14716
rect 13554 14656 13618 14660
rect 18259 14716 18323 14720
rect 18259 14660 18263 14716
rect 18263 14660 18319 14716
rect 18319 14660 18323 14716
rect 18259 14656 18323 14660
rect 18339 14716 18403 14720
rect 18339 14660 18343 14716
rect 18343 14660 18399 14716
rect 18399 14660 18403 14716
rect 18339 14656 18403 14660
rect 18419 14716 18483 14720
rect 18419 14660 18423 14716
rect 18423 14660 18479 14716
rect 18479 14660 18483 14716
rect 18419 14656 18483 14660
rect 18499 14716 18563 14720
rect 18499 14660 18503 14716
rect 18503 14660 18559 14716
rect 18559 14660 18563 14716
rect 18499 14656 18563 14660
rect 5896 14172 5960 14176
rect 5896 14116 5900 14172
rect 5900 14116 5956 14172
rect 5956 14116 5960 14172
rect 5896 14112 5960 14116
rect 5976 14172 6040 14176
rect 5976 14116 5980 14172
rect 5980 14116 6036 14172
rect 6036 14116 6040 14172
rect 5976 14112 6040 14116
rect 6056 14172 6120 14176
rect 6056 14116 6060 14172
rect 6060 14116 6116 14172
rect 6116 14116 6120 14172
rect 6056 14112 6120 14116
rect 6136 14172 6200 14176
rect 6136 14116 6140 14172
rect 6140 14116 6196 14172
rect 6196 14116 6200 14172
rect 6136 14112 6200 14116
rect 10841 14172 10905 14176
rect 10841 14116 10845 14172
rect 10845 14116 10901 14172
rect 10901 14116 10905 14172
rect 10841 14112 10905 14116
rect 10921 14172 10985 14176
rect 10921 14116 10925 14172
rect 10925 14116 10981 14172
rect 10981 14116 10985 14172
rect 10921 14112 10985 14116
rect 11001 14172 11065 14176
rect 11001 14116 11005 14172
rect 11005 14116 11061 14172
rect 11061 14116 11065 14172
rect 11001 14112 11065 14116
rect 11081 14172 11145 14176
rect 11081 14116 11085 14172
rect 11085 14116 11141 14172
rect 11141 14116 11145 14172
rect 11081 14112 11145 14116
rect 15786 14172 15850 14176
rect 15786 14116 15790 14172
rect 15790 14116 15846 14172
rect 15846 14116 15850 14172
rect 15786 14112 15850 14116
rect 15866 14172 15930 14176
rect 15866 14116 15870 14172
rect 15870 14116 15926 14172
rect 15926 14116 15930 14172
rect 15866 14112 15930 14116
rect 15946 14172 16010 14176
rect 15946 14116 15950 14172
rect 15950 14116 16006 14172
rect 16006 14116 16010 14172
rect 15946 14112 16010 14116
rect 16026 14172 16090 14176
rect 16026 14116 16030 14172
rect 16030 14116 16086 14172
rect 16086 14116 16090 14172
rect 16026 14112 16090 14116
rect 20731 14172 20795 14176
rect 20731 14116 20735 14172
rect 20735 14116 20791 14172
rect 20791 14116 20795 14172
rect 20731 14112 20795 14116
rect 20811 14172 20875 14176
rect 20811 14116 20815 14172
rect 20815 14116 20871 14172
rect 20871 14116 20875 14172
rect 20811 14112 20875 14116
rect 20891 14172 20955 14176
rect 20891 14116 20895 14172
rect 20895 14116 20951 14172
rect 20951 14116 20955 14172
rect 20891 14112 20955 14116
rect 20971 14172 21035 14176
rect 20971 14116 20975 14172
rect 20975 14116 21031 14172
rect 21031 14116 21035 14172
rect 20971 14112 21035 14116
rect 3424 13628 3488 13632
rect 3424 13572 3428 13628
rect 3428 13572 3484 13628
rect 3484 13572 3488 13628
rect 3424 13568 3488 13572
rect 3504 13628 3568 13632
rect 3504 13572 3508 13628
rect 3508 13572 3564 13628
rect 3564 13572 3568 13628
rect 3504 13568 3568 13572
rect 3584 13628 3648 13632
rect 3584 13572 3588 13628
rect 3588 13572 3644 13628
rect 3644 13572 3648 13628
rect 3584 13568 3648 13572
rect 3664 13628 3728 13632
rect 3664 13572 3668 13628
rect 3668 13572 3724 13628
rect 3724 13572 3728 13628
rect 3664 13568 3728 13572
rect 8369 13628 8433 13632
rect 8369 13572 8373 13628
rect 8373 13572 8429 13628
rect 8429 13572 8433 13628
rect 8369 13568 8433 13572
rect 8449 13628 8513 13632
rect 8449 13572 8453 13628
rect 8453 13572 8509 13628
rect 8509 13572 8513 13628
rect 8449 13568 8513 13572
rect 8529 13628 8593 13632
rect 8529 13572 8533 13628
rect 8533 13572 8589 13628
rect 8589 13572 8593 13628
rect 8529 13568 8593 13572
rect 8609 13628 8673 13632
rect 8609 13572 8613 13628
rect 8613 13572 8669 13628
rect 8669 13572 8673 13628
rect 8609 13568 8673 13572
rect 13314 13628 13378 13632
rect 13314 13572 13318 13628
rect 13318 13572 13374 13628
rect 13374 13572 13378 13628
rect 13314 13568 13378 13572
rect 13394 13628 13458 13632
rect 13394 13572 13398 13628
rect 13398 13572 13454 13628
rect 13454 13572 13458 13628
rect 13394 13568 13458 13572
rect 13474 13628 13538 13632
rect 13474 13572 13478 13628
rect 13478 13572 13534 13628
rect 13534 13572 13538 13628
rect 13474 13568 13538 13572
rect 13554 13628 13618 13632
rect 13554 13572 13558 13628
rect 13558 13572 13614 13628
rect 13614 13572 13618 13628
rect 13554 13568 13618 13572
rect 18259 13628 18323 13632
rect 18259 13572 18263 13628
rect 18263 13572 18319 13628
rect 18319 13572 18323 13628
rect 18259 13568 18323 13572
rect 18339 13628 18403 13632
rect 18339 13572 18343 13628
rect 18343 13572 18399 13628
rect 18399 13572 18403 13628
rect 18339 13568 18403 13572
rect 18419 13628 18483 13632
rect 18419 13572 18423 13628
rect 18423 13572 18479 13628
rect 18479 13572 18483 13628
rect 18419 13568 18483 13572
rect 18499 13628 18563 13632
rect 18499 13572 18503 13628
rect 18503 13572 18559 13628
rect 18559 13572 18563 13628
rect 18499 13568 18563 13572
rect 5896 13084 5960 13088
rect 5896 13028 5900 13084
rect 5900 13028 5956 13084
rect 5956 13028 5960 13084
rect 5896 13024 5960 13028
rect 5976 13084 6040 13088
rect 5976 13028 5980 13084
rect 5980 13028 6036 13084
rect 6036 13028 6040 13084
rect 5976 13024 6040 13028
rect 6056 13084 6120 13088
rect 6056 13028 6060 13084
rect 6060 13028 6116 13084
rect 6116 13028 6120 13084
rect 6056 13024 6120 13028
rect 6136 13084 6200 13088
rect 6136 13028 6140 13084
rect 6140 13028 6196 13084
rect 6196 13028 6200 13084
rect 6136 13024 6200 13028
rect 10841 13084 10905 13088
rect 10841 13028 10845 13084
rect 10845 13028 10901 13084
rect 10901 13028 10905 13084
rect 10841 13024 10905 13028
rect 10921 13084 10985 13088
rect 10921 13028 10925 13084
rect 10925 13028 10981 13084
rect 10981 13028 10985 13084
rect 10921 13024 10985 13028
rect 11001 13084 11065 13088
rect 11001 13028 11005 13084
rect 11005 13028 11061 13084
rect 11061 13028 11065 13084
rect 11001 13024 11065 13028
rect 11081 13084 11145 13088
rect 11081 13028 11085 13084
rect 11085 13028 11141 13084
rect 11141 13028 11145 13084
rect 11081 13024 11145 13028
rect 15786 13084 15850 13088
rect 15786 13028 15790 13084
rect 15790 13028 15846 13084
rect 15846 13028 15850 13084
rect 15786 13024 15850 13028
rect 15866 13084 15930 13088
rect 15866 13028 15870 13084
rect 15870 13028 15926 13084
rect 15926 13028 15930 13084
rect 15866 13024 15930 13028
rect 15946 13084 16010 13088
rect 15946 13028 15950 13084
rect 15950 13028 16006 13084
rect 16006 13028 16010 13084
rect 15946 13024 16010 13028
rect 16026 13084 16090 13088
rect 16026 13028 16030 13084
rect 16030 13028 16086 13084
rect 16086 13028 16090 13084
rect 16026 13024 16090 13028
rect 20731 13084 20795 13088
rect 20731 13028 20735 13084
rect 20735 13028 20791 13084
rect 20791 13028 20795 13084
rect 20731 13024 20795 13028
rect 20811 13084 20875 13088
rect 20811 13028 20815 13084
rect 20815 13028 20871 13084
rect 20871 13028 20875 13084
rect 20811 13024 20875 13028
rect 20891 13084 20955 13088
rect 20891 13028 20895 13084
rect 20895 13028 20951 13084
rect 20951 13028 20955 13084
rect 20891 13024 20955 13028
rect 20971 13084 21035 13088
rect 20971 13028 20975 13084
rect 20975 13028 21031 13084
rect 21031 13028 21035 13084
rect 20971 13024 21035 13028
rect 3424 12540 3488 12544
rect 3424 12484 3428 12540
rect 3428 12484 3484 12540
rect 3484 12484 3488 12540
rect 3424 12480 3488 12484
rect 3504 12540 3568 12544
rect 3504 12484 3508 12540
rect 3508 12484 3564 12540
rect 3564 12484 3568 12540
rect 3504 12480 3568 12484
rect 3584 12540 3648 12544
rect 3584 12484 3588 12540
rect 3588 12484 3644 12540
rect 3644 12484 3648 12540
rect 3584 12480 3648 12484
rect 3664 12540 3728 12544
rect 3664 12484 3668 12540
rect 3668 12484 3724 12540
rect 3724 12484 3728 12540
rect 3664 12480 3728 12484
rect 8369 12540 8433 12544
rect 8369 12484 8373 12540
rect 8373 12484 8429 12540
rect 8429 12484 8433 12540
rect 8369 12480 8433 12484
rect 8449 12540 8513 12544
rect 8449 12484 8453 12540
rect 8453 12484 8509 12540
rect 8509 12484 8513 12540
rect 8449 12480 8513 12484
rect 8529 12540 8593 12544
rect 8529 12484 8533 12540
rect 8533 12484 8589 12540
rect 8589 12484 8593 12540
rect 8529 12480 8593 12484
rect 8609 12540 8673 12544
rect 8609 12484 8613 12540
rect 8613 12484 8669 12540
rect 8669 12484 8673 12540
rect 8609 12480 8673 12484
rect 13314 12540 13378 12544
rect 13314 12484 13318 12540
rect 13318 12484 13374 12540
rect 13374 12484 13378 12540
rect 13314 12480 13378 12484
rect 13394 12540 13458 12544
rect 13394 12484 13398 12540
rect 13398 12484 13454 12540
rect 13454 12484 13458 12540
rect 13394 12480 13458 12484
rect 13474 12540 13538 12544
rect 13474 12484 13478 12540
rect 13478 12484 13534 12540
rect 13534 12484 13538 12540
rect 13474 12480 13538 12484
rect 13554 12540 13618 12544
rect 13554 12484 13558 12540
rect 13558 12484 13614 12540
rect 13614 12484 13618 12540
rect 13554 12480 13618 12484
rect 18259 12540 18323 12544
rect 18259 12484 18263 12540
rect 18263 12484 18319 12540
rect 18319 12484 18323 12540
rect 18259 12480 18323 12484
rect 18339 12540 18403 12544
rect 18339 12484 18343 12540
rect 18343 12484 18399 12540
rect 18399 12484 18403 12540
rect 18339 12480 18403 12484
rect 18419 12540 18483 12544
rect 18419 12484 18423 12540
rect 18423 12484 18479 12540
rect 18479 12484 18483 12540
rect 18419 12480 18483 12484
rect 18499 12540 18563 12544
rect 18499 12484 18503 12540
rect 18503 12484 18559 12540
rect 18559 12484 18563 12540
rect 18499 12480 18563 12484
rect 5896 11996 5960 12000
rect 5896 11940 5900 11996
rect 5900 11940 5956 11996
rect 5956 11940 5960 11996
rect 5896 11936 5960 11940
rect 5976 11996 6040 12000
rect 5976 11940 5980 11996
rect 5980 11940 6036 11996
rect 6036 11940 6040 11996
rect 5976 11936 6040 11940
rect 6056 11996 6120 12000
rect 6056 11940 6060 11996
rect 6060 11940 6116 11996
rect 6116 11940 6120 11996
rect 6056 11936 6120 11940
rect 6136 11996 6200 12000
rect 6136 11940 6140 11996
rect 6140 11940 6196 11996
rect 6196 11940 6200 11996
rect 6136 11936 6200 11940
rect 10841 11996 10905 12000
rect 10841 11940 10845 11996
rect 10845 11940 10901 11996
rect 10901 11940 10905 11996
rect 10841 11936 10905 11940
rect 10921 11996 10985 12000
rect 10921 11940 10925 11996
rect 10925 11940 10981 11996
rect 10981 11940 10985 11996
rect 10921 11936 10985 11940
rect 11001 11996 11065 12000
rect 11001 11940 11005 11996
rect 11005 11940 11061 11996
rect 11061 11940 11065 11996
rect 11001 11936 11065 11940
rect 11081 11996 11145 12000
rect 11081 11940 11085 11996
rect 11085 11940 11141 11996
rect 11141 11940 11145 11996
rect 11081 11936 11145 11940
rect 15786 11996 15850 12000
rect 15786 11940 15790 11996
rect 15790 11940 15846 11996
rect 15846 11940 15850 11996
rect 15786 11936 15850 11940
rect 15866 11996 15930 12000
rect 15866 11940 15870 11996
rect 15870 11940 15926 11996
rect 15926 11940 15930 11996
rect 15866 11936 15930 11940
rect 15946 11996 16010 12000
rect 15946 11940 15950 11996
rect 15950 11940 16006 11996
rect 16006 11940 16010 11996
rect 15946 11936 16010 11940
rect 16026 11996 16090 12000
rect 16026 11940 16030 11996
rect 16030 11940 16086 11996
rect 16086 11940 16090 11996
rect 16026 11936 16090 11940
rect 20731 11996 20795 12000
rect 20731 11940 20735 11996
rect 20735 11940 20791 11996
rect 20791 11940 20795 11996
rect 20731 11936 20795 11940
rect 20811 11996 20875 12000
rect 20811 11940 20815 11996
rect 20815 11940 20871 11996
rect 20871 11940 20875 11996
rect 20811 11936 20875 11940
rect 20891 11996 20955 12000
rect 20891 11940 20895 11996
rect 20895 11940 20951 11996
rect 20951 11940 20955 11996
rect 20891 11936 20955 11940
rect 20971 11996 21035 12000
rect 20971 11940 20975 11996
rect 20975 11940 21031 11996
rect 21031 11940 21035 11996
rect 20971 11936 21035 11940
rect 3424 11452 3488 11456
rect 3424 11396 3428 11452
rect 3428 11396 3484 11452
rect 3484 11396 3488 11452
rect 3424 11392 3488 11396
rect 3504 11452 3568 11456
rect 3504 11396 3508 11452
rect 3508 11396 3564 11452
rect 3564 11396 3568 11452
rect 3504 11392 3568 11396
rect 3584 11452 3648 11456
rect 3584 11396 3588 11452
rect 3588 11396 3644 11452
rect 3644 11396 3648 11452
rect 3584 11392 3648 11396
rect 3664 11452 3728 11456
rect 3664 11396 3668 11452
rect 3668 11396 3724 11452
rect 3724 11396 3728 11452
rect 3664 11392 3728 11396
rect 8369 11452 8433 11456
rect 8369 11396 8373 11452
rect 8373 11396 8429 11452
rect 8429 11396 8433 11452
rect 8369 11392 8433 11396
rect 8449 11452 8513 11456
rect 8449 11396 8453 11452
rect 8453 11396 8509 11452
rect 8509 11396 8513 11452
rect 8449 11392 8513 11396
rect 8529 11452 8593 11456
rect 8529 11396 8533 11452
rect 8533 11396 8589 11452
rect 8589 11396 8593 11452
rect 8529 11392 8593 11396
rect 8609 11452 8673 11456
rect 8609 11396 8613 11452
rect 8613 11396 8669 11452
rect 8669 11396 8673 11452
rect 8609 11392 8673 11396
rect 13314 11452 13378 11456
rect 13314 11396 13318 11452
rect 13318 11396 13374 11452
rect 13374 11396 13378 11452
rect 13314 11392 13378 11396
rect 13394 11452 13458 11456
rect 13394 11396 13398 11452
rect 13398 11396 13454 11452
rect 13454 11396 13458 11452
rect 13394 11392 13458 11396
rect 13474 11452 13538 11456
rect 13474 11396 13478 11452
rect 13478 11396 13534 11452
rect 13534 11396 13538 11452
rect 13474 11392 13538 11396
rect 13554 11452 13618 11456
rect 13554 11396 13558 11452
rect 13558 11396 13614 11452
rect 13614 11396 13618 11452
rect 13554 11392 13618 11396
rect 18259 11452 18323 11456
rect 18259 11396 18263 11452
rect 18263 11396 18319 11452
rect 18319 11396 18323 11452
rect 18259 11392 18323 11396
rect 18339 11452 18403 11456
rect 18339 11396 18343 11452
rect 18343 11396 18399 11452
rect 18399 11396 18403 11452
rect 18339 11392 18403 11396
rect 18419 11452 18483 11456
rect 18419 11396 18423 11452
rect 18423 11396 18479 11452
rect 18479 11396 18483 11452
rect 18419 11392 18483 11396
rect 18499 11452 18563 11456
rect 18499 11396 18503 11452
rect 18503 11396 18559 11452
rect 18559 11396 18563 11452
rect 18499 11392 18563 11396
rect 5896 10908 5960 10912
rect 5896 10852 5900 10908
rect 5900 10852 5956 10908
rect 5956 10852 5960 10908
rect 5896 10848 5960 10852
rect 5976 10908 6040 10912
rect 5976 10852 5980 10908
rect 5980 10852 6036 10908
rect 6036 10852 6040 10908
rect 5976 10848 6040 10852
rect 6056 10908 6120 10912
rect 6056 10852 6060 10908
rect 6060 10852 6116 10908
rect 6116 10852 6120 10908
rect 6056 10848 6120 10852
rect 6136 10908 6200 10912
rect 6136 10852 6140 10908
rect 6140 10852 6196 10908
rect 6196 10852 6200 10908
rect 6136 10848 6200 10852
rect 10841 10908 10905 10912
rect 10841 10852 10845 10908
rect 10845 10852 10901 10908
rect 10901 10852 10905 10908
rect 10841 10848 10905 10852
rect 10921 10908 10985 10912
rect 10921 10852 10925 10908
rect 10925 10852 10981 10908
rect 10981 10852 10985 10908
rect 10921 10848 10985 10852
rect 11001 10908 11065 10912
rect 11001 10852 11005 10908
rect 11005 10852 11061 10908
rect 11061 10852 11065 10908
rect 11001 10848 11065 10852
rect 11081 10908 11145 10912
rect 11081 10852 11085 10908
rect 11085 10852 11141 10908
rect 11141 10852 11145 10908
rect 11081 10848 11145 10852
rect 15786 10908 15850 10912
rect 15786 10852 15790 10908
rect 15790 10852 15846 10908
rect 15846 10852 15850 10908
rect 15786 10848 15850 10852
rect 15866 10908 15930 10912
rect 15866 10852 15870 10908
rect 15870 10852 15926 10908
rect 15926 10852 15930 10908
rect 15866 10848 15930 10852
rect 15946 10908 16010 10912
rect 15946 10852 15950 10908
rect 15950 10852 16006 10908
rect 16006 10852 16010 10908
rect 15946 10848 16010 10852
rect 16026 10908 16090 10912
rect 16026 10852 16030 10908
rect 16030 10852 16086 10908
rect 16086 10852 16090 10908
rect 16026 10848 16090 10852
rect 20731 10908 20795 10912
rect 20731 10852 20735 10908
rect 20735 10852 20791 10908
rect 20791 10852 20795 10908
rect 20731 10848 20795 10852
rect 20811 10908 20875 10912
rect 20811 10852 20815 10908
rect 20815 10852 20871 10908
rect 20871 10852 20875 10908
rect 20811 10848 20875 10852
rect 20891 10908 20955 10912
rect 20891 10852 20895 10908
rect 20895 10852 20951 10908
rect 20951 10852 20955 10908
rect 20891 10848 20955 10852
rect 20971 10908 21035 10912
rect 20971 10852 20975 10908
rect 20975 10852 21031 10908
rect 21031 10852 21035 10908
rect 20971 10848 21035 10852
rect 3424 10364 3488 10368
rect 3424 10308 3428 10364
rect 3428 10308 3484 10364
rect 3484 10308 3488 10364
rect 3424 10304 3488 10308
rect 3504 10364 3568 10368
rect 3504 10308 3508 10364
rect 3508 10308 3564 10364
rect 3564 10308 3568 10364
rect 3504 10304 3568 10308
rect 3584 10364 3648 10368
rect 3584 10308 3588 10364
rect 3588 10308 3644 10364
rect 3644 10308 3648 10364
rect 3584 10304 3648 10308
rect 3664 10364 3728 10368
rect 3664 10308 3668 10364
rect 3668 10308 3724 10364
rect 3724 10308 3728 10364
rect 3664 10304 3728 10308
rect 8369 10364 8433 10368
rect 8369 10308 8373 10364
rect 8373 10308 8429 10364
rect 8429 10308 8433 10364
rect 8369 10304 8433 10308
rect 8449 10364 8513 10368
rect 8449 10308 8453 10364
rect 8453 10308 8509 10364
rect 8509 10308 8513 10364
rect 8449 10304 8513 10308
rect 8529 10364 8593 10368
rect 8529 10308 8533 10364
rect 8533 10308 8589 10364
rect 8589 10308 8593 10364
rect 8529 10304 8593 10308
rect 8609 10364 8673 10368
rect 8609 10308 8613 10364
rect 8613 10308 8669 10364
rect 8669 10308 8673 10364
rect 8609 10304 8673 10308
rect 13314 10364 13378 10368
rect 13314 10308 13318 10364
rect 13318 10308 13374 10364
rect 13374 10308 13378 10364
rect 13314 10304 13378 10308
rect 13394 10364 13458 10368
rect 13394 10308 13398 10364
rect 13398 10308 13454 10364
rect 13454 10308 13458 10364
rect 13394 10304 13458 10308
rect 13474 10364 13538 10368
rect 13474 10308 13478 10364
rect 13478 10308 13534 10364
rect 13534 10308 13538 10364
rect 13474 10304 13538 10308
rect 13554 10364 13618 10368
rect 13554 10308 13558 10364
rect 13558 10308 13614 10364
rect 13614 10308 13618 10364
rect 13554 10304 13618 10308
rect 18259 10364 18323 10368
rect 18259 10308 18263 10364
rect 18263 10308 18319 10364
rect 18319 10308 18323 10364
rect 18259 10304 18323 10308
rect 18339 10364 18403 10368
rect 18339 10308 18343 10364
rect 18343 10308 18399 10364
rect 18399 10308 18403 10364
rect 18339 10304 18403 10308
rect 18419 10364 18483 10368
rect 18419 10308 18423 10364
rect 18423 10308 18479 10364
rect 18479 10308 18483 10364
rect 18419 10304 18483 10308
rect 18499 10364 18563 10368
rect 18499 10308 18503 10364
rect 18503 10308 18559 10364
rect 18559 10308 18563 10364
rect 18499 10304 18563 10308
rect 5896 9820 5960 9824
rect 5896 9764 5900 9820
rect 5900 9764 5956 9820
rect 5956 9764 5960 9820
rect 5896 9760 5960 9764
rect 5976 9820 6040 9824
rect 5976 9764 5980 9820
rect 5980 9764 6036 9820
rect 6036 9764 6040 9820
rect 5976 9760 6040 9764
rect 6056 9820 6120 9824
rect 6056 9764 6060 9820
rect 6060 9764 6116 9820
rect 6116 9764 6120 9820
rect 6056 9760 6120 9764
rect 6136 9820 6200 9824
rect 6136 9764 6140 9820
rect 6140 9764 6196 9820
rect 6196 9764 6200 9820
rect 6136 9760 6200 9764
rect 10841 9820 10905 9824
rect 10841 9764 10845 9820
rect 10845 9764 10901 9820
rect 10901 9764 10905 9820
rect 10841 9760 10905 9764
rect 10921 9820 10985 9824
rect 10921 9764 10925 9820
rect 10925 9764 10981 9820
rect 10981 9764 10985 9820
rect 10921 9760 10985 9764
rect 11001 9820 11065 9824
rect 11001 9764 11005 9820
rect 11005 9764 11061 9820
rect 11061 9764 11065 9820
rect 11001 9760 11065 9764
rect 11081 9820 11145 9824
rect 11081 9764 11085 9820
rect 11085 9764 11141 9820
rect 11141 9764 11145 9820
rect 11081 9760 11145 9764
rect 15786 9820 15850 9824
rect 15786 9764 15790 9820
rect 15790 9764 15846 9820
rect 15846 9764 15850 9820
rect 15786 9760 15850 9764
rect 15866 9820 15930 9824
rect 15866 9764 15870 9820
rect 15870 9764 15926 9820
rect 15926 9764 15930 9820
rect 15866 9760 15930 9764
rect 15946 9820 16010 9824
rect 15946 9764 15950 9820
rect 15950 9764 16006 9820
rect 16006 9764 16010 9820
rect 15946 9760 16010 9764
rect 16026 9820 16090 9824
rect 16026 9764 16030 9820
rect 16030 9764 16086 9820
rect 16086 9764 16090 9820
rect 16026 9760 16090 9764
rect 20731 9820 20795 9824
rect 20731 9764 20735 9820
rect 20735 9764 20791 9820
rect 20791 9764 20795 9820
rect 20731 9760 20795 9764
rect 20811 9820 20875 9824
rect 20811 9764 20815 9820
rect 20815 9764 20871 9820
rect 20871 9764 20875 9820
rect 20811 9760 20875 9764
rect 20891 9820 20955 9824
rect 20891 9764 20895 9820
rect 20895 9764 20951 9820
rect 20951 9764 20955 9820
rect 20891 9760 20955 9764
rect 20971 9820 21035 9824
rect 20971 9764 20975 9820
rect 20975 9764 21031 9820
rect 21031 9764 21035 9820
rect 20971 9760 21035 9764
rect 3424 9276 3488 9280
rect 3424 9220 3428 9276
rect 3428 9220 3484 9276
rect 3484 9220 3488 9276
rect 3424 9216 3488 9220
rect 3504 9276 3568 9280
rect 3504 9220 3508 9276
rect 3508 9220 3564 9276
rect 3564 9220 3568 9276
rect 3504 9216 3568 9220
rect 3584 9276 3648 9280
rect 3584 9220 3588 9276
rect 3588 9220 3644 9276
rect 3644 9220 3648 9276
rect 3584 9216 3648 9220
rect 3664 9276 3728 9280
rect 3664 9220 3668 9276
rect 3668 9220 3724 9276
rect 3724 9220 3728 9276
rect 3664 9216 3728 9220
rect 8369 9276 8433 9280
rect 8369 9220 8373 9276
rect 8373 9220 8429 9276
rect 8429 9220 8433 9276
rect 8369 9216 8433 9220
rect 8449 9276 8513 9280
rect 8449 9220 8453 9276
rect 8453 9220 8509 9276
rect 8509 9220 8513 9276
rect 8449 9216 8513 9220
rect 8529 9276 8593 9280
rect 8529 9220 8533 9276
rect 8533 9220 8589 9276
rect 8589 9220 8593 9276
rect 8529 9216 8593 9220
rect 8609 9276 8673 9280
rect 8609 9220 8613 9276
rect 8613 9220 8669 9276
rect 8669 9220 8673 9276
rect 8609 9216 8673 9220
rect 13314 9276 13378 9280
rect 13314 9220 13318 9276
rect 13318 9220 13374 9276
rect 13374 9220 13378 9276
rect 13314 9216 13378 9220
rect 13394 9276 13458 9280
rect 13394 9220 13398 9276
rect 13398 9220 13454 9276
rect 13454 9220 13458 9276
rect 13394 9216 13458 9220
rect 13474 9276 13538 9280
rect 13474 9220 13478 9276
rect 13478 9220 13534 9276
rect 13534 9220 13538 9276
rect 13474 9216 13538 9220
rect 13554 9276 13618 9280
rect 13554 9220 13558 9276
rect 13558 9220 13614 9276
rect 13614 9220 13618 9276
rect 13554 9216 13618 9220
rect 18259 9276 18323 9280
rect 18259 9220 18263 9276
rect 18263 9220 18319 9276
rect 18319 9220 18323 9276
rect 18259 9216 18323 9220
rect 18339 9276 18403 9280
rect 18339 9220 18343 9276
rect 18343 9220 18399 9276
rect 18399 9220 18403 9276
rect 18339 9216 18403 9220
rect 18419 9276 18483 9280
rect 18419 9220 18423 9276
rect 18423 9220 18479 9276
rect 18479 9220 18483 9276
rect 18419 9216 18483 9220
rect 18499 9276 18563 9280
rect 18499 9220 18503 9276
rect 18503 9220 18559 9276
rect 18559 9220 18563 9276
rect 18499 9216 18563 9220
rect 5896 8732 5960 8736
rect 5896 8676 5900 8732
rect 5900 8676 5956 8732
rect 5956 8676 5960 8732
rect 5896 8672 5960 8676
rect 5976 8732 6040 8736
rect 5976 8676 5980 8732
rect 5980 8676 6036 8732
rect 6036 8676 6040 8732
rect 5976 8672 6040 8676
rect 6056 8732 6120 8736
rect 6056 8676 6060 8732
rect 6060 8676 6116 8732
rect 6116 8676 6120 8732
rect 6056 8672 6120 8676
rect 6136 8732 6200 8736
rect 6136 8676 6140 8732
rect 6140 8676 6196 8732
rect 6196 8676 6200 8732
rect 6136 8672 6200 8676
rect 10841 8732 10905 8736
rect 10841 8676 10845 8732
rect 10845 8676 10901 8732
rect 10901 8676 10905 8732
rect 10841 8672 10905 8676
rect 10921 8732 10985 8736
rect 10921 8676 10925 8732
rect 10925 8676 10981 8732
rect 10981 8676 10985 8732
rect 10921 8672 10985 8676
rect 11001 8732 11065 8736
rect 11001 8676 11005 8732
rect 11005 8676 11061 8732
rect 11061 8676 11065 8732
rect 11001 8672 11065 8676
rect 11081 8732 11145 8736
rect 11081 8676 11085 8732
rect 11085 8676 11141 8732
rect 11141 8676 11145 8732
rect 11081 8672 11145 8676
rect 15786 8732 15850 8736
rect 15786 8676 15790 8732
rect 15790 8676 15846 8732
rect 15846 8676 15850 8732
rect 15786 8672 15850 8676
rect 15866 8732 15930 8736
rect 15866 8676 15870 8732
rect 15870 8676 15926 8732
rect 15926 8676 15930 8732
rect 15866 8672 15930 8676
rect 15946 8732 16010 8736
rect 15946 8676 15950 8732
rect 15950 8676 16006 8732
rect 16006 8676 16010 8732
rect 15946 8672 16010 8676
rect 16026 8732 16090 8736
rect 16026 8676 16030 8732
rect 16030 8676 16086 8732
rect 16086 8676 16090 8732
rect 16026 8672 16090 8676
rect 20731 8732 20795 8736
rect 20731 8676 20735 8732
rect 20735 8676 20791 8732
rect 20791 8676 20795 8732
rect 20731 8672 20795 8676
rect 20811 8732 20875 8736
rect 20811 8676 20815 8732
rect 20815 8676 20871 8732
rect 20871 8676 20875 8732
rect 20811 8672 20875 8676
rect 20891 8732 20955 8736
rect 20891 8676 20895 8732
rect 20895 8676 20951 8732
rect 20951 8676 20955 8732
rect 20891 8672 20955 8676
rect 20971 8732 21035 8736
rect 20971 8676 20975 8732
rect 20975 8676 21031 8732
rect 21031 8676 21035 8732
rect 20971 8672 21035 8676
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 3584 8188 3648 8192
rect 3584 8132 3588 8188
rect 3588 8132 3644 8188
rect 3644 8132 3648 8188
rect 3584 8128 3648 8132
rect 3664 8188 3728 8192
rect 3664 8132 3668 8188
rect 3668 8132 3724 8188
rect 3724 8132 3728 8188
rect 3664 8128 3728 8132
rect 8369 8188 8433 8192
rect 8369 8132 8373 8188
rect 8373 8132 8429 8188
rect 8429 8132 8433 8188
rect 8369 8128 8433 8132
rect 8449 8188 8513 8192
rect 8449 8132 8453 8188
rect 8453 8132 8509 8188
rect 8509 8132 8513 8188
rect 8449 8128 8513 8132
rect 8529 8188 8593 8192
rect 8529 8132 8533 8188
rect 8533 8132 8589 8188
rect 8589 8132 8593 8188
rect 8529 8128 8593 8132
rect 8609 8188 8673 8192
rect 8609 8132 8613 8188
rect 8613 8132 8669 8188
rect 8669 8132 8673 8188
rect 8609 8128 8673 8132
rect 13314 8188 13378 8192
rect 13314 8132 13318 8188
rect 13318 8132 13374 8188
rect 13374 8132 13378 8188
rect 13314 8128 13378 8132
rect 13394 8188 13458 8192
rect 13394 8132 13398 8188
rect 13398 8132 13454 8188
rect 13454 8132 13458 8188
rect 13394 8128 13458 8132
rect 13474 8188 13538 8192
rect 13474 8132 13478 8188
rect 13478 8132 13534 8188
rect 13534 8132 13538 8188
rect 13474 8128 13538 8132
rect 13554 8188 13618 8192
rect 13554 8132 13558 8188
rect 13558 8132 13614 8188
rect 13614 8132 13618 8188
rect 13554 8128 13618 8132
rect 18259 8188 18323 8192
rect 18259 8132 18263 8188
rect 18263 8132 18319 8188
rect 18319 8132 18323 8188
rect 18259 8128 18323 8132
rect 18339 8188 18403 8192
rect 18339 8132 18343 8188
rect 18343 8132 18399 8188
rect 18399 8132 18403 8188
rect 18339 8128 18403 8132
rect 18419 8188 18483 8192
rect 18419 8132 18423 8188
rect 18423 8132 18479 8188
rect 18479 8132 18483 8188
rect 18419 8128 18483 8132
rect 18499 8188 18563 8192
rect 18499 8132 18503 8188
rect 18503 8132 18559 8188
rect 18559 8132 18563 8188
rect 18499 8128 18563 8132
rect 5896 7644 5960 7648
rect 5896 7588 5900 7644
rect 5900 7588 5956 7644
rect 5956 7588 5960 7644
rect 5896 7584 5960 7588
rect 5976 7644 6040 7648
rect 5976 7588 5980 7644
rect 5980 7588 6036 7644
rect 6036 7588 6040 7644
rect 5976 7584 6040 7588
rect 6056 7644 6120 7648
rect 6056 7588 6060 7644
rect 6060 7588 6116 7644
rect 6116 7588 6120 7644
rect 6056 7584 6120 7588
rect 6136 7644 6200 7648
rect 6136 7588 6140 7644
rect 6140 7588 6196 7644
rect 6196 7588 6200 7644
rect 6136 7584 6200 7588
rect 10841 7644 10905 7648
rect 10841 7588 10845 7644
rect 10845 7588 10901 7644
rect 10901 7588 10905 7644
rect 10841 7584 10905 7588
rect 10921 7644 10985 7648
rect 10921 7588 10925 7644
rect 10925 7588 10981 7644
rect 10981 7588 10985 7644
rect 10921 7584 10985 7588
rect 11001 7644 11065 7648
rect 11001 7588 11005 7644
rect 11005 7588 11061 7644
rect 11061 7588 11065 7644
rect 11001 7584 11065 7588
rect 11081 7644 11145 7648
rect 11081 7588 11085 7644
rect 11085 7588 11141 7644
rect 11141 7588 11145 7644
rect 11081 7584 11145 7588
rect 15786 7644 15850 7648
rect 15786 7588 15790 7644
rect 15790 7588 15846 7644
rect 15846 7588 15850 7644
rect 15786 7584 15850 7588
rect 15866 7644 15930 7648
rect 15866 7588 15870 7644
rect 15870 7588 15926 7644
rect 15926 7588 15930 7644
rect 15866 7584 15930 7588
rect 15946 7644 16010 7648
rect 15946 7588 15950 7644
rect 15950 7588 16006 7644
rect 16006 7588 16010 7644
rect 15946 7584 16010 7588
rect 16026 7644 16090 7648
rect 16026 7588 16030 7644
rect 16030 7588 16086 7644
rect 16086 7588 16090 7644
rect 16026 7584 16090 7588
rect 20731 7644 20795 7648
rect 20731 7588 20735 7644
rect 20735 7588 20791 7644
rect 20791 7588 20795 7644
rect 20731 7584 20795 7588
rect 20811 7644 20875 7648
rect 20811 7588 20815 7644
rect 20815 7588 20871 7644
rect 20871 7588 20875 7644
rect 20811 7584 20875 7588
rect 20891 7644 20955 7648
rect 20891 7588 20895 7644
rect 20895 7588 20951 7644
rect 20951 7588 20955 7644
rect 20891 7584 20955 7588
rect 20971 7644 21035 7648
rect 20971 7588 20975 7644
rect 20975 7588 21031 7644
rect 21031 7588 21035 7644
rect 20971 7584 21035 7588
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 3584 7100 3648 7104
rect 3584 7044 3588 7100
rect 3588 7044 3644 7100
rect 3644 7044 3648 7100
rect 3584 7040 3648 7044
rect 3664 7100 3728 7104
rect 3664 7044 3668 7100
rect 3668 7044 3724 7100
rect 3724 7044 3728 7100
rect 3664 7040 3728 7044
rect 8369 7100 8433 7104
rect 8369 7044 8373 7100
rect 8373 7044 8429 7100
rect 8429 7044 8433 7100
rect 8369 7040 8433 7044
rect 8449 7100 8513 7104
rect 8449 7044 8453 7100
rect 8453 7044 8509 7100
rect 8509 7044 8513 7100
rect 8449 7040 8513 7044
rect 8529 7100 8593 7104
rect 8529 7044 8533 7100
rect 8533 7044 8589 7100
rect 8589 7044 8593 7100
rect 8529 7040 8593 7044
rect 8609 7100 8673 7104
rect 8609 7044 8613 7100
rect 8613 7044 8669 7100
rect 8669 7044 8673 7100
rect 8609 7040 8673 7044
rect 13314 7100 13378 7104
rect 13314 7044 13318 7100
rect 13318 7044 13374 7100
rect 13374 7044 13378 7100
rect 13314 7040 13378 7044
rect 13394 7100 13458 7104
rect 13394 7044 13398 7100
rect 13398 7044 13454 7100
rect 13454 7044 13458 7100
rect 13394 7040 13458 7044
rect 13474 7100 13538 7104
rect 13474 7044 13478 7100
rect 13478 7044 13534 7100
rect 13534 7044 13538 7100
rect 13474 7040 13538 7044
rect 13554 7100 13618 7104
rect 13554 7044 13558 7100
rect 13558 7044 13614 7100
rect 13614 7044 13618 7100
rect 13554 7040 13618 7044
rect 18259 7100 18323 7104
rect 18259 7044 18263 7100
rect 18263 7044 18319 7100
rect 18319 7044 18323 7100
rect 18259 7040 18323 7044
rect 18339 7100 18403 7104
rect 18339 7044 18343 7100
rect 18343 7044 18399 7100
rect 18399 7044 18403 7100
rect 18339 7040 18403 7044
rect 18419 7100 18483 7104
rect 18419 7044 18423 7100
rect 18423 7044 18479 7100
rect 18479 7044 18483 7100
rect 18419 7040 18483 7044
rect 18499 7100 18563 7104
rect 18499 7044 18503 7100
rect 18503 7044 18559 7100
rect 18559 7044 18563 7100
rect 18499 7040 18563 7044
rect 5896 6556 5960 6560
rect 5896 6500 5900 6556
rect 5900 6500 5956 6556
rect 5956 6500 5960 6556
rect 5896 6496 5960 6500
rect 5976 6556 6040 6560
rect 5976 6500 5980 6556
rect 5980 6500 6036 6556
rect 6036 6500 6040 6556
rect 5976 6496 6040 6500
rect 6056 6556 6120 6560
rect 6056 6500 6060 6556
rect 6060 6500 6116 6556
rect 6116 6500 6120 6556
rect 6056 6496 6120 6500
rect 6136 6556 6200 6560
rect 6136 6500 6140 6556
rect 6140 6500 6196 6556
rect 6196 6500 6200 6556
rect 6136 6496 6200 6500
rect 10841 6556 10905 6560
rect 10841 6500 10845 6556
rect 10845 6500 10901 6556
rect 10901 6500 10905 6556
rect 10841 6496 10905 6500
rect 10921 6556 10985 6560
rect 10921 6500 10925 6556
rect 10925 6500 10981 6556
rect 10981 6500 10985 6556
rect 10921 6496 10985 6500
rect 11001 6556 11065 6560
rect 11001 6500 11005 6556
rect 11005 6500 11061 6556
rect 11061 6500 11065 6556
rect 11001 6496 11065 6500
rect 11081 6556 11145 6560
rect 11081 6500 11085 6556
rect 11085 6500 11141 6556
rect 11141 6500 11145 6556
rect 11081 6496 11145 6500
rect 15786 6556 15850 6560
rect 15786 6500 15790 6556
rect 15790 6500 15846 6556
rect 15846 6500 15850 6556
rect 15786 6496 15850 6500
rect 15866 6556 15930 6560
rect 15866 6500 15870 6556
rect 15870 6500 15926 6556
rect 15926 6500 15930 6556
rect 15866 6496 15930 6500
rect 15946 6556 16010 6560
rect 15946 6500 15950 6556
rect 15950 6500 16006 6556
rect 16006 6500 16010 6556
rect 15946 6496 16010 6500
rect 16026 6556 16090 6560
rect 16026 6500 16030 6556
rect 16030 6500 16086 6556
rect 16086 6500 16090 6556
rect 16026 6496 16090 6500
rect 20731 6556 20795 6560
rect 20731 6500 20735 6556
rect 20735 6500 20791 6556
rect 20791 6500 20795 6556
rect 20731 6496 20795 6500
rect 20811 6556 20875 6560
rect 20811 6500 20815 6556
rect 20815 6500 20871 6556
rect 20871 6500 20875 6556
rect 20811 6496 20875 6500
rect 20891 6556 20955 6560
rect 20891 6500 20895 6556
rect 20895 6500 20951 6556
rect 20951 6500 20955 6556
rect 20891 6496 20955 6500
rect 20971 6556 21035 6560
rect 20971 6500 20975 6556
rect 20975 6500 21031 6556
rect 21031 6500 21035 6556
rect 20971 6496 21035 6500
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 3584 6012 3648 6016
rect 3584 5956 3588 6012
rect 3588 5956 3644 6012
rect 3644 5956 3648 6012
rect 3584 5952 3648 5956
rect 3664 6012 3728 6016
rect 3664 5956 3668 6012
rect 3668 5956 3724 6012
rect 3724 5956 3728 6012
rect 3664 5952 3728 5956
rect 8369 6012 8433 6016
rect 8369 5956 8373 6012
rect 8373 5956 8429 6012
rect 8429 5956 8433 6012
rect 8369 5952 8433 5956
rect 8449 6012 8513 6016
rect 8449 5956 8453 6012
rect 8453 5956 8509 6012
rect 8509 5956 8513 6012
rect 8449 5952 8513 5956
rect 8529 6012 8593 6016
rect 8529 5956 8533 6012
rect 8533 5956 8589 6012
rect 8589 5956 8593 6012
rect 8529 5952 8593 5956
rect 8609 6012 8673 6016
rect 8609 5956 8613 6012
rect 8613 5956 8669 6012
rect 8669 5956 8673 6012
rect 8609 5952 8673 5956
rect 13314 6012 13378 6016
rect 13314 5956 13318 6012
rect 13318 5956 13374 6012
rect 13374 5956 13378 6012
rect 13314 5952 13378 5956
rect 13394 6012 13458 6016
rect 13394 5956 13398 6012
rect 13398 5956 13454 6012
rect 13454 5956 13458 6012
rect 13394 5952 13458 5956
rect 13474 6012 13538 6016
rect 13474 5956 13478 6012
rect 13478 5956 13534 6012
rect 13534 5956 13538 6012
rect 13474 5952 13538 5956
rect 13554 6012 13618 6016
rect 13554 5956 13558 6012
rect 13558 5956 13614 6012
rect 13614 5956 13618 6012
rect 13554 5952 13618 5956
rect 18259 6012 18323 6016
rect 18259 5956 18263 6012
rect 18263 5956 18319 6012
rect 18319 5956 18323 6012
rect 18259 5952 18323 5956
rect 18339 6012 18403 6016
rect 18339 5956 18343 6012
rect 18343 5956 18399 6012
rect 18399 5956 18403 6012
rect 18339 5952 18403 5956
rect 18419 6012 18483 6016
rect 18419 5956 18423 6012
rect 18423 5956 18479 6012
rect 18479 5956 18483 6012
rect 18419 5952 18483 5956
rect 18499 6012 18563 6016
rect 18499 5956 18503 6012
rect 18503 5956 18559 6012
rect 18559 5956 18563 6012
rect 18499 5952 18563 5956
rect 5896 5468 5960 5472
rect 5896 5412 5900 5468
rect 5900 5412 5956 5468
rect 5956 5412 5960 5468
rect 5896 5408 5960 5412
rect 5976 5468 6040 5472
rect 5976 5412 5980 5468
rect 5980 5412 6036 5468
rect 6036 5412 6040 5468
rect 5976 5408 6040 5412
rect 6056 5468 6120 5472
rect 6056 5412 6060 5468
rect 6060 5412 6116 5468
rect 6116 5412 6120 5468
rect 6056 5408 6120 5412
rect 6136 5468 6200 5472
rect 6136 5412 6140 5468
rect 6140 5412 6196 5468
rect 6196 5412 6200 5468
rect 6136 5408 6200 5412
rect 10841 5468 10905 5472
rect 10841 5412 10845 5468
rect 10845 5412 10901 5468
rect 10901 5412 10905 5468
rect 10841 5408 10905 5412
rect 10921 5468 10985 5472
rect 10921 5412 10925 5468
rect 10925 5412 10981 5468
rect 10981 5412 10985 5468
rect 10921 5408 10985 5412
rect 11001 5468 11065 5472
rect 11001 5412 11005 5468
rect 11005 5412 11061 5468
rect 11061 5412 11065 5468
rect 11001 5408 11065 5412
rect 11081 5468 11145 5472
rect 11081 5412 11085 5468
rect 11085 5412 11141 5468
rect 11141 5412 11145 5468
rect 11081 5408 11145 5412
rect 15786 5468 15850 5472
rect 15786 5412 15790 5468
rect 15790 5412 15846 5468
rect 15846 5412 15850 5468
rect 15786 5408 15850 5412
rect 15866 5468 15930 5472
rect 15866 5412 15870 5468
rect 15870 5412 15926 5468
rect 15926 5412 15930 5468
rect 15866 5408 15930 5412
rect 15946 5468 16010 5472
rect 15946 5412 15950 5468
rect 15950 5412 16006 5468
rect 16006 5412 16010 5468
rect 15946 5408 16010 5412
rect 16026 5468 16090 5472
rect 16026 5412 16030 5468
rect 16030 5412 16086 5468
rect 16086 5412 16090 5468
rect 16026 5408 16090 5412
rect 20731 5468 20795 5472
rect 20731 5412 20735 5468
rect 20735 5412 20791 5468
rect 20791 5412 20795 5468
rect 20731 5408 20795 5412
rect 20811 5468 20875 5472
rect 20811 5412 20815 5468
rect 20815 5412 20871 5468
rect 20871 5412 20875 5468
rect 20811 5408 20875 5412
rect 20891 5468 20955 5472
rect 20891 5412 20895 5468
rect 20895 5412 20951 5468
rect 20951 5412 20955 5468
rect 20891 5408 20955 5412
rect 20971 5468 21035 5472
rect 20971 5412 20975 5468
rect 20975 5412 21031 5468
rect 21031 5412 21035 5468
rect 20971 5408 21035 5412
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 3584 4924 3648 4928
rect 3584 4868 3588 4924
rect 3588 4868 3644 4924
rect 3644 4868 3648 4924
rect 3584 4864 3648 4868
rect 3664 4924 3728 4928
rect 3664 4868 3668 4924
rect 3668 4868 3724 4924
rect 3724 4868 3728 4924
rect 3664 4864 3728 4868
rect 8369 4924 8433 4928
rect 8369 4868 8373 4924
rect 8373 4868 8429 4924
rect 8429 4868 8433 4924
rect 8369 4864 8433 4868
rect 8449 4924 8513 4928
rect 8449 4868 8453 4924
rect 8453 4868 8509 4924
rect 8509 4868 8513 4924
rect 8449 4864 8513 4868
rect 8529 4924 8593 4928
rect 8529 4868 8533 4924
rect 8533 4868 8589 4924
rect 8589 4868 8593 4924
rect 8529 4864 8593 4868
rect 8609 4924 8673 4928
rect 8609 4868 8613 4924
rect 8613 4868 8669 4924
rect 8669 4868 8673 4924
rect 8609 4864 8673 4868
rect 13314 4924 13378 4928
rect 13314 4868 13318 4924
rect 13318 4868 13374 4924
rect 13374 4868 13378 4924
rect 13314 4864 13378 4868
rect 13394 4924 13458 4928
rect 13394 4868 13398 4924
rect 13398 4868 13454 4924
rect 13454 4868 13458 4924
rect 13394 4864 13458 4868
rect 13474 4924 13538 4928
rect 13474 4868 13478 4924
rect 13478 4868 13534 4924
rect 13534 4868 13538 4924
rect 13474 4864 13538 4868
rect 13554 4924 13618 4928
rect 13554 4868 13558 4924
rect 13558 4868 13614 4924
rect 13614 4868 13618 4924
rect 13554 4864 13618 4868
rect 18259 4924 18323 4928
rect 18259 4868 18263 4924
rect 18263 4868 18319 4924
rect 18319 4868 18323 4924
rect 18259 4864 18323 4868
rect 18339 4924 18403 4928
rect 18339 4868 18343 4924
rect 18343 4868 18399 4924
rect 18399 4868 18403 4924
rect 18339 4864 18403 4868
rect 18419 4924 18483 4928
rect 18419 4868 18423 4924
rect 18423 4868 18479 4924
rect 18479 4868 18483 4924
rect 18419 4864 18483 4868
rect 18499 4924 18563 4928
rect 18499 4868 18503 4924
rect 18503 4868 18559 4924
rect 18559 4868 18563 4924
rect 18499 4864 18563 4868
rect 5896 4380 5960 4384
rect 5896 4324 5900 4380
rect 5900 4324 5956 4380
rect 5956 4324 5960 4380
rect 5896 4320 5960 4324
rect 5976 4380 6040 4384
rect 5976 4324 5980 4380
rect 5980 4324 6036 4380
rect 6036 4324 6040 4380
rect 5976 4320 6040 4324
rect 6056 4380 6120 4384
rect 6056 4324 6060 4380
rect 6060 4324 6116 4380
rect 6116 4324 6120 4380
rect 6056 4320 6120 4324
rect 6136 4380 6200 4384
rect 6136 4324 6140 4380
rect 6140 4324 6196 4380
rect 6196 4324 6200 4380
rect 6136 4320 6200 4324
rect 10841 4380 10905 4384
rect 10841 4324 10845 4380
rect 10845 4324 10901 4380
rect 10901 4324 10905 4380
rect 10841 4320 10905 4324
rect 10921 4380 10985 4384
rect 10921 4324 10925 4380
rect 10925 4324 10981 4380
rect 10981 4324 10985 4380
rect 10921 4320 10985 4324
rect 11001 4380 11065 4384
rect 11001 4324 11005 4380
rect 11005 4324 11061 4380
rect 11061 4324 11065 4380
rect 11001 4320 11065 4324
rect 11081 4380 11145 4384
rect 11081 4324 11085 4380
rect 11085 4324 11141 4380
rect 11141 4324 11145 4380
rect 11081 4320 11145 4324
rect 15786 4380 15850 4384
rect 15786 4324 15790 4380
rect 15790 4324 15846 4380
rect 15846 4324 15850 4380
rect 15786 4320 15850 4324
rect 15866 4380 15930 4384
rect 15866 4324 15870 4380
rect 15870 4324 15926 4380
rect 15926 4324 15930 4380
rect 15866 4320 15930 4324
rect 15946 4380 16010 4384
rect 15946 4324 15950 4380
rect 15950 4324 16006 4380
rect 16006 4324 16010 4380
rect 15946 4320 16010 4324
rect 16026 4380 16090 4384
rect 16026 4324 16030 4380
rect 16030 4324 16086 4380
rect 16086 4324 16090 4380
rect 16026 4320 16090 4324
rect 20731 4380 20795 4384
rect 20731 4324 20735 4380
rect 20735 4324 20791 4380
rect 20791 4324 20795 4380
rect 20731 4320 20795 4324
rect 20811 4380 20875 4384
rect 20811 4324 20815 4380
rect 20815 4324 20871 4380
rect 20871 4324 20875 4380
rect 20811 4320 20875 4324
rect 20891 4380 20955 4384
rect 20891 4324 20895 4380
rect 20895 4324 20951 4380
rect 20951 4324 20955 4380
rect 20891 4320 20955 4324
rect 20971 4380 21035 4384
rect 20971 4324 20975 4380
rect 20975 4324 21031 4380
rect 21031 4324 21035 4380
rect 20971 4320 21035 4324
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 3584 3836 3648 3840
rect 3584 3780 3588 3836
rect 3588 3780 3644 3836
rect 3644 3780 3648 3836
rect 3584 3776 3648 3780
rect 3664 3836 3728 3840
rect 3664 3780 3668 3836
rect 3668 3780 3724 3836
rect 3724 3780 3728 3836
rect 3664 3776 3728 3780
rect 8369 3836 8433 3840
rect 8369 3780 8373 3836
rect 8373 3780 8429 3836
rect 8429 3780 8433 3836
rect 8369 3776 8433 3780
rect 8449 3836 8513 3840
rect 8449 3780 8453 3836
rect 8453 3780 8509 3836
rect 8509 3780 8513 3836
rect 8449 3776 8513 3780
rect 8529 3836 8593 3840
rect 8529 3780 8533 3836
rect 8533 3780 8589 3836
rect 8589 3780 8593 3836
rect 8529 3776 8593 3780
rect 8609 3836 8673 3840
rect 8609 3780 8613 3836
rect 8613 3780 8669 3836
rect 8669 3780 8673 3836
rect 8609 3776 8673 3780
rect 13314 3836 13378 3840
rect 13314 3780 13318 3836
rect 13318 3780 13374 3836
rect 13374 3780 13378 3836
rect 13314 3776 13378 3780
rect 13394 3836 13458 3840
rect 13394 3780 13398 3836
rect 13398 3780 13454 3836
rect 13454 3780 13458 3836
rect 13394 3776 13458 3780
rect 13474 3836 13538 3840
rect 13474 3780 13478 3836
rect 13478 3780 13534 3836
rect 13534 3780 13538 3836
rect 13474 3776 13538 3780
rect 13554 3836 13618 3840
rect 13554 3780 13558 3836
rect 13558 3780 13614 3836
rect 13614 3780 13618 3836
rect 13554 3776 13618 3780
rect 18259 3836 18323 3840
rect 18259 3780 18263 3836
rect 18263 3780 18319 3836
rect 18319 3780 18323 3836
rect 18259 3776 18323 3780
rect 18339 3836 18403 3840
rect 18339 3780 18343 3836
rect 18343 3780 18399 3836
rect 18399 3780 18403 3836
rect 18339 3776 18403 3780
rect 18419 3836 18483 3840
rect 18419 3780 18423 3836
rect 18423 3780 18479 3836
rect 18479 3780 18483 3836
rect 18419 3776 18483 3780
rect 18499 3836 18563 3840
rect 18499 3780 18503 3836
rect 18503 3780 18559 3836
rect 18559 3780 18563 3836
rect 18499 3776 18563 3780
rect 5896 3292 5960 3296
rect 5896 3236 5900 3292
rect 5900 3236 5956 3292
rect 5956 3236 5960 3292
rect 5896 3232 5960 3236
rect 5976 3292 6040 3296
rect 5976 3236 5980 3292
rect 5980 3236 6036 3292
rect 6036 3236 6040 3292
rect 5976 3232 6040 3236
rect 6056 3292 6120 3296
rect 6056 3236 6060 3292
rect 6060 3236 6116 3292
rect 6116 3236 6120 3292
rect 6056 3232 6120 3236
rect 6136 3292 6200 3296
rect 6136 3236 6140 3292
rect 6140 3236 6196 3292
rect 6196 3236 6200 3292
rect 6136 3232 6200 3236
rect 10841 3292 10905 3296
rect 10841 3236 10845 3292
rect 10845 3236 10901 3292
rect 10901 3236 10905 3292
rect 10841 3232 10905 3236
rect 10921 3292 10985 3296
rect 10921 3236 10925 3292
rect 10925 3236 10981 3292
rect 10981 3236 10985 3292
rect 10921 3232 10985 3236
rect 11001 3292 11065 3296
rect 11001 3236 11005 3292
rect 11005 3236 11061 3292
rect 11061 3236 11065 3292
rect 11001 3232 11065 3236
rect 11081 3292 11145 3296
rect 11081 3236 11085 3292
rect 11085 3236 11141 3292
rect 11141 3236 11145 3292
rect 11081 3232 11145 3236
rect 15786 3292 15850 3296
rect 15786 3236 15790 3292
rect 15790 3236 15846 3292
rect 15846 3236 15850 3292
rect 15786 3232 15850 3236
rect 15866 3292 15930 3296
rect 15866 3236 15870 3292
rect 15870 3236 15926 3292
rect 15926 3236 15930 3292
rect 15866 3232 15930 3236
rect 15946 3292 16010 3296
rect 15946 3236 15950 3292
rect 15950 3236 16006 3292
rect 16006 3236 16010 3292
rect 15946 3232 16010 3236
rect 16026 3292 16090 3296
rect 16026 3236 16030 3292
rect 16030 3236 16086 3292
rect 16086 3236 16090 3292
rect 16026 3232 16090 3236
rect 20731 3292 20795 3296
rect 20731 3236 20735 3292
rect 20735 3236 20791 3292
rect 20791 3236 20795 3292
rect 20731 3232 20795 3236
rect 20811 3292 20875 3296
rect 20811 3236 20815 3292
rect 20815 3236 20871 3292
rect 20871 3236 20875 3292
rect 20811 3232 20875 3236
rect 20891 3292 20955 3296
rect 20891 3236 20895 3292
rect 20895 3236 20951 3292
rect 20951 3236 20955 3292
rect 20891 3232 20955 3236
rect 20971 3292 21035 3296
rect 20971 3236 20975 3292
rect 20975 3236 21031 3292
rect 21031 3236 21035 3292
rect 20971 3232 21035 3236
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 3584 2748 3648 2752
rect 3584 2692 3588 2748
rect 3588 2692 3644 2748
rect 3644 2692 3648 2748
rect 3584 2688 3648 2692
rect 3664 2748 3728 2752
rect 3664 2692 3668 2748
rect 3668 2692 3724 2748
rect 3724 2692 3728 2748
rect 3664 2688 3728 2692
rect 8369 2748 8433 2752
rect 8369 2692 8373 2748
rect 8373 2692 8429 2748
rect 8429 2692 8433 2748
rect 8369 2688 8433 2692
rect 8449 2748 8513 2752
rect 8449 2692 8453 2748
rect 8453 2692 8509 2748
rect 8509 2692 8513 2748
rect 8449 2688 8513 2692
rect 8529 2748 8593 2752
rect 8529 2692 8533 2748
rect 8533 2692 8589 2748
rect 8589 2692 8593 2748
rect 8529 2688 8593 2692
rect 8609 2748 8673 2752
rect 8609 2692 8613 2748
rect 8613 2692 8669 2748
rect 8669 2692 8673 2748
rect 8609 2688 8673 2692
rect 13314 2748 13378 2752
rect 13314 2692 13318 2748
rect 13318 2692 13374 2748
rect 13374 2692 13378 2748
rect 13314 2688 13378 2692
rect 13394 2748 13458 2752
rect 13394 2692 13398 2748
rect 13398 2692 13454 2748
rect 13454 2692 13458 2748
rect 13394 2688 13458 2692
rect 13474 2748 13538 2752
rect 13474 2692 13478 2748
rect 13478 2692 13534 2748
rect 13534 2692 13538 2748
rect 13474 2688 13538 2692
rect 13554 2748 13618 2752
rect 13554 2692 13558 2748
rect 13558 2692 13614 2748
rect 13614 2692 13618 2748
rect 13554 2688 13618 2692
rect 18259 2748 18323 2752
rect 18259 2692 18263 2748
rect 18263 2692 18319 2748
rect 18319 2692 18323 2748
rect 18259 2688 18323 2692
rect 18339 2748 18403 2752
rect 18339 2692 18343 2748
rect 18343 2692 18399 2748
rect 18399 2692 18403 2748
rect 18339 2688 18403 2692
rect 18419 2748 18483 2752
rect 18419 2692 18423 2748
rect 18423 2692 18479 2748
rect 18479 2692 18483 2748
rect 18419 2688 18483 2692
rect 18499 2748 18563 2752
rect 18499 2692 18503 2748
rect 18503 2692 18559 2748
rect 18559 2692 18563 2748
rect 18499 2688 18563 2692
rect 5896 2204 5960 2208
rect 5896 2148 5900 2204
rect 5900 2148 5956 2204
rect 5956 2148 5960 2204
rect 5896 2144 5960 2148
rect 5976 2204 6040 2208
rect 5976 2148 5980 2204
rect 5980 2148 6036 2204
rect 6036 2148 6040 2204
rect 5976 2144 6040 2148
rect 6056 2204 6120 2208
rect 6056 2148 6060 2204
rect 6060 2148 6116 2204
rect 6116 2148 6120 2204
rect 6056 2144 6120 2148
rect 6136 2204 6200 2208
rect 6136 2148 6140 2204
rect 6140 2148 6196 2204
rect 6196 2148 6200 2204
rect 6136 2144 6200 2148
rect 10841 2204 10905 2208
rect 10841 2148 10845 2204
rect 10845 2148 10901 2204
rect 10901 2148 10905 2204
rect 10841 2144 10905 2148
rect 10921 2204 10985 2208
rect 10921 2148 10925 2204
rect 10925 2148 10981 2204
rect 10981 2148 10985 2204
rect 10921 2144 10985 2148
rect 11001 2204 11065 2208
rect 11001 2148 11005 2204
rect 11005 2148 11061 2204
rect 11061 2148 11065 2204
rect 11001 2144 11065 2148
rect 11081 2204 11145 2208
rect 11081 2148 11085 2204
rect 11085 2148 11141 2204
rect 11141 2148 11145 2204
rect 11081 2144 11145 2148
rect 15786 2204 15850 2208
rect 15786 2148 15790 2204
rect 15790 2148 15846 2204
rect 15846 2148 15850 2204
rect 15786 2144 15850 2148
rect 15866 2204 15930 2208
rect 15866 2148 15870 2204
rect 15870 2148 15926 2204
rect 15926 2148 15930 2204
rect 15866 2144 15930 2148
rect 15946 2204 16010 2208
rect 15946 2148 15950 2204
rect 15950 2148 16006 2204
rect 16006 2148 16010 2204
rect 15946 2144 16010 2148
rect 16026 2204 16090 2208
rect 16026 2148 16030 2204
rect 16030 2148 16086 2204
rect 16086 2148 16090 2204
rect 16026 2144 16090 2148
rect 20731 2204 20795 2208
rect 20731 2148 20735 2204
rect 20735 2148 20791 2204
rect 20791 2148 20795 2204
rect 20731 2144 20795 2148
rect 20811 2204 20875 2208
rect 20811 2148 20815 2204
rect 20815 2148 20871 2204
rect 20871 2148 20875 2204
rect 20811 2144 20875 2148
rect 20891 2204 20955 2208
rect 20891 2148 20895 2204
rect 20895 2148 20951 2204
rect 20951 2148 20955 2204
rect 20891 2144 20955 2148
rect 20971 2204 21035 2208
rect 20971 2148 20975 2204
rect 20975 2148 21031 2204
rect 21031 2148 21035 2204
rect 20971 2144 21035 2148
<< metal4 >>
rect 3416 19072 3736 19632
rect 3416 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3736 19072
rect 3416 17984 3736 19008
rect 3416 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3736 17984
rect 3416 16896 3736 17920
rect 3416 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3736 16896
rect 3416 15808 3736 16832
rect 3416 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3736 15808
rect 3416 14720 3736 15744
rect 3416 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3736 14720
rect 3416 13632 3736 14656
rect 3416 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3736 13632
rect 3416 12544 3736 13568
rect 3416 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3736 12544
rect 3416 11456 3736 12480
rect 3416 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3736 11456
rect 3416 10368 3736 11392
rect 3416 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3736 10368
rect 3416 9280 3736 10304
rect 3416 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3736 9280
rect 3416 8192 3736 9216
rect 3416 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3736 8192
rect 3416 7104 3736 8128
rect 3416 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3736 7104
rect 3416 6016 3736 7040
rect 3416 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3736 6016
rect 3416 4928 3736 5952
rect 3416 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3736 4928
rect 3416 3840 3736 4864
rect 3416 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3736 3840
rect 3416 2752 3736 3776
rect 3416 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3736 2752
rect 3416 2128 3736 2688
rect 5888 19616 6208 19632
rect 5888 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6208 19616
rect 5888 18528 6208 19552
rect 5888 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6208 18528
rect 5888 17440 6208 18464
rect 5888 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6208 17440
rect 5888 16352 6208 17376
rect 5888 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6208 16352
rect 5888 15264 6208 16288
rect 5888 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6208 15264
rect 5888 14176 6208 15200
rect 5888 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6208 14176
rect 5888 13088 6208 14112
rect 5888 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6208 13088
rect 5888 12000 6208 13024
rect 5888 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6208 12000
rect 5888 10912 6208 11936
rect 5888 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6208 10912
rect 5888 9824 6208 10848
rect 5888 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6208 9824
rect 5888 8736 6208 9760
rect 5888 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6208 8736
rect 5888 7648 6208 8672
rect 5888 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6208 7648
rect 5888 6560 6208 7584
rect 5888 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6208 6560
rect 5888 5472 6208 6496
rect 5888 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6208 5472
rect 5888 4384 6208 5408
rect 5888 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6208 4384
rect 5888 3296 6208 4320
rect 5888 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6208 3296
rect 5888 2208 6208 3232
rect 5888 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6208 2208
rect 5888 2128 6208 2144
rect 8361 19072 8681 19632
rect 8361 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8681 19072
rect 8361 17984 8681 19008
rect 8361 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8681 17984
rect 8361 16896 8681 17920
rect 8361 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8681 16896
rect 8361 15808 8681 16832
rect 8361 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8681 15808
rect 8361 14720 8681 15744
rect 8361 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8681 14720
rect 8361 13632 8681 14656
rect 8361 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8681 13632
rect 8361 12544 8681 13568
rect 8361 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8681 12544
rect 8361 11456 8681 12480
rect 8361 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8681 11456
rect 8361 10368 8681 11392
rect 8361 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8681 10368
rect 8361 9280 8681 10304
rect 8361 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8681 9280
rect 8361 8192 8681 9216
rect 8361 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8681 8192
rect 8361 7104 8681 8128
rect 8361 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8681 7104
rect 8361 6016 8681 7040
rect 8361 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8681 6016
rect 8361 4928 8681 5952
rect 8361 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8681 4928
rect 8361 3840 8681 4864
rect 8361 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8681 3840
rect 8361 2752 8681 3776
rect 8361 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8681 2752
rect 8361 2128 8681 2688
rect 10833 19616 11153 19632
rect 10833 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11153 19616
rect 10833 18528 11153 19552
rect 10833 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11153 18528
rect 10833 17440 11153 18464
rect 10833 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11153 17440
rect 10833 16352 11153 17376
rect 10833 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11153 16352
rect 10833 15264 11153 16288
rect 10833 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11153 15264
rect 10833 14176 11153 15200
rect 10833 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11153 14176
rect 10833 13088 11153 14112
rect 10833 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11153 13088
rect 10833 12000 11153 13024
rect 10833 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11153 12000
rect 10833 10912 11153 11936
rect 10833 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11153 10912
rect 10833 9824 11153 10848
rect 10833 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11153 9824
rect 10833 8736 11153 9760
rect 10833 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11153 8736
rect 10833 7648 11153 8672
rect 10833 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11153 7648
rect 10833 6560 11153 7584
rect 10833 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11153 6560
rect 10833 5472 11153 6496
rect 10833 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11153 5472
rect 10833 4384 11153 5408
rect 10833 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11153 4384
rect 10833 3296 11153 4320
rect 10833 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11153 3296
rect 10833 2208 11153 3232
rect 10833 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11153 2208
rect 10833 2128 11153 2144
rect 13306 19072 13626 19632
rect 13306 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13626 19072
rect 13306 17984 13626 19008
rect 13306 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13626 17984
rect 13306 16896 13626 17920
rect 13306 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13626 16896
rect 13306 15808 13626 16832
rect 13306 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13626 15808
rect 13306 14720 13626 15744
rect 13306 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13626 14720
rect 13306 13632 13626 14656
rect 13306 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13626 13632
rect 13306 12544 13626 13568
rect 13306 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13626 12544
rect 13306 11456 13626 12480
rect 13306 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13626 11456
rect 13306 10368 13626 11392
rect 13306 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13626 10368
rect 13306 9280 13626 10304
rect 13306 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13626 9280
rect 13306 8192 13626 9216
rect 13306 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13626 8192
rect 13306 7104 13626 8128
rect 13306 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13626 7104
rect 13306 6016 13626 7040
rect 13306 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13626 6016
rect 13306 4928 13626 5952
rect 13306 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13626 4928
rect 13306 3840 13626 4864
rect 13306 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13626 3840
rect 13306 2752 13626 3776
rect 13306 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13626 2752
rect 13306 2128 13626 2688
rect 15778 19616 16098 19632
rect 15778 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16098 19616
rect 15778 18528 16098 19552
rect 15778 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16098 18528
rect 15778 17440 16098 18464
rect 15778 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16098 17440
rect 15778 16352 16098 17376
rect 15778 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16098 16352
rect 15778 15264 16098 16288
rect 15778 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16098 15264
rect 15778 14176 16098 15200
rect 15778 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16098 14176
rect 15778 13088 16098 14112
rect 15778 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16098 13088
rect 15778 12000 16098 13024
rect 15778 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16098 12000
rect 15778 10912 16098 11936
rect 15778 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16098 10912
rect 15778 9824 16098 10848
rect 15778 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16098 9824
rect 15778 8736 16098 9760
rect 15778 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16098 8736
rect 15778 7648 16098 8672
rect 15778 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16098 7648
rect 15778 6560 16098 7584
rect 15778 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16098 6560
rect 15778 5472 16098 6496
rect 15778 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16098 5472
rect 15778 4384 16098 5408
rect 15778 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16098 4384
rect 15778 3296 16098 4320
rect 15778 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16098 3296
rect 15778 2208 16098 3232
rect 15778 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16098 2208
rect 15778 2128 16098 2144
rect 18251 19072 18571 19632
rect 18251 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18571 19072
rect 18251 17984 18571 19008
rect 18251 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18571 17984
rect 18251 16896 18571 17920
rect 18251 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18571 16896
rect 18251 15808 18571 16832
rect 18251 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18571 15808
rect 18251 14720 18571 15744
rect 18251 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18571 14720
rect 18251 13632 18571 14656
rect 18251 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18571 13632
rect 18251 12544 18571 13568
rect 18251 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18571 12544
rect 18251 11456 18571 12480
rect 18251 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18571 11456
rect 18251 10368 18571 11392
rect 18251 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18571 10368
rect 18251 9280 18571 10304
rect 18251 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18571 9280
rect 18251 8192 18571 9216
rect 18251 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18571 8192
rect 18251 7104 18571 8128
rect 18251 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18571 7104
rect 18251 6016 18571 7040
rect 18251 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18571 6016
rect 18251 4928 18571 5952
rect 18251 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18571 4928
rect 18251 3840 18571 4864
rect 18251 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18571 3840
rect 18251 2752 18571 3776
rect 18251 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18571 2752
rect 18251 2128 18571 2688
rect 20723 19616 21043 19632
rect 20723 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21043 19616
rect 20723 18528 21043 19552
rect 20723 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21043 18528
rect 20723 17440 21043 18464
rect 20723 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21043 17440
rect 20723 16352 21043 17376
rect 20723 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21043 16352
rect 20723 15264 21043 16288
rect 20723 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21043 15264
rect 20723 14176 21043 15200
rect 20723 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21043 14176
rect 20723 13088 21043 14112
rect 20723 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21043 13088
rect 20723 12000 21043 13024
rect 20723 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21043 12000
rect 20723 10912 21043 11936
rect 20723 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21043 10912
rect 20723 9824 21043 10848
rect 20723 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21043 9824
rect 20723 8736 21043 9760
rect 20723 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21043 8736
rect 20723 7648 21043 8672
rect 20723 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21043 7648
rect 20723 6560 21043 7584
rect 20723 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21043 6560
rect 20723 5472 21043 6496
rect 20723 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21043 5472
rect 20723 4384 21043 5408
rect 20723 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21043 4384
rect 20723 3296 21043 4320
rect 20723 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21043 3296
rect 20723 2208 21043 3232
rect 20723 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21043 2208
rect 20723 2128 21043 2144
use sky130_fd_sc_hd__decap_3  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99
timestamp 1676037725
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_157
timestamp 1676037725
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp 1676037725
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_186
timestamp 1676037725
transform 1 0 18216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1676037725
transform 1 0 19780 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_210
timestamp 1676037725
transform 1 0 20424 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_119
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_130
timestamp 1676037725
transform 1 0 13064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_142
timestamp 1676037725
transform 1 0 14168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_154
timestamp 1676037725
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_211
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_44
timestamp 1676037725
transform 1 0 5152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1676037725
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1676037725
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1676037725
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_107
timestamp 1676037725
transform 1 0 10948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_120
timestamp 1676037725
transform 1 0 12144 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_126
timestamp 1676037725
transform 1 0 12696 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_149
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_161
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_173
timestamp 1676037725
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_185
timestamp 1676037725
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_12
timestamp 1676037725
transform 1 0 2208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_18
timestamp 1676037725
transform 1 0 2760 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_22
timestamp 1676037725
transform 1 0 3128 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_34
timestamp 1676037725
transform 1 0 4232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1676037725
transform 1 0 5336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_50
timestamp 1676037725
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1676037725
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1676037725
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_74
timestamp 1676037725
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_86
timestamp 1676037725
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_98
timestamp 1676037725
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_118
timestamp 1676037725
transform 1 0 11960 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_130
timestamp 1676037725
transform 1 0 13064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_143
timestamp 1676037725
transform 1 0 14260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_211
timestamp 1676037725
transform 1 0 20516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_16
timestamp 1676037725
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1676037725
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_60
timestamp 1676037725
transform 1 0 6624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_68
timestamp 1676037725
transform 1 0 7360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1676037725
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_100
timestamp 1676037725
transform 1 0 10304 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_108
timestamp 1676037725
transform 1 0 11040 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_120
timestamp 1676037725
transform 1 0 12144 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1676037725
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1676037725
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_183
timestamp 1676037725
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1676037725
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_36
timestamp 1676037725
transform 1 0 4416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp 1676037725
transform 1 0 5244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1676037725
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1676037725
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1676037725
transform 1 0 8372 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1676037725
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_99
timestamp 1676037725
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_103
timestamp 1676037725
transform 1 0 10580 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_123
timestamp 1676037725
transform 1 0 12420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_131
timestamp 1676037725
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_140
timestamp 1676037725
transform 1 0 13984 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_152
timestamp 1676037725
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1676037725
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_176
timestamp 1676037725
transform 1 0 17296 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_185
timestamp 1676037725
transform 1 0 18124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_200
timestamp 1676037725
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_51
timestamp 1676037725
transform 1 0 5796 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_61
timestamp 1676037725
transform 1 0 6716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1676037725
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_103
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_111
timestamp 1676037725
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1676037725
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_152
timestamp 1676037725
transform 1 0 15088 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_164
timestamp 1676037725
transform 1 0 16192 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1676037725
transform 1 0 16928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1676037725
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1676037725
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_18
timestamp 1676037725
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_30
timestamp 1676037725
transform 1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1676037725
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_42
timestamp 1676037725
transform 1 0 4968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1676037725
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1676037725
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_133
timestamp 1676037725
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1676037725
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1676037725
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1676037725
transform 1 0 17572 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_200
timestamp 1676037725
transform 1 0 19504 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1676037725
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_43
timestamp 1676037725
transform 1 0 5060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_51
timestamp 1676037725
transform 1 0 5796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1676037725
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1676037725
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_112
timestamp 1676037725
transform 1 0 11408 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1676037725
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_150
timestamp 1676037725
transform 1 0 14904 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_162
timestamp 1676037725
transform 1 0 16008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1676037725
transform 1 0 16744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1676037725
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1676037725
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1676037725
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1676037725
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_75
timestamp 1676037725
transform 1 0 8004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1676037725
transform 1 0 8740 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_90
timestamp 1676037725
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1676037725
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_104
timestamp 1676037725
transform 1 0 10672 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_120
timestamp 1676037725
transform 1 0 12144 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_138
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_162
timestamp 1676037725
transform 1 0 16008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_179
timestamp 1676037725
transform 1 0 17572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_195
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_201
timestamp 1676037725
transform 1 0 19596 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_209
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1676037725
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_36
timestamp 1676037725
transform 1 0 4416 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_60
timestamp 1676037725
transform 1 0 6624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1676037725
transform 1 0 6992 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1676037725
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_90
timestamp 1676037725
transform 1 0 9384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_110
timestamp 1676037725
transform 1 0 11224 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1676037725
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1676037725
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_149
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_159
timestamp 1676037725
transform 1 0 15732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1676037725
transform 1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_178
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_205
timestamp 1676037725
transform 1 0 19964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_211
timestamp 1676037725
transform 1 0 20516 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1676037725
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_88
timestamp 1676037725
transform 1 0 9200 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_154
timestamp 1676037725
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1676037725
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_185
timestamp 1676037725
transform 1 0 18124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_197
timestamp 1676037725
transform 1 0 19228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_211
timestamp 1676037725
transform 1 0 20516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1676037725
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1676037725
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1676037725
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_71
timestamp 1676037725
transform 1 0 7636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1676037725
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1676037725
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_156
timestamp 1676037725
transform 1 0 15456 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1676037725
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_211
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_16
timestamp 1676037725
transform 1 0 2576 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1676037725
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_43
timestamp 1676037725
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_94
timestamp 1676037725
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1676037725
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_177
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1676037725
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_203
timestamp 1676037725
transform 1 0 19780 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_211
timestamp 1676037725
transform 1 0 20516 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_13
timestamp 1676037725
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1676037725
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_63
timestamp 1676037725
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1676037725
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_157
timestamp 1676037725
transform 1 0 15548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_178
timestamp 1676037725
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_10
timestamp 1676037725
transform 1 0 2024 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_22
timestamp 1676037725
transform 1 0 3128 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1676037725
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_75
timestamp 1676037725
transform 1 0 8004 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_87
timestamp 1676037725
transform 1 0 9108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_99
timestamp 1676037725
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1676037725
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_138
timestamp 1676037725
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_150
timestamp 1676037725
transform 1 0 14904 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_182
timestamp 1676037725
transform 1 0 17848 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_12
timestamp 1676037725
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1676037725
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_50
timestamp 1676037725
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1676037725
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1676037725
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1676037725
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1676037725
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1676037725
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_206
timestamp 1676037725
transform 1 0 20056 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1676037725
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_12
timestamp 1676037725
transform 1 0 2208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_24
timestamp 1676037725
transform 1 0 3312 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_32
timestamp 1676037725
transform 1 0 4048 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1676037725
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_96
timestamp 1676037725
transform 1 0 9936 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1676037725
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1676037725
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_186
timestamp 1676037725
transform 1 0 18216 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_202
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1676037725
transform 1 0 20424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_14
timestamp 1676037725
transform 1 0 2392 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1676037725
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_69
timestamp 1676037725
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1676037725
transform 1 0 20056 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1676037725
transform 1 0 3312 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1676037725
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_75
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1676037725
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1676037725
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_136
timestamp 1676037725
transform 1 0 13616 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_148
timestamp 1676037725
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_179
timestamp 1676037725
transform 1 0 17572 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_187
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1676037725
transform 1 0 20516 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1676037725
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_50
timestamp 1676037725
transform 1 0 5704 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_62
timestamp 1676037725
transform 1 0 6808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_111
timestamp 1676037725
transform 1 0 11316 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_119
timestamp 1676037725
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1676037725
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1676037725
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1676037725
transform 1 0 20148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1676037725
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_16
timestamp 1676037725
transform 1 0 2576 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_28
timestamp 1676037725
transform 1 0 3680 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_40
timestamp 1676037725
transform 1 0 4784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1676037725
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_77
timestamp 1676037725
transform 1 0 8188 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_98
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_131
timestamp 1676037725
transform 1 0 13156 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_143
timestamp 1676037725
transform 1 0 14260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_156
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1676037725
transform 1 0 19412 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_203
timestamp 1676037725
transform 1 0 19780 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1676037725
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_13
timestamp 1676037725
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1676037725
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1676037725
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_156
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_168
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_174
timestamp 1676037725
transform 1 0 17112 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_180
timestamp 1676037725
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1676037725
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1676037725
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_13
timestamp 1676037725
transform 1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1676037725
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1676037725
transform 1 0 4232 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_92
timestamp 1676037725
transform 1 0 9568 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1676037725
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_136
timestamp 1676037725
transform 1 0 13616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_146
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_183
timestamp 1676037725
transform 1 0 17940 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_204
timestamp 1676037725
transform 1 0 19872 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_14
timestamp 1676037725
transform 1 0 2392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1676037725
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1676037725
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_105
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_117
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_156
timestamp 1676037725
transform 1 0 15456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_176
timestamp 1676037725
transform 1 0 17296 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1676037725
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1676037725
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1676037725
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_211
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1676037725
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_14
timestamp 1676037725
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1676037725
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1676037725
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_131
timestamp 1676037725
transform 1 0 13156 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_143
timestamp 1676037725
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_155
timestamp 1676037725
transform 1 0 15364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_192
timestamp 1676037725
transform 1 0 18768 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_198
timestamp 1676037725
transform 1 0 19320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1676037725
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_12
timestamp 1676037725
transform 1 0 2208 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1676037725
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_48
timestamp 1676037725
transform 1 0 5520 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1676037725
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_164
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_172
timestamp 1676037725
transform 1 0 16928 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_184
timestamp 1676037725
transform 1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_204
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_14
timestamp 1676037725
transform 1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_23
timestamp 1676037725
transform 1 0 3220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1676037725
transform 1 0 9016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1676037725
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1676037725
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_153
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_176
timestamp 1676037725
transform 1 0 17296 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_184
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1676037725
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1676037725
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_63
timestamp 1676037725
transform 1 0 6900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_105
timestamp 1676037725
transform 1 0 10764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1676037725
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1676037725
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1676037725
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_169
timestamp 1676037725
transform 1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1676037725
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_16
timestamp 1676037725
transform 1 0 2576 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1676037725
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_134
timestamp 1676037725
transform 1 0 13432 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_141
timestamp 1676037725
transform 1 0 14076 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1676037725
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1676037725
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_209
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 20884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1676037725
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1676037725
transform 1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1676037725
transform 1 0 16376 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1676037725
transform -1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 3036 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _193_
timestamp 1676037725
transform 1 0 1748 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19136 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _198_
timestamp 1676037725
transform -1 0 19780 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp 1676037725
transform 1 0 14996 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _201_
timestamp 1676037725
transform 1 0 14996 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 13340 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1676037725
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _204_
timestamp 1676037725
transform 1 0 17756 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1676037725
transform 1 0 19412 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14628 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16192 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15732 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _209_
timestamp 1676037725
transform 1 0 14904 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _210_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16652 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _212_
timestamp 1676037725
transform -1 0 15824 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _213_
timestamp 1676037725
transform -1 0 17572 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1676037725
transform -1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16652 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _218_
timestamp 1676037725
transform -1 0 17388 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__o21ai_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15456 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _225_
timestamp 1676037725
transform -1 0 16192 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _229_
timestamp 1676037725
transform -1 0 13984 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _231_
timestamp 1676037725
transform -1 0 15548 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _233_
timestamp 1676037725
transform -1 0 15916 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 1676037725
transform -1 0 3404 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1676037725
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp 1676037725
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _239_
timestamp 1676037725
transform 1 0 4784 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _240_
timestamp 1676037725
transform 1 0 7452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_4  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8004 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1676037725
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17940 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8464 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 4416 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 6900 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_2  _248_
timestamp 1676037725
transform -1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 8648 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _250_
timestamp 1676037725
transform 1 0 7268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _251_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp 1676037725
transform -1 0 5336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1676037725
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _257_
timestamp 1676037725
transform 1 0 5152 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5060 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1676037725
transform -1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _260_
timestamp 1676037725
transform -1 0 8004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _261_
timestamp 1676037725
transform -1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1676037725
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _263_
timestamp 1676037725
transform -1 0 7084 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _265_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2208 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _267_
timestamp 1676037725
transform -1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _268_
timestamp 1676037725
transform -1 0 2576 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1676037725
transform -1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _270_
timestamp 1676037725
transform 1 0 9568 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13340 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _272_
timestamp 1676037725
transform -1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _273_
timestamp 1676037725
transform 1 0 12788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _274_
timestamp 1676037725
transform -1 0 13340 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _275_
timestamp 1676037725
transform -1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10580 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _277_
timestamp 1676037725
transform 1 0 11500 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _278_
timestamp 1676037725
transform -1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _279_
timestamp 1676037725
transform 1 0 10672 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 1676037725
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 10304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _284_
timestamp 1676037725
transform -1 0 12328 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _286_
timestamp 1676037725
transform 1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _287_
timestamp 1676037725
transform 1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _288_
timestamp 1676037725
transform -1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _289_
timestamp 1676037725
transform -1 0 12144 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1676037725
transform -1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _291_
timestamp 1676037725
transform -1 0 11224 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _292_
timestamp 1676037725
transform -1 0 18492 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _293_
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _295_
timestamp 1676037725
transform -1 0 19872 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 1676037725
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _297_
timestamp 1676037725
transform 1 0 16836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17572 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _299_
timestamp 1676037725
transform 1 0 17664 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _300_
timestamp 1676037725
transform -1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _301_
timestamp 1676037725
transform -1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _302_
timestamp 1676037725
transform 1 0 17020 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1676037725
transform 1 0 17848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _304_
timestamp 1676037725
transform -1 0 17572 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _305_
timestamp 1676037725
transform -1 0 17388 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _306_
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _307_
timestamp 1676037725
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _308_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17664 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _309_
timestamp 1676037725
transform -1 0 17388 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _310_
timestamp 1676037725
transform 1 0 17020 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _311_
timestamp 1676037725
transform -1 0 17572 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _312_
timestamp 1676037725
transform -1 0 18952 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp 1676037725
transform -1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _314_
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _315_
timestamp 1676037725
transform 1 0 18400 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _316_
timestamp 1676037725
transform 1 0 18308 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _317_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp 1676037725
transform 1 0 18400 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _319_
timestamp 1676037725
transform -1 0 19688 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _320_
timestamp 1676037725
transform -1 0 20056 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _321_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _323_
timestamp 1676037725
transform 1 0 19228 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _324_
timestamp 1676037725
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _325_
timestamp 1676037725
transform -1 0 20148 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1676037725
transform 1 0 18308 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _327_
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _328_
timestamp 1676037725
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 1676037725
transform -1 0 17204 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _330_
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _331_
timestamp 1676037725
transform -1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _332_
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _334_
timestamp 1676037725
transform -1 0 19872 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _335_
timestamp 1676037725
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _336_
timestamp 1676037725
transform 1 0 17020 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 17296 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 16928 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _340_
timestamp 1676037725
transform 1 0 14260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1676037725
transform -1 0 15732 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _342_
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _343_
timestamp 1676037725
transform 1 0 1932 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _344_
timestamp 1676037725
transform 1 0 2852 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _345_
timestamp 1676037725
transform 1 0 1932 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _346_
timestamp 1676037725
transform -1 0 2576 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _348_
timestamp 1676037725
transform -1 0 15088 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _349_
timestamp 1676037725
transform 1 0 14720 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _350_
timestamp 1676037725
transform 1 0 15548 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _351_
timestamp 1676037725
transform -1 0 15180 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _352_
timestamp 1676037725
transform 1 0 2760 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _353_
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _354_
timestamp 1676037725
transform -1 0 2576 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _355_
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1676037725
transform 1 0 1840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _357_
timestamp 1676037725
transform -1 0 2392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _358_
timestamp 1676037725
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _359_
timestamp 1676037725
transform -1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _360_
timestamp 1676037725
transform 1 0 2024 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _361_
timestamp 1676037725
transform 1 0 1840 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5244 0 -1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _364_
timestamp 1676037725
transform -1 0 5704 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5060 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1676037725
transform 1 0 4140 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 1676037725
transform -1 0 4968 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1676037725
transform 1 0 7176 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1676037725
transform 1 0 7176 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1676037725
transform 1 0 7728 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1676037725
transform 1 0 6532 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _372_
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1676037725
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _374_
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _375_
timestamp 1676037725
transform -1 0 10488 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _376_
timestamp 1676037725
transform 1 0 9568 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _377_
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1676037725
transform 1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _379_
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1676037725
transform 1 0 9752 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _381_
timestamp 1676037725
transform 1 0 9200 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1676037725
transform 1 0 12236 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _388_
timestamp 1676037725
transform 1 0 12144 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1676037725
transform 1 0 12144 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _390_
timestamp 1676037725
transform 1 0 12052 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _394_
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _397_
timestamp 1676037725
transform -1 0 5704 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _398_
timestamp 1676037725
transform -1 0 5428 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _399_
timestamp 1676037725
transform -1 0 5520 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1676037725
transform -1 0 5244 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _401_
timestamp 1676037725
transform -1 0 8464 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _402_
timestamp 1676037725
transform 1 0 9292 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _403_
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _404_
timestamp 1676037725
transform 1 0 7544 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _405_
timestamp 1676037725
transform 1 0 9384 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _406_
timestamp 1676037725
transform 1 0 5888 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1676037725
transform -1 0 5428 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1676037725
transform -1 0 6072 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1676037725
transform -1 0 4232 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1676037725
transform -1 0 5152 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _411_
timestamp 1676037725
transform -1 0 8004 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _412_
timestamp 1676037725
transform -1 0 6716 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _413_
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _414_
timestamp 1676037725
transform 1 0 5428 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1676037725
transform 1 0 5152 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8280 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1676037725
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1676037725
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1676037725
transform 1 0 10396 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1676037725
transform 1 0 19504 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 18308 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1676037725
transform 1 0 15180 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1676037725
transform -1 0 15548 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1676037725
transform 1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1676037725
transform -1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1676037725
transform -1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output3
timestamp 1676037725
transform -1 0 2208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1676037725
transform -1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1676037725
transform -1 0 7544 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1676037725
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp 1676037725
transform 1 0 17664 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp 1676037725
transform 1 0 19872 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal2 s 3698 21200 3754 22000 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 18234 21200 18290 22000 0 FreeSans 224 90 0 0 io_in
port 1 nsew signal input
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 io_out[0]
port 2 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 io_out[1]
port 3 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 io_out[2]
port 4 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 io_out[3]
port 5 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_out[4]
port 6 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 io_out[5]
port 7 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 io_out[6]
port 8 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 io_out[7]
port 9 nsew signal tristate
flabel metal2 s 10966 21200 11022 22000 0 FreeSans 224 90 0 0 rst
port 10 nsew signal input
flabel metal4 s 3416 2128 3736 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 8361 2128 8681 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 13306 2128 13626 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 18251 2128 18571 19632 0 FreeSans 1920 90 0 0 vccd1
port 11 nsew power bidirectional
flabel metal4 s 5888 2128 6208 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 10833 2128 11153 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 15778 2128 16098 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
flabel metal4 s 20723 2128 21043 19632 0 FreeSans 1920 90 0 0 vssd1
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22000 22000
<< end >>
