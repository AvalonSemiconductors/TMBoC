magic
tech sky130B
magscale 1 2
timestamp 1682098769
<< obsli1 >>
rect 1104 2159 20884 19601
<< obsm1 >>
rect 1104 2128 21043 19632
<< obsm2 >>
rect 1584 2139 21037 19621
<< metal3 >>
rect 0 18232 800 18352
rect 0 10888 800 11008
rect 0 3544 800 3664
<< obsm3 >>
rect 800 18432 21041 19617
rect 880 18152 21041 18432
rect 800 11088 21041 18152
rect 880 10808 21041 11088
rect 800 3744 21041 10808
rect 880 3464 21041 3744
rect 800 2143 21041 3464
<< metal4 >>
rect 3416 2128 3736 19632
rect 5888 2128 6208 19632
rect 8361 2128 8681 19632
rect 10833 2128 11153 19632
rect 13306 2128 13626 19632
rect 15778 2128 16098 19632
rect 18251 2128 18571 19632
rect 20723 2128 21043 19632
<< labels >>
rlabel metal3 s 0 18232 800 18352 6 OP
port 1 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 clk
port 2 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 rst
port 3 nsew signal input
rlabel metal4 s 3416 2128 3736 19632 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 8361 2128 8681 19632 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 13306 2128 13626 19632 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 18251 2128 18571 19632 6 vccd1
port 4 nsew power bidirectional
rlabel metal4 s 5888 2128 6208 19632 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 10833 2128 11153 19632 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 15778 2128 16098 19632 6 vssd1
port 5 nsew ground bidirectional
rlabel metal4 s 20723 2128 21043 19632 6 vssd1
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 22000 22000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1349658
string GDS_FILE /run/media/tholin/Data/Projects/MPW/TMBoC/openlane/TunePlayer/runs/23_04_21_19_38/results/signoff/tune_player.magic.gds
string GDS_START 549934
<< end >>

