* NGSPICE file created from tholin_avalonsemi_5401.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt tholin_avalonsemi_5401 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] rst vccd1
+ vssd1
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0985_ _0501_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_24.result sky130_fd_sc_hd__buf_1
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1115__B1 _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0770_ _0305_ _0308_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__and2_1
XANTENNA__1106__B1 _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1184_ net45 _0058_ vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0968_ CIRCUIT_1957.MEMORY_66.s_currentState _0469_ CIRCUIT_1957.MEMORY_62.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__mux2_1
X_0899_ _0292_ _0375_ _0431_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0822_ _0353_ _0299_ _0358_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0684_ _0211_ _0212_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__nor2_1
X_0753_ _0291_ _0277_ _0288_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__a21o_2
X_1098_ CIRCUIT_1957.int_memory_1.mul2_1.A2 _0532_ _0514_ vssd1 vssd1 vccd1 vccd1
+ _0079_ sky130_fd_sc_hd__a21o_1
X_1167_ CIRCUIT_1957.GATES_41.result CIRCUIT_1957.GATES_28.result _0011_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_73.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1030__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__clkbuf_4
X_0805_ _0337_ _0169_ _0339_ _0340_ _0343_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__a41o_1
X_0598_ net7 net3 _0144_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__mux2_1
X_0667_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A3 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__nor2_1
X_0736_ _0273_ _0274_ _0231_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__a21o_1
X_1219_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result _0093_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.B0 sky130_fd_sc_hd__dfxtp_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1004_ clknet_1_0__leaf_clk _0119_ _0341_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__and3_2
X_0719_ _0233_ _0246_ _0257_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__a21oi_2
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__0502_ clknet_0__0502_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0502_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0984_ clknet_1_1__leaf__0498_ _0496_ _0321_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__and3_2
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0874__B1 _0333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result
+ sky130_fd_sc_hd__clkbuf_16
X_1183_ net44 _0057_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1042__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0967_ _0491_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_30.result sky130_fd_sc_hd__dlymetal6s2s_1
X_0898_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[0\] _0333_ _0341_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[0\]
+ _0436_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__a221o_1
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1033__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0821_ _0359_ _0309_ _0348_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__o21a_1
X_0752_ _0281_ _0282_ _0168_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__a21o_1
XANTENNA__1024__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0683_ _0200_ _0221_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__xor2_2
X_1166_ CIRCUIT_1957.GATES_41.result CIRCUIT_1957.GATES_30.result _0010_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_74.s_currentState sky130_fd_sc_hd__dfrtp_1
X_1097_ _0511_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__buf_2
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1015__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1020_ _0521_ _0511_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__nor2_2
X_0735_ _0272_ _0258_ _0259_ _0267_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__nand4_1
X_0804_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[3\] _0341_ _0342_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a22o_1
X_0597_ _0146_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.D1 sky130_fd_sc_hd__clkbuf_1
X_0666_ _0202_ _0204_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1218_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result _0092_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A7 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1149_ CIRCUIT_1957.clock_gen_2_1.CLK1 CIRCUIT_1957.D1 _0005_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState sky130_fd_sc_hd__dfrtp_4
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result CIRCUIT_1957.int_memory_1.GATES_21.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result sky130_fd_sc_hd__clkbuf_16
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1003_ _0509_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_50.result sky130_fd_sc_hd__buf_1
X_0718_ _0166_ _0246_ CIRCUIT_1957.int_memory_1.div_1.A2 vssd1 vssd1 vccd1 vccd1 _0257_
+ sky130_fd_sc_hd__a21boi_1
X_0649_ _0175_ _0186_ _0187_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__mux2_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0598__S _0144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1073__8 clknet_1_1__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__inv_2
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0983_ _0500_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_23.result sky130_fd_sc_hd__buf_1
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0580__A0 CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1115__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result
+ sky130_fd_sc_hd__clkbuf_16
X_1182_ net43 _0056_ vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0897_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[0\] _0334_ _0433_ _0435_ vssd1 vssd1
+ vccd1 vccd1 _0436_ sky130_fd_sc_hd__a211o_1
X_0966_ CIRCUIT_1957.MEMORY_67.s_currentState _0398_ CIRCUIT_1957.MEMORY_62.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__mux2_1
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0820_ CIRCUIT_1957.int_memory_1.mul2_1.A3 CIRCUIT_1957.int_memory_1.mul2_1.B1 vssd1
+ vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__and2_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0751_ _0281_ _0282_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__nand2_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0682_ _0215_ _0219_ _0220_ _0208_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__a211o_1
X_1096_ CIRCUIT_1957.int_memory_1.mul2_1.A1 _0531_ _0523_ vssd1 vssd1 vccd1 vccd1
+ _0078_ sky130_fd_sc_hd__a21o_1
X_1165_ CIRCUIT_1957.GATES_41.result CIRCUIT_1957.GATES_35.result _0009_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_75.s_currentState sky130_fd_sc_hd__dfrtp_1
X_0949_ _0482_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.clock_gen_2_1.GATES_3.result sky130_fd_sc_hd__clkbuf_1
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0665_ _0188_ _0203_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__xor2_1
X_0803_ _0295_ _0319_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__nor2_1
X_0734_ _0272_ _0259_ _0267_ _0258_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__a31o_1
Xclkbuf_1_0__f__0526_ clknet_0__0526_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0526_
+ sky130_fd_sc_hd__clkbuf_16
X_0596_ net6 net2 _0144_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__mux2_1
X_1217_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result _0091_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A6 sky130_fd_sc_hd__dfxtp_1
X_1079_ _0527_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
X_1148_ CIRCUIT_1957.clock_gen_2_1.CLK1 CIRCUIT_1957.D0 _0004_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1002_ clknet_1_1__leaf__0498_ _0119_ _0342_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__and3_2
X_0648_ _0173_ _0176_ _0182_ _0181_ _0168_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__a32o_1
X_0717_ _0162_ _0255_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__and2_1
X_0579_ _0135_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0968__A0 CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1118__B1 _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0982_ clknet_1_1__leaf__0498_ _0496_ _0333_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__and3_2
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1181_ net42 _0055_ vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__0502_ _0502_ vssd1 vssd1 vccd1 vccd1 clknet_0__0502_ sky130_fd_sc_hd__clkbuf_16
X_0965_ _0490_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_35.result sky130_fd_sc_hd__dlymetal6s2s_1
X_0896_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[0\] _0328_ _0342_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[0\]
+ _0434_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__a221o_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1033__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0681_ _0207_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
X_0750_ _0277_ _0288_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__and2b_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1095_ CIRCUIT_1957.int_memory_1.mul2_1.A0 _0531_ _0520_ vssd1 vssd1 vccd1 vccd1
+ _0077_ sky130_fd_sc_hd__a21o_1
X_1164_ CIRCUIT_1957.GATES_39.result CIRCUIT_1957.GATES_27.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_76.s_currentState sky130_fd_sc_hd__dfxtp_1
X_0948_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState vssd1 vssd1 vccd1 vccd1
+ _0482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0879_ _0409_ _0415_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__or3_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0802_ _0324_ _0319_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__nor2_1
X_0664_ _0185_ _0189_ _0197_ _0198_ CIRCUIT_1957.int_memory_1.div_1.B2 vssd1 vssd1
+ vccd1 vccd1 _0203_ sky130_fd_sc_hd__o311a_1
X_0733_ _0162_ _0255_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__nand2_1
X_0595_ _0145_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.D0 sky130_fd_sc_hd__clkbuf_1
X_1216_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result _0090_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A5 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result CIRCUIT_1957.int_memory_1.GATES_50.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result sky130_fd_sc_hd__clkbuf_16
X_1078_ net25 net11 vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__or2_1
X_1147_ _0003_ CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 _0002_ vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1001_ _0508_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_33.result sky130_fd_sc_hd__buf_1
XANTENNA__1000__A clknet_1_0__leaf__0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0647_ _0171_ _0176_ _0172_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__a21o_1
X_0716_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A1 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__nor2_1
X_0578_ net26 net15 _0108_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__mux2_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1090__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_2
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A io_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0981_ _0499_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_22.result sky130_fd_sc_hd__buf_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1045__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result CIRCUIT_1957.int_memory_1.GATES_27.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result sky130_fd_sc_hd__clkbuf_16
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1036__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1180_ net41 _0054_ vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1027__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0617__A3 _0149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0964_ CIRCUIT_1957.MEMORY_63.s_currentState _0378_ CIRCUIT_1957.MEMORY_62.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__mux2_1
X_0895_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[0\] _0323_ _0332_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__a22o_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1018__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0680_ _0167_ _0205_ _0218_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__o21a_1
X_1094_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[3\] _0531_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0076_ sky130_fd_sc_hd__a21o_1
X_1163_ CIRCUIT_1957.GATES_39.result CIRCUIT_1957.GATES_28.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_77.s_currentState sky130_fd_sc_hd__dfxtp_1
X_0947_ _0478_ _0480_ _0481_ _0458_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.MEMORY_63.d
+ sky130_fd_sc_hd__a2bb2o_1
X_0878_ _0347_ _0416_ _0339_ _0187_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__a2bb2o_1
Xtholin_avalonsemi_5401_30 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_30/HI io_out[6]
+ sky130_fd_sc_hd__conb_1
X_0801_ _0166_ _0177_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__nand2_1
X_0594_ net5 net1 _0144_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0663_ _0191_ _0196_ _0201_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__or3_1
X_0732_ _0165_ _0268_ _0269_ _0270_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__o31a_1
X_1215_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result _0089_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A4 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1146_ clknet_1_0__leaf_clk CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d _0001_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState sky130_fd_sc_hd__dfrtp_4
X_1077_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[3\] _0525_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0064_ sky130_fd_sc_hd__a21o_1
XFILLER_29_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ clknet_1_0__leaf__0498_ _0119_ _0331_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__and3_2
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1000__B _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0715_ _0231_ _0253_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__nand2_1
X_0646_ _0168_ _0184_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__and2_1
X_0577_ _0134_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1129_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result _0037_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_6.input2\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_2
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_2
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0629_ CIRCUIT_1957.int_memory_1.div_1.B3 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1118__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0980_ clknet_1_0__leaf__0498_ _0496_ _0334_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__and3_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1109__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0859__B2 _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0963_ _0489_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_38.result sky130_fd_sc_hd__clkbuf_1
X_0894_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[0\] _0327_ _0325_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[0\]
+ _0432_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__a221o_1
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result CIRCUIT_1957.int_memory_1.GATES_33.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result sky130_fd_sc_hd__clkbuf_16
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1162_ CIRCUIT_1957.GATES_39.result CIRCUIT_1957.GATES_30.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_78.s_currentState sky130_fd_sc_hd__dfxtp_1
X_1093_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[2\] _0531_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0075_ sky130_fd_sc_hd__a21o_1
X_0877_ _0363_ _0370_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0946_ _0400_ _0456_ _0457_ _0459_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o31a_1
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtholin_avalonsemi_5401_31 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_31/HI io_out[7]
+ sky130_fd_sc_hd__conb_1
X_0800_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
X_0731_ _0162_ _0164_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__or2_1
X_0662_ _0185_ _0189_ _0197_ _0198_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__o31ai_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0593_ net22 net25 net24 net21 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__or4b_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1014__A _0517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1214_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result _0088_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A3 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1145_ CIRCUIT_1957.clock_gen_2_1.GATES_3.result CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
+ _0000_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState
+ sky130_fd_sc_hd__dfstp_1
X_1076_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[2\] _0525_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0063_ sky130_fd_sc_hd__a21o_1
X_0929_ _0465_ _0449_ _0466_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1000__C _0331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0645_ _0173_ _0176_ _0182_ _0183_ _0177_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__a311oi_2
X_0714_ _0236_ _0252_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__xnor2_2
X_0576_ CIRCUIT_1957.MEMORY_67.s_currentState CIRCUIT_1957.MEMORY_70.s_currentState
+ CIRCUIT_1957.MEMORY_86.s_currentState CIRCUIT_1957.MEMORY_78.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__mux4_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1059_ _0140_ clknet_1_0__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__nand2_2
X_1128_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result _0036_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_5.input2\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_2
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_2
XFILLER_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0628_ CIRCUIT_1957.int_memory_1.div_1.B3 vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0559_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState _0099_ _0120_ vssd1 vssd1
+ vccd1 vccd1 _0121_ sky130_fd_sc_hd__or3b_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0861__A CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1036__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0893_ CIRCUIT_1957.int_memory_1.mul2_1.A0 CIRCUIT_1957.int_memory_1.mul2_1.B0 _0321_
+ _0331_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[0\] vssd1 vssd1 vccd1 vccd1 _0432_
+ sky130_fd_sc_hd__a32o_1
X_0962_ _0128_ _0120_ _0149_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__and3_1
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1092_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[1\] _0531_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0074_ sky130_fd_sc_hd__a21o_1
X_1161_ CIRCUIT_1957.GATES_39.result CIRCUIT_1957.GATES_35.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_79.s_currentState sky130_fd_sc_hd__dfxtp_1
X_0876_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[1\] _0327_ _0341_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[1\]
+ _0414_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__a221o_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0945_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState CIRCUIT_1957.MEMORY_63.s_currentState
+ _0378_ _0459_ _0479_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__a311o_1
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtholin_avalonsemi_5401_32 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_32/HI io_out[8]
+ sky130_fd_sc_hd__conb_1
X_0661_ CIRCUIT_1957.int_memory_1.div_1.A4 _0199_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__xor2_2
X_0730_ _0166_ _0267_ CIRCUIT_1957.int_memory_1.div_1.A1 vssd1 vssd1 vccd1 vccd1 _0269_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1213_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result _0087_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A2 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1084__A_N net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0592_ _0141_ clknet_1_1__leaf__0143_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__nand2_2
X_1075_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[1\] _0525_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0062_ sky130_fd_sc_hd__a21o_1
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result _0052_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_49.input2\[3\] sky130_fd_sc_hd__dfxtp_1
X_0928_ _0465_ _0449_ _0459_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__o21ai_1
X_0859_ _0115_ CIRCUIT_1957.D2 _0397_ _0119_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__a22o_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1093__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1066__1 clknet_1_0__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__inv_2
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0644_ _0178_ _0169_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__and2b_1
X_0713_ _0234_ _0237_ _0246_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__nand3b_1
XANTENNA__1009__B _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0575_ _0133_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__1075__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1058_ _0140_ clknet_1_0__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__nand2_2
X_1127_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result _0035_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_5.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_2
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_2
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0627_ CIRCUIT_1957.int_memory_1.div_1.B0 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__buf_2
X_0558_ CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__nor2_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1039__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input6_A io_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0961_ _0488_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_39.result sky130_fd_sc_hd__clkbuf_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0892_ _0201_ _0338_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__nor2_1
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0940__A2 CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1091_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[0\] _0531_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0073_ sky130_fd_sc_hd__a21o_1
X_1160_ CIRCUIT_1957.GATES_40.result CIRCUIT_1957.GATES_27.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_80.s_currentState sky130_fd_sc_hd__dfxtp_1
X_0944_ _0099_ _0378_ _0161_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__a21oi_1
X_0875_ _0410_ _0321_ _0411_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__a31o_1
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result
+ sky130_fd_sc_hd__clkbuf_16
Xtholin_avalonsemi_5401_33 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_33/HI io_out[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0660_ _0185_ _0189_ _0197_ _0198_ _0166_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__o311a_1
X_0591_ clknet_1_0__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__buf_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1212_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result _0086_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1074_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[0\] _0525_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0061_ sky130_fd_sc_hd__a21o_1
X_1143_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result _0051_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_49.input2\[2\] sky130_fd_sc_hd__dfxtp_1
X_0927_ _0450_ _0446_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__and2b_1
X_0858_ _0246_ _0375_ _0384_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__a211o_1
X_0789_ _0117_ _0322_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__nor2_2
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0643_ CIRCUIT_1957.int_memory_1.div_1.B2 _0177_ _0181_ CIRCUIT_1957.int_memory_1.div_1.B3
+ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__a211oi_1
X_0712_ _0167_ _0250_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__nand2_1
X_0574_ net27 net16 _0108_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__mux2_1
X_1126_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result _0034_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_5.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1057_ _0141_ clknet_1_0__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__nand2_2
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_2
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_2
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0626_ _0162_ _0164_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__and2_1
X_0557_ _0115_ _0118_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__nor2_4
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1109_ CIRCUIT_1957.int_memory_1.div_1.A4 _0533_ _0519_ vssd1 vssd1 vccd1 vccd1 _0089_
+ sky130_fd_sc_hd__a21o_1
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result CIRCUIT_1957.int_memory_1.GATES_22.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result sky130_fd_sc_hd__clkbuf_16
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0609_ _0154_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 _0152_ net11 vssd1
+ vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__a31o_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ _0154_ _0156_ _0484_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__and3_1
X_0891_ _0317_ _0368_ _0429_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1111__B1 _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1102__B1 _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1090_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[3\] _0531_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0072_ sky130_fd_sc_hd__a21o_1
X_0874_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[1\] _0328_ _0333_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[1\]
+ _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__a221o_1
X_0943_ _0099_ _0378_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__nor2_1
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtholin_avalonsemi_5401_34 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_34/HI io_out[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0590_ clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__buf_1
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1211_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result _0085_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.A0 sky130_fd_sc_hd__dfxtp_1
X_1142_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result _0050_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_49.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0857_ _0386_ _0388_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or3_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0926_ _0462_ _0463_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState vssd1 vssd1
+ vccd1 vccd1 _0464_ sky130_fd_sc_hd__or3b_1
X_0788_ _0324_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__nor2_2
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1146__CLK clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0711_ _0222_ _0249_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__xnor2_1
XANTENNA__0898__A2 _0333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0642_ CIRCUIT_1957.int_memory_1.div_1.B3 _0178_ _0179_ _0180_ CIRCUIT_1957.int_memory_1.div_1.A7
+ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__o311a_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0573_ _0132_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1125_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result _0033_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_5.input2\[0\] sky130_fd_sc_hd__dfxtp_1
X_1056_ _0141_ clknet_1_0__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__nand2_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_2
X_0909_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState _0447_ vssd1 vssd1 vccd1
+ vccd1 _0448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0625_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A0 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__nor2_1
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0556_ _0116_ _0117_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__nor2_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1039_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[1\] _0524_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0046_ sky130_fd_sc_hd__a21o_1
X_1108_ _0511_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__buf_2
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1039__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0976__A _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0608_ CIRCUIT_1957.GATES_33.input2 vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__inv_2
X_0539_ CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState _0103_ CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__nor3b_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0890_ _0347_ _0369_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__or2_1
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0962__C _0149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0873_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[1\] _0331_ _0332_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__a22o_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0942_ _0456_ _0473_ _0475_ _0477_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.MEMORY_67.d
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1096__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xtholin_avalonsemi_5401_35 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_35/HI io_out[23]
+ sky130_fd_sc_hd__conb_1
XANTENNA__0793__B _0322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1210_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result _0084_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.B3 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1141_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result _0049_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_49.input2\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1087__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0856_ _0316_ _0321_ _0389_ _0394_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__a31o_1
X_0787_ CIRCUIT_1957.MEMORY_71.s_currentState CIRCUIT_1957.MEMORY_70.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__nand2b_2
X_0925_ CIRCUIT_1957.MEMORY_65.s_currentState vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
XANTENNA__1011__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0788__B _0326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0641_ CIRCUIT_1957.int_memory_1.div_1.B2 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_0710_ _0246_ _0248_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__nand2_1
XANTENNA__0979__A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__0502_ clknet_0__0502_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0502_
+ sky130_fd_sc_hd__clkbuf_16
X_0572_ CIRCUIT_1957.MEMORY_63.s_currentState CIRCUIT_1957.MEMORY_71.s_currentState
+ CIRCUIT_1957.MEMORY_87.s_currentState CIRCUIT_1957.MEMORY_79.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__mux4_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1055_ _0141_ clknet_1_1__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__nand2_2
X_1124_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result _0032_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_4.input2\[3\] sky130_fd_sc_hd__dfxtp_1
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_2
X_0908_ CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__and2b_1
X_0839_ _0115_ CIRCUIT_1957.D3 _0377_ _0119_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__a22o_2
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ CIRCUIT_1957.int_memory_1.div_1.B0 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkinv_2
XFILLER_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0555_ CIRCUIT_1957.MEMORY_68.s_currentState CIRCUIT_1957.MEMORY_69.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__nand2_2
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1107_ CIRCUIT_1957.int_memory_1.div_1.A3 _0532_ _0517_ vssd1 vssd1 vccd1 vccd1 _0088_
+ sky130_fd_sc_hd__a21o_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1038_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[0\] _0524_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0045_ sky130_fd_sc_hd__a21o_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0992__A clknet_1_0__leaf__0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0607_ CIRCUIT_1957.GATES_33.input2 _0152_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2
+ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__a21o_1
X_0538_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState _0100_ _0101_ _0102_ vssd1
+ vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__o22a_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A io_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1111__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1069__4 clknet_1_0__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__inv_2
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0941_ _0102_ _0474_ _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__a21oi_1
X_0872_ CIRCUIT_1957.int_memory_1.mul2_1.A1 CIRCUIT_1957.int_memory_1.mul2_1.B0 CIRCUIT_1957.int_memory_1.mul2_1.B1
+ CIRCUIT_1957.int_memory_1.mul2_1.A0 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__a22o_1
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtholin_avalonsemi_5401_36 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_36/HI io_out[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0984__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result CIRCUIT_1957.int_memory_1.GATES_28.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result sky130_fd_sc_hd__clkbuf_16
XFILLER_1_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1140_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result _0048_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_8.input2\[3\] sky130_fd_sc_hd__dfxtp_1
X_0924_ _0439_ _0442_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__and2_1
X_0855_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[2\] _0333_ _0334_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[2\]
+ _0393_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__a221o_1
X_0786_ _0324_ _0322_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__nor2_1
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0640_ CIRCUIT_1957.int_memory_1.div_1.A6 CIRCUIT_1957.int_memory_1.div_1.B1 CIRCUIT_1957.int_memory_1.div_1.B0
+ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__and3b_1
X_0571_ _0131_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1123_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result _0031_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_4.input2\[2\] sky130_fd_sc_hd__dfxtp_1
X_1054_ _0141_ clknet_1_1__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__nand2_2
X_0907_ _0443_ _0444_ _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__nand3_1
X_0769_ _0306_ _0307_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__nor2_1
X_0838_ _0298_ _0346_ _0376_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__or3_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0623_ CIRCUIT_1957.int_memory_1.div_1.B1 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__buf_2
X_0554_ CIRCUIT_1957.MEMORY_70.s_currentState CIRCUIT_1957.MEMORY_71.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__nand2_1
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1106_ CIRCUIT_1957.int_memory_1.div_1.A2 _0532_ _0514_ vssd1 vssd1 vccd1 vccd1 _0087_
+ sky130_fd_sc_hd__a21o_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1037_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[3\] _0524_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0044_ sky130_fd_sc_hd__a21o_1
XANTENNA__0964__A0 CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0992__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0606_ _0149_ _0151_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__nand2_1
X_0537_ CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState vssd1 vssd1 vccd1 vccd1 _0102_
+ sky130_fd_sc_hd__buf_2
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1114__B1 _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1105__B1 _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0940_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState CIRCUIT_1957.MEMORY_67.s_currentState
+ _0398_ _0459_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__a31o_1
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result
+ sky130_fd_sc_hd__clkbuf_16
X_0871_ _0304_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XANTENNA__0998__A clknet_1_0__leaf__0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0852__A2 _0331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071__6 clknet_1_1__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__inv_2
Xtholin_avalonsemi_5401_37 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_37/HI io_out[25]
+ sky130_fd_sc_hd__conb_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0854_ _0169_ _0390_ _0339_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__a31o_1
X_0923_ _0443_ _0445_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__nand2_1
X_0785_ CIRCUIT_1957.MEMORY_69.s_currentState CIRCUIT_1957.MEMORY_68.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__nand2b_2
X_1199_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result _0073_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_2.input2\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0606__A _0149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0570_ _0130_ net17 _0108_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__mux2_1
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1122_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result _0030_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_4.input2\[1\] sky130_fd_sc_hd__dfxtp_1
X_1053_ _0141_ clknet_1_1__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__nand2_2
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0837_ _0347_ _0373_ _0374_ _0375_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__a2bb2o_1
X_0906_ CIRCUIT_1957.MEMORY_65.s_currentState _0160_ vssd1 vssd1 vccd1 vccd1 _0445_
+ sky130_fd_sc_hd__nand2_1
X_0768_ CIRCUIT_1957.int_memory_1.mul2_1.B0 CIRCUIT_1957.int_memory_1.mul2_1.A3 _0303_
+ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__a21oi_1
X_0699_ _0234_ _0236_ _0222_ _0231_ _0237_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__o221ai_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0553_ CIRCUIT_1957.MEMORY_62.s_currentState _0114_ CIRCUIT_1957.MEMORY_72.s_currentState
+ CIRCUIT_1957.MEMORY_73.s_currentState vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__or4bb_4
X_0622_ CIRCUIT_1957.MEMORY_63.s_currentState _0160_ vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__and2_1
X_1105_ CIRCUIT_1957.int_memory_1.div_1.A1 _0532_ _0522_ vssd1 vssd1 vccd1 vccd1 _0086_
+ sky130_fd_sc_hd__a21o_1
X_1036_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[2\] _0524_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0043_ sky130_fd_sc_hd__a21o_1
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0605_ _0150_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__dlymetal6s2s_1
X_0536_ CIRCUIT_1957.MEMORY_66.s_currentState CIRCUIT_1957.MEMORY_65.s_currentState
+ CIRCUIT_1957.MEMORY_63.s_currentState CIRCUIT_1957.MEMORY_67.s_currentState vssd1
+ vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__or4_1
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1019_ CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__inv_2
XFILLER_43_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1041__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1032__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1099__B1 _0517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0870_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[1\] _0325_ _0342_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[1\]
+ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__a221o_1
XANTENNA__0998__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1023__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0999_ _0507_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_32.result sky130_fd_sc_hd__buf_1
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtholin_avalonsemi_5401_38 vssd1 vssd1 vccd1 vccd1 io_oeb tholin_avalonsemi_5401_38/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0853_ CIRCUIT_1957.int_memory_1.GATES_51.input2\[2\] _0341_ _0342_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[2\]
+ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a221o_1
X_0922_ _0380_ _0458_ _0460_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.MEMORY_64.d sky130_fd_sc_hd__a21oi_1
X_0784_ _0295_ _0322_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__nor2_1
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
X_1198_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result _0072_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_1.input2\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0622__A CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1121_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result _0029_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_4.input2\[0\] sky130_fd_sc_hd__dfxtp_1
X_1052_ _0141_ clknet_1_1__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__nand2_2
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0767_ CIRCUIT_1957.int_memory_1.mul2_1.B0 CIRCUIT_1957.int_memory_1.mul2_1.A3 _0303_
+ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__and3_1
X_0836_ _0116_ _0324_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__nor2_2
X_0905_ _0102_ _0439_ _0442_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__nand3_1
X_0698_ _0162_ _0233_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__or2_1
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0621_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState _0102_ CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState
+ CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__or4_2
X_0552_ CIRCUIT_1957.MEMORY_75.s_currentState CIRCUIT_1957.MEMORY_74.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__nand2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1035_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[1\] _0524_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0042_ sky130_fd_sc_hd__a21o_1
X_1104_ CIRCUIT_1957.int_memory_1.div_1.A0 _0532_ _0519_ vssd1 vssd1 vccd1 vccd1 _0085_
+ sky130_fd_sc_hd__a21o_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0819_ _0353_ _0299_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__xor2_1
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0604_ CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState
+ _0128_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__and3b_1
X_0535_ _0099_ CIRCUIT_1957.MEMORY_64.s_currentState vssd1 vssd1 vccd1 vccd1 _0100_
+ sky130_fd_sc_hd__nor2_1
XFILLER_34_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[0\] _0512_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0029_ sky130_fd_sc_hd__a21o_1
XANTENNA__1114__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0596__S _0144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A io_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0998_ clknet_1_0__leaf__0498_ _0496_ _0328_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__and3_2
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_input2_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtholin_avalonsemi_5401_39 vssd1 vssd1 vccd1 vccd1 io_out[26] tholin_avalonsemi_5401_39/LO
+ sky130_fd_sc_hd__conb_1
Xtholin_avalonsemi_5401_28 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_28/HI io_out[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0921_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
X_0852_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[2\] _0331_ _0332_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__a22o_1
X_0783_ CIRCUIT_1957.MEMORY_70.s_currentState CIRCUIT_1957.MEMORY_71.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__or2_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_1197_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result _0071_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_1.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1120_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result _0028_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_3.input2\[3\] sky130_fd_sc_hd__dfxtp_1
X_1051_ _0141_ clknet_1_1__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__nand2_2
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0904_ _0439_ _0442_ _0102_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__a21o_1
X_0766_ CIRCUIT_1957.int_memory_1.mul2_1.A1 CIRCUIT_1957.int_memory_1.mul2_1.B0 _0303_
+ _0304_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__a31o_1
X_0835_ _0215_ _0219_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__nand2_1
X_0697_ CIRCUIT_1957.int_memory_1.div_1.A3 _0235_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__xnor2_2
XANTENNA__0900__B1 _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0551_ CIRCUIT_1957.MEMORY_73.s_currentState CIRCUIT_1957.MEMORY_81.s_currentState
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__mux2_1
X_0620_ _0151_ _0159_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_53.result sky130_fd_sc_hd__nor2_1
XFILLER_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1103_ CIRCUIT_1957.int_memory_1.mul2_1.B3 _0532_ _0517_ vssd1 vssd1 vccd1 vccd1
+ _0084_ sky130_fd_sc_hd__a21o_1
X_1034_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[0\] _0524_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0041_ sky130_fd_sc_hd__a21o_1
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0818_ _0356_ _0348_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__or2b_1
X_0749_ _0168_ _0281_ _0282_ _0287_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__a31o_1
XFILLER_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0603_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState CIRCUIT_1957.clock_gen_2_1.GATES_1.input2
+ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__nand2_2
X_0534_ CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState vssd1 vssd1 vccd1 vccd1 _0099_
+ sky130_fd_sc_hd__clkinv_2
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1017_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__0873__A2 _0331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0855__A2 _0333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1032__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result CIRCUIT_1957.int_memory_1.GATES_23.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result sky130_fd_sc_hd__clkbuf_16
X_0997_ _0506_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_31.result sky130_fd_sc_hd__buf_1
Xtholin_avalonsemi_5401_29 vssd1 vssd1 vccd1 vccd1 tholin_avalonsemi_5401_29/HI io_out[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0920_ _0126_ _0160_ _0128_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__a21o_2
X_0851_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A6 _0174_ vssd1 vssd1 vccd1 vccd1 _0390_
+ sky130_fd_sc_hd__o21a_1
X_0782_ _0319_ _0320_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__nor2_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1196_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result _0070_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_1.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1050_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState vssd1 vssd1 vccd1 vccd1
+ _0003_ sky130_fd_sc_hd__clkinv_2
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0834_ _0355_ _0372_ _0354_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0903_ _0440_ _0115_ _0402_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__o31a_1
X_0765_ CIRCUIT_1957.int_memory_1.mul2_1.A0 CIRCUIT_1957.int_memory_1.mul2_1.A1 CIRCUIT_1957.int_memory_1.mul2_1.B0
+ CIRCUIT_1957.int_memory_1.mul2_1.B1 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__and4_1
X_0696_ _0215_ _0219_ _0163_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1179_ net40 _0053_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0550_ net19 _0108_ _0112_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__a21o_1
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1102_ CIRCUIT_1957.int_memory_1.mul2_1.B2 _0532_ _0514_ vssd1 vssd1 vccd1 vccd1
+ _0083_ sky130_fd_sc_hd__a21o_1
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1033_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[3\] _0524_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0040_ sky130_fd_sc_hd__a21o_1
X_0817_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nor2_1
X_0679_ _0168_ _0216_ _0217_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__mux2_1
X_0748_ _0283_ _0284_ _0286_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1080__A_N net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0602_ CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 sky130_fd_sc_hd__inv_2
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1016_ _0463_ _0511_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__nor2_2
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1044__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1035__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1026__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0996_ clknet_1_0__leaf__0498_ _0496_ _0332_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__and3_2
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0850_ _0300_ _0313_ _0315_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__nand3_1
X_0781_ CIRCUIT_1957.MEMORY_68.s_currentState CIRCUIT_1957.MEMORY_69.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__nand2b_2
Xinput4 io_in[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1195_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result _0069_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_1.input2\[0\] sky130_fd_sc_hd__dfxtp_1
X_0979_ clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__buf_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ _0351_ _0357_ _0361_ _0371_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__a31o_1
XFILLER_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0902_ _0115_ CIRCUIT_1957.D0 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__nand2_1
X_0764_ CIRCUIT_1957.int_memory_1.mul2_1.A2 CIRCUIT_1957.int_memory_1.mul2_1.B1 vssd1
+ vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__and2_1
X_0695_ _0162_ _0233_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__and2_1
X_1178_ CIRCUIT_1957.GATES_60.result CIRCUIT_1957.MEMORY_62.d _0018_ vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_62.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1101_ CIRCUIT_1957.int_memory_1.mul2_1.B1 _0532_ _0522_ vssd1 vssd1 vccd1 vccd1
+ _0082_ sky130_fd_sc_hd__a21o_1
X_1032_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[2\] _0524_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0039_ sky130_fd_sc_hd__a21o_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0816_ _0351_ _0352_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__a21oi_1
X_0747_ _0168_ _0285_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__xnor2_1
X_0678_ _0189_ _0197_ _0184_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__or3b_1
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1117__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0601_ _0148_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.D3 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1015_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[3\] _0512_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0028_ sky130_fd_sc_hd__a21o_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0995_ _0505_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_30.result sky130_fd_sc_hd__buf_1
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0780_ CIRCUIT_1957.MEMORY_70.s_currentState CIRCUIT_1957.MEMORY_71.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__nand2b_1
XFILLER_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 io_in[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1194_ clknet_1_1__leaf_clk _0068_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dfxtp_1
XANTENNA__1004__A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0978_ _0497_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_21.result sky130_fd_sc_hd__buf_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__0143_ clknet_0__0143_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0143_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0901_ net9 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
X_0832_ _0363_ _0370_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__and2_1
X_0763_ _0299_ _0300_ _0301_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__o21ba_1
X_0694_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A2 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__nor2_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1177_ CIRCUIT_1957.GATES_9.result CIRCUIT_1957.MEMORY_63.d vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.MEMORY_63.s_currentState sky130_fd_sc_hd__dfxtp_2
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1100_ CIRCUIT_1957.int_memory_1.mul2_1.B0 _0532_ _0519_ vssd1 vssd1 vccd1 vccd1
+ _0081_ sky130_fd_sc_hd__a21o_1
X_1031_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[1\] _0524_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0038_ sky130_fd_sc_hd__a21o_1
X_0815_ _0353_ _0351_ _0352_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__a21oi_1
X_0746_ _0254_ _0260_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__nand2_1
X_0677_ _0168_ _0184_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__nand2_1
XFILLER_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result CIRCUIT_1957.int_memory_1.GATES_29.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result sky130_fd_sc_hd__clkbuf_16
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0600_ net8 net4 _0144_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__mux2_1
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1014_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__1012__A CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0729_ _0166_ CIRCUIT_1957.int_memory_1.div_1.A1 _0267_ vssd1 vssd1 vccd1 vccd1 _0268_
+ sky130_fd_sc_hd__and3_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1035__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1007__A _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0994_ clknet_1_0__leaf__0498_ _0496_ _0325_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__and3_2
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 io_in[5] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1004__B _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1193_ clknet_1_1__leaf_clk _0067_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__dfxtp_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0977_ clknet_1_1__leaf__0142_ _0496_ _0327_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and3_2
XFILLER_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1092__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f__0142_ clknet_0__0142_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0142_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0900_ _0428_ _0430_ _0438_ _0119_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__o31ai_2
X_0831_ _0366_ _0367_ _0369_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__o21bai_1
X_0762_ CIRCUIT_1957.int_memory_1.mul2_1.B3 CIRCUIT_1957.int_memory_1.mul2_1.A0 CIRCUIT_1957.int_memory_1.mul2_1.B2
+ CIRCUIT_1957.int_memory_1.mul2_1.A1 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__a22oi_1
X_0693_ _0231_ _0222_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__nand2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result
+ sky130_fd_sc_hd__clkbuf_16
X_1176_ CIRCUIT_1957.GATES_10.result CIRCUIT_1957.MEMORY_64.d _0017_ vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_64.s_currentState sky130_fd_sc_hd__dfrtp_1
XANTENNA__1074__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1030_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[0\] _0524_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0037_ sky130_fd_sc_hd__a21o_1
X_0814_ CIRCUIT_1957.int_memory_1.mul2_1.B2 CIRCUIT_1957.int_memory_1.mul2_1.A2 vssd1
+ vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result
+ sky130_fd_sc_hd__clkbuf_16
X_0676_ _0167_ _0205_ _0209_ _0213_ _0214_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__a221o_1
X_0745_ _0283_ _0265_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__nor2_1
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1159_ CIRCUIT_1957.GATES_40.result CIRCUIT_1957.GATES_28.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_81.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1038__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1013_ _0516_ _0511_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__nor2_2
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0659_ _0167_ _0177_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__nand2_1
X_0728_ _0251_ _0254_ _0260_ _0266_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__a31o_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1108__A _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0993_ _0504_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_29.result sky130_fd_sc_hd__buf_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 io_in[6] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_1192_ clknet_1_1__leaf_clk _0066_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dfxtp_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0976_ _0119_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__buf_2
XANTENNA__1020__B _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _0317_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__nor2_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0761_ CIRCUIT_1957.int_memory_1.mul2_1.A0 CIRCUIT_1957.int_memory_1.mul2_1.B2 vssd1
+ vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__nand2_1
X_0692_ CIRCUIT_1957.int_memory_1.div_1.B2 vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1175_ CIRCUIT_1957.GATES_9.result CIRCUIT_1957.MEMORY_65.d vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.MEMORY_65.s_currentState sky130_fd_sc_hd__dfxtp_1
X_0959_ _0487_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_40.result sky130_fd_sc_hd__clkbuf_1
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0576__A0 CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 io_in[9] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_0813_ CIRCUIT_1957.int_memory_1.mul2_1.B3 CIRCUIT_1957.int_memory_1.mul2_1.A3 vssd1
+ vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__nand2_1
X_0675_ _0211_ _0212_ CIRCUIT_1957.int_memory_1.div_1.B2 vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__o21a_1
X_0744_ _0250_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
X_1158_ CIRCUIT_1957.GATES_40.result CIRCUIT_1957.GATES_30.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_82.s_currentState sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__0143_ _0143_ vssd1 vssd1 vccd1 vccd1 clknet_0__0143_ sky130_fd_sc_hd__clkbuf_16
X_1089_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[2\] _0531_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0071_ sky130_fd_sc_hd__a21o_1
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1012_ CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__inv_2
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0727_ _0167_ _0250_ _0265_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0658_ CIRCUIT_1957.int_memory_1.div_1.B2 _0188_ _0191_ _0196_ vssd1 vssd1 vccd1
+ vccd1 _0197_ sky130_fd_sc_hd__o2bb2a_1
X_0589_ _0140_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__buf_4
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1110__B1 _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1101__B1 _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0992_ clknet_1_0__leaf__0498_ _0496_ _0323_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__and3_2
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 io_in[7] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_1191_ clknet_1_1__leaf_clk _0065_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dfxtp_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0975_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState
+ _0460_ CIRCUIT_1957.GATES_10.result vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_9.result
+ sky130_fd_sc_hd__a31o_1
XANTENNA__1029__A _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0760_ CIRCUIT_1957.int_memory_1.mul2_1.B3 CIRCUIT_1957.int_memory_1.mul2_1.A1 vssd1
+ vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__nand2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0691_ _0167_ _0229_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__nand2_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1174_ CIRCUIT_1957.GATES_9.result CIRCUIT_1957.MEMORY_66.d vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.MEMORY_66.s_currentState sky130_fd_sc_hd__dfxtp_2
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0889_ _0426_ _0427_ _0296_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a21oi_1
X_0958_ CIRCUIT_1957.GATES_33.input2 _0484_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__and2_1
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1067__2 clknet_1_0__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__inv_2
XFILLER_46_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 rst vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
X_0812_ _0348_ _0349_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__or3_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0743_ _0279_ _0280_ _0278_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__a21o_1
X_0674_ CIRCUIT_1957.int_memory_1.div_1.B2 _0211_ _0212_ vssd1 vssd1 vccd1 vccd1 _0213_
+ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1157_ CIRCUIT_1957.GATES_40.result CIRCUIT_1957.GATES_35.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_83.s_currentState sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__0142_ _0142_ vssd1 vssd1 vccd1 vccd1 clknet_0__0142_ sky130_fd_sc_hd__clkbuf_16
X_1088_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[1\] _0531_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0070_ sky130_fd_sc_hd__a21o_1
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1038__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[2\] _0512_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0027_ sky130_fd_sc_hd__a21o_1
XFILLER_19_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0726_ _0229_ _0261_ _0264_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__mux2_1
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0657_ _0193_ _0194_ _0195_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__o21ba_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0588_ net11 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1209_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result _0083_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.B2 sky130_fd_sc_hd__dfxtp_1
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0709_ _0231_ _0247_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input9_A io_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0991_ _0338_ clknet_1_1__leaf__0502_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_28.result
+ sky130_fd_sc_hd__nor2_2
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1095__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 io_in[8] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_1190_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result _0064_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_51.input2\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ _0495_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_10.result sky130_fd_sc_hd__clkbuf_1
XFILLER_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1077__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0690_ _0223_ _0228_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1173_ CIRCUIT_1957.GATES_9.result CIRCUIT_1957.MEMORY_67.d vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.MEMORY_67.s_currentState sky130_fd_sc_hd__dfxtp_2
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0888_ _0166_ _0292_ CIRCUIT_1957.int_memory_1.div_1.A0 vssd1 vssd1 vccd1 vccd1 _0427_
+ sky130_fd_sc_hd__a21bo_1
X_0957_ _0486_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_41.result sky130_fd_sc_hd__clkbuf_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result CIRCUIT_1957.int_memory_1.GATES_24.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result sky130_fd_sc_hd__clkbuf_16
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0811_ CIRCUIT_1957.int_memory_1.mul2_1.B3 CIRCUIT_1957.int_memory_1.mul2_1.B2 CIRCUIT_1957.int_memory_1.mul2_1.A3
+ CIRCUIT_1957.int_memory_1.mul2_1.A2 vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__and4_1
X_0673_ _0210_ _0191_ _0195_ _0201_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__nor4_1
X_0742_ _0278_ _0279_ _0280_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__nand3_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1087_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[0\] _0531_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0069_ sky130_fd_sc_hd__a21o_1
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1156_ CIRCUIT_1957.GATES_42.result CIRCUIT_1957.GATES_27.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_84.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0797__A2 _0331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1010_ _0514_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0656_ CIRCUIT_1957.int_memory_1.div_1.B1 _0190_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__and2_1
X_0725_ _0262_ _0263_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__nor2_1
XFILLER_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1208_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result _0082_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.B1 sky130_fd_sc_hd__dfxtp_1
X_0587_ _0139_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1139_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result _0047_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_8.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0786__B _0322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0639_ CIRCUIT_1957.int_memory_1.div_1.B0 CIRCUIT_1957.int_memory_1.div_1.B1 vssd1
+ vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__nor2_1
X_0708_ _0234_ _0236_ _0237_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__o21ai_1
XANTENNA__0933__A2 CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1110__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0990_ _0503_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_27.result sky130_fd_sc_hd__buf_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState
+ _0447_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__and3_1
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0794__B _0326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1172_ CIRCUIT_1957.GATES_38.result CIRCUIT_1957.GATES_27.result _0016_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_68.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0956_ _0128_ _0127_ _0149_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__and3_1
X_0887_ _0164_ _0292_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__nand2_1
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0789__B _0322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0810_ CIRCUIT_1957.int_memory_1.mul2_1.B2 CIRCUIT_1957.int_memory_1.mul2_1.A3 CIRCUIT_1957.int_memory_1.mul2_1.A2
+ CIRCUIT_1957.int_memory_1.mul2_1.B3 vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__a22oi_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0672_ _0191_ _0195_ _0201_ _0210_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__o31a_1
X_0741_ _0231_ _0253_ _0267_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__nand3_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1224_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result _0098_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_3.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1155_ CIRCUIT_1957.GATES_42.result CIRCUIT_1957.GATES_28.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_85.s_currentState sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result CIRCUIT_1957.int_memory_1.GATES_30.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result sky130_fd_sc_hd__clkbuf_16
X_1086_ _0511_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__buf_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0939_ _0102_ _0474_ _0454_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0982__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0655_ _0166_ _0187_ _0192_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__a21oi_1
X_0724_ _0232_ _0238_ _0168_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__a21oi_1
X_0586_ net12 net13 _0108_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__mux2_1
X_1207_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result _0081_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.B0 sky130_fd_sc_hd__dfxtp_1
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1138_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result _0046_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_8.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0977__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ _0230_ _0232_ _0238_ _0245_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__a31o_2
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0638_ CIRCUIT_1957.int_memory_1.div_1.A7 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
X_0569_ _0125_ _0129_ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState vssd1 vssd1
+ vccd1 vccd1 _0130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__0498_ clknet_0__0498_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0498_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0972_ _0494_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_27.result sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1171_ CIRCUIT_1957.GATES_38.result CIRCUIT_1957.GATES_28.result _0015_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_69.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0955_ _0485_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_42.result sky130_fd_sc_hd__clkbuf_1
X_0886_ _0423_ _0424_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result CIRCUIT_1957.int_memory_1.GATES_53.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result sky130_fd_sc_hd__clkbuf_16
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0740_ _0231_ _0267_ _0253_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__a21o_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0671_ _0193_ _0194_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__nor2_1
XANTENNA__0996__A clknet_1_0__leaf__0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1154_ CIRCUIT_1957.GATES_42.result CIRCUIT_1957.GATES_30.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_86.s_currentState sky130_fd_sc_hd__dfxtp_1
X_1223_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result _0097_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_3.input2\[0\] sky130_fd_sc_hd__dfxtp_1
X_1085_ _0530_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
X_0938_ _0398_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__inv_2
X_0869_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[1\] _0323_ _0334_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__a22o_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0982__C _0333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0723_ _0168_ _0232_ _0238_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__and3_1
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0654_ _0166_ _0192_ _0187_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__and3_1
X_0585_ _0138_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_1206_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result _0080_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.A3 sky130_fd_sc_hd__dfxtp_1
X_1137_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result _0045_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_8.input2\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0881__B1 _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0706_ _0167_ _0229_ _0244_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__o21bai_1
X_0637_ CIRCUIT_1957.int_memory_1.div_1.B1 _0175_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__nand2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0568_ _0120_ _0127_ _0128_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__o21a_1
XANTENNA__1031__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1098__B1 _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1022__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1089__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A io_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ CIRCUIT_1957.MEMORY_65.s_currentState _0493_ CIRCUIT_1957.MEMORY_62.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__mux2_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0612__A _0149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1170_ CIRCUIT_1957.GATES_38.result CIRCUIT_1957.GATES_30.result _0014_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_70.s_currentState sky130_fd_sc_hd__dfrtp_1
X_0954_ _0154_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 _0484_ vssd1 vssd1
+ vccd1 vccd1 _0485_ sky130_fd_sc_hd__and3_1
X_0885_ CIRCUIT_1957.MEMORY_66.s_currentState _0160_ vssd1 vssd1 vccd1 vccd1 _0424_
+ sky130_fd_sc_hd__and2_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0670_ _0207_ _0200_ _0208_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0996__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1222_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result _0096_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.B3 sky130_fd_sc_hd__dfxtp_1
X_1153_ CIRCUIT_1957.GATES_42.result CIRCUIT_1957.GATES_35.result vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_87.s_currentState sky130_fd_sc_hd__dfxtp_1
X_1084_ net11 net24 vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__and2b_1
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0799_ _0116_ _0320_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__or2_1
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0937_ _0425_ _0453_ _0455_ _0460_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__a31o_1
X_0868_ _0405_ _0406_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__and2b_1
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0653_ CIRCUIT_1957.int_memory_1.div_1.A5 vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
X_0722_ _0229_ _0244_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__nand2_1
XANTENNA__0945__A2 CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0584_ CIRCUIT_1957.MEMORY_65.s_currentState CIRCUIT_1957.MEMORY_68.s_currentState
+ CIRCUIT_1957.MEMORY_84.s_currentState CIRCUIT_1957.MEMORY_76.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__mux4_1
X_1205_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result _0079_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.A2 sky130_fd_sc_hd__dfxtp_1
X_1136_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result _0044_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_7.input2\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1113__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0636_ CIRCUIT_1957.int_memory_1.div_1.B0 _0169_ _0174_ _0170_ vssd1 vssd1 vccd1
+ vccd1 _0175_ sky130_fd_sc_hd__a31o_1
X_0705_ _0239_ _0240_ _0243_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__mux2_1
X_0567_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState _0102_ vssd1 vssd1 vccd1
+ vccd1 _0128_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result
+ sky130_fd_sc_hd__clkbuf_16
X_1119_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result _0027_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_3.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0619_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__nand2_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0970_ _0462_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__inv_2
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1086__A _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__0498_ _0498_ vssd1 vssd1 vccd1 vccd1 clknet_0__0498_ sky130_fd_sc_hd__clkbuf_16
X_1072__7 clknet_1_1__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__inv_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0803__A _0295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0953_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState
+ _0151_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__and3_1
X_0884_ _0102_ _0422_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__xnor2_1
XANTENNA__0966__A0 CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0594__S _0144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1221_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result _0095_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.B2 sky130_fd_sc_hd__dfxtp_2
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1083_ _0529_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
X_1152_ clknet_1_1__leaf_clk CIRCUIT_1957.GATES_53.result _0008_ vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_1957.MEMORY_88.s_currentState sky130_fd_sc_hd__dfrtp_1
X_0936_ _0453_ _0459_ _0468_ _0471_ _0472_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.MEMORY_66.d
+ sky130_fd_sc_hd__a32o_1
X_0798_ _0162_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_0867_ _0403_ _0270_ _0292_ _0404_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__a31o_1
XFILLER_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1116__B1 _0517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0652_ CIRCUIT_1957.int_memory_1.div_1.B1 _0190_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__nor2_1
X_0721_ _0256_ _0258_ _0253_ _0231_ _0259_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__o221ai_2
X_0583_ _0137_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1204_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result _0078_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1107__B1 _0517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1135_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result _0043_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_7.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1078__B net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0919_ _0400_ _0456_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0635_ CIRCUIT_1957.int_memory_1.div_1.A7 CIRCUIT_1957.int_memory_1.div_1.B1 vssd1
+ vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__or2b_1
X_0704_ _0168_ _0242_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__xnor2_1
X_0566_ _0126_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result
+ sky130_fd_sc_hd__clkbuf_16
X_1049_ _0141_ clknet_1_1__leaf__0526_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__nand2_2
X_1118_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[1\] _0533_ _0522_ vssd1 vssd1 vccd1
+ vccd1 _0098_ sky130_fd_sc_hd__a21o_1
XANTENNA__1031__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__0143_ clknet_0__0143_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0143_
+ sky130_fd_sc_hd__clkbuf_16
X_0549_ _0110_ _0111_ _0108_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__a21oi_1
X_0618_ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d sky130_fd_sc_hd__clkinv_2
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0536__A CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ _0151_ _0159_ CIRCUIT_1957.MEMORY_88.s_currentState vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.GATES_60.result sky130_fd_sc_hd__o21a_1
X_0883_ _0401_ _0115_ _0402_ _0420_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__o311a_1
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1097__A _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1220_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result _0094_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.div_1.B1 sky130_fd_sc_hd__dfxtp_2
X_1151_ CIRCUIT_1957.clock_gen_2_1.CLK1 CIRCUIT_1957.D3 _0007_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__0893__B1 _0331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1082_ net11 net22 vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and2b_1
X_0866_ _0403_ _0270_ _0404_ _0292_ _0296_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__a41o_1
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0935_ _0099_ _0469_ _0424_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__a21o_1
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0797_ CIRCUIT_1957.int_memory_1.GATES_7.input2\[3\] _0331_ _0332_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[3\]
+ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__a221o_1
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0720_ _0162_ _0255_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__or2_1
XFILLER_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0651_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A4 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__nor2_1
X_0582_ net23 net14 _0108_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__mux2_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1203_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result _0077_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.mul2_1.A0 sky130_fd_sc_hd__dfxtp_1
X_1134_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result _0042_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_7.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1065_ _0140_ clknet_1_0__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__nand2_2
XANTENNA__1043__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0918_ _0161_ _0379_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__xor2_1
X_0849_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[2\] _0328_ _0325_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[2\]
+ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__a221o_1
XANTENNA__0609__B1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1034__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0703_ _0223_ _0241_ _0226_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1025__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0634_ _0171_ _0172_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__nand2_1
X_0565_ CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__nand2_1
X_1117_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[0\] _0533_ _0519_ vssd1 vssd1 vccd1
+ vccd1 _0097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1048_ clknet_1_1__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__buf_1
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__0142_ clknet_0__0142_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0142_
+ sky130_fd_sc_hd__clkbuf_16
X_0548_ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState CIRCUIT_1957.MEMORY_82.s_currentState
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__o21ai_1
X_0617_ _0154_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result _0149_ _0151_ _0155_
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result sky130_fd_sc_hd__a41o_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input5_A io_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0951_ _0483_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.MEMORY_62.d sky130_fd_sc_hd__clkbuf_1
X_0882_ _0115_ CIRCUIT_1957.D1 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result
+ sky130_fd_sc_hd__clkbuf_16
X_1150_ CIRCUIT_1957.clock_gen_2_1.CLK1 CIRCUIT_1957.D2 _0006_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1081_ _0528_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0934_ _0102_ _0422_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__a21oi_1
X_0865_ _0268_ _0269_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__nor2_1
X_0796_ CIRCUIT_1957.int_memory_1.GATES_2.input2\[3\] _0333_ _0334_ CIRCUIT_1957.int_memory_1.GATES_1.input2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__a22o_1
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1116__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0572__A0 CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0915__A CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0650_ CIRCUIT_1957.int_memory_1.div_1.B2 _0188_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__nor2_1
X_0581_ _0136_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1133_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result _0041_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_7.input2\[0\] sky130_fd_sc_hd__dfxtp_1
X_1202_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result _0076_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_2.input2\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1064_ _0140_ clknet_1_0__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__nand2_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0779_ _0312_ _0316_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__nand2_1
XANTENNA__0560__A _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0917_ _0425_ _0453_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__a21oi_1
X_0848_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[2\] _0327_ _0323_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__a22o_1
XFILLER_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result CIRCUIT_1957.int_memory_1.GATES_25.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result sky130_fd_sc_hd__clkbuf_16
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0633_ _0163_ CIRCUIT_1957.int_memory_1.div_1.A5 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__nor2_1
X_0702_ _0207_ _0200_ _0208_ _0180_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__a211o_1
X_0564_ CIRCUIT_1957.MEMORY_72.s_currentState CIRCUIT_1957.MEMORY_80.s_currentState
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__mux2_1
X_1116_ _0167_ _0533_ _0517_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__a21o_1
X_1047_ _0141_ clknet_1_1__leaf__0143_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__nand2_2
XANTENNA__0839__B2 _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0616_ _0158_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_33.input2 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0547_ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState _0104_ CIRCUIT_1957.MEMORY_74.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__or3b_1
XFILLER_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0536__C CIRCUIT_1957.MEMORY_63.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0950_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState _0099_ _0120_ vssd1 vssd1
+ vccd1 vccd1 _0483_ sky130_fd_sc_hd__and3_1
X_0881_ _0407_ _0419_ _0119_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1080_ net11 net21 vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and2b_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0933_ CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState CIRCUIT_1957.MEMORY_66.s_currentState
+ _0469_ _0459_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__a31o_1
X_0795_ _0320_ _0326_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__nor2_2
X_0864_ _0165_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1201_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result _0075_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_2.input2\[2\] sky130_fd_sc_hd__dfxtp_1
X_0580_ CIRCUIT_1957.MEMORY_66.s_currentState CIRCUIT_1957.MEMORY_69.s_currentState
+ CIRCUIT_1957.MEMORY_85.s_currentState CIRCUIT_1957.MEMORY_77.s_currentState CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__mux4_1
X_1132_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result _0040_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_6.input2\[3\] sky130_fd_sc_hd__dfxtp_1
X_1063_ _0140_ clknet_1_1__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__nand2_2
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0916_ _0399_ _0454_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__xor2_1
X_0778_ _0312_ _0316_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__or2_1
X_0847_ _0347_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__nor2_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1034__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0632_ _0166_ _0169_ _0170_ CIRCUIT_1957.int_memory_1.div_1.B1 vssd1 vssd1 vccd1
+ vccd1 _0171_ sky130_fd_sc_hd__a211o_1
X_0701_ _0239_ _0218_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__nor2_1
X_0563_ _0124_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__0600__S _0144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1115_ _0231_ _0533_ _0514_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1046_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[3\] _0525_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0052_ sky130_fd_sc_hd__a21o_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result CIRCUIT_1957.int_memory_1.GATES_31.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result sky130_fd_sc_hd__clkbuf_16
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0546_ _0109_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0615_ _0140_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 _0157_ vssd1 vssd1
+ vccd1 vccd1 _0158_ sky130_fd_sc_hd__and3b_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1029_ _0511_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__buf_2
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0536__D CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1010__A _0514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1091__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1082__A_N net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0880_ _0267_ _0375_ _0418_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__a21o_1
XFILLER_11_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0932_ _0422_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__inv_2
X_0794_ _0117_ _0326_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__nor2_2
X_0863_ _0118_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1046__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1037__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1200_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result _0074_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_2.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1062_ _0140_ clknet_1_0__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__nand2_2
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1131_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result _0039_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_6.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1028__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1002__B _0119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0915_ CIRCUIT_1957.MEMORY_67.s_currentState _0160_ vssd1 vssd1 vccd1 vccd1 _0454_
+ sky130_fd_sc_hd__nand2_1
X_0846_ _0355_ _0372_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__xnor2_1
X_0777_ _0313_ _0315_ _0300_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__a21o_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0700_ _0205_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
X_0631_ CIRCUIT_1957.int_memory_1.div_1.A6 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
X_0562_ _0123_ net18 _0108_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__mux2_1
X_1114_ _0162_ _0533_ _0522_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__a21o_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1045_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[2\] _0525_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0051_ sky130_fd_sc_hd__a21o_1
X_0829_ _0366_ _0367_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1008__A CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0545_ _0106_ net20 _0108_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__mux2_1
X_0614_ _0156_ CIRCUIT_1957.GATES_33.input2 _0152_ vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__mux2_1
X_1028_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[3\] _0512_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0036_ sky130_fd_sc_hd__a21o_1
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input11_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__0526_ clknet_0__0526_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__0526_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1021__A _0522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_A io_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0862_ net10 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
X_0931_ _0451_ _0452_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__or2_1
X_0793_ _0320_ _0322_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__nor2_2
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0590__A clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1130_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result _0038_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_6.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061_ _0140_ clknet_1_0__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__nand2_2
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0845_ _0382_ _0383_ _0296_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__o21ba_1
X_0914_ _0451_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__nand2_1
X_0776_ _0305_ _0314_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__or2_1
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0630_ CIRCUIT_1957.int_memory_1.div_1.B3 CIRCUIT_1957.int_memory_1.div_1.B2 vssd1
+ vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__nor2_2
X_0561_ _0113_ _0122_ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState vssd1 vssd1
+ vccd1 vccd1 _0123_ sky130_fd_sc_hd__mux2_1
X_1113_ _0166_ _0533_ _0519_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__a21o_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1044_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[1\] _0525_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1013__B _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0828_ _0299_ _0300_ _0301_ _0311_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__o22a_1
X_0759_ _0289_ _0294_ _0297_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__o21a_1
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0613_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 vssd1 vssd1 vccd1 vccd1 _0156_
+ sky130_fd_sc_hd__inv_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0544_ _0107_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__buf_2
X_1027_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[2\] _0512_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0035_ sky130_fd_sc_hd__a21o_1
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0757__B _0295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1019__A CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0588__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0792_ _0295_ _0326_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__nor2_2
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0861_ CIRCUIT_1957.MEMORY_67.s_currentState _0160_ _0399_ vssd1 vssd1 vccd1 vccd1
+ _0400_ sky130_fd_sc_hd__and3_1
X_0930_ _0444_ _0460_ _0461_ _0464_ _0467_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.MEMORY_65.d
+ sky130_fd_sc_hd__a41o_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1016__B _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1037__A2 _0524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1060_ _0140_ clknet_1_0__leaf__0142_ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__nand2_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0775_ CIRCUIT_1957.int_memory_1.mul2_1.B0 CIRCUIT_1957.int_memory_1.mul2_1.A2 CIRCUIT_1957.int_memory_1.mul2_1.B1
+ CIRCUIT_1957.int_memory_1.mul2_1.A1 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__a22oi_1
X_0844_ _0273_ _0274_ _0292_ _0381_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__a22oi_1
Xclkbuf_1_0__f__0498_ clknet_0__0498_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__0498_
+ sky130_fd_sc_hd__clkbuf_16
X_0913_ _0423_ _0424_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__xor2_1
X_1189_ clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result _0063_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_51.input2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0560_ _0119_ _0121_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__nor2_1
X_1112_ CIRCUIT_1957.int_memory_1.div_1.A7 _0533_ _0517_ vssd1 vssd1 vccd1 vccd1 _0092_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1043_ CIRCUIT_1957.int_memory_1.GATES_49.input2\[0\] _0525_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0049_ sky130_fd_sc_hd__a21o_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0827_ _0364_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__or2_1
X_0758_ _0289_ _0294_ _0296_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__a21oi_1
X_0689_ _0215_ _0219_ _0226_ _0227_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__a211oi_1
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0612_ _0149_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.clock_gen_2_1.CLK1 sky130_fd_sc_hd__inv_2
X_0543_ net22 net21 net25 net24 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__or4b_1
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1026_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[1\] _0512_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0034_ sky130_fd_sc_hd__a21o_1
XANTENNA__1040__A _0511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1094__B1 _0518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1076__B1 _0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _0513_ _0511_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nor2_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0784__A _0295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result
+ sky130_fd_sc_hd__clkbuf_16
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0860_ _0099_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__xnor2_1
X_0791_ CIRCUIT_1957.int_memory_1.GATES_3.input2\[3\] _0323_ _0325_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[3\]
+ _0329_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__a221o_1
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0989_ clknet_1_1__leaf__0498_ _0496_ _0375_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__and3_2
Xclkbuf_0__0526_ _0526_ vssd1 vssd1 vccd1 vccd1 clknet_0__0526_ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0796__A2 _0333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0912_ _0446_ _0449_ _0450_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__a21o_1
X_0774_ _0303_ _0304_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__nand2_1
X_0843_ _0273_ _0274_ _0292_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__and4_1
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1188_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result _0062_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_51.input2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0792__A _0295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1111_ CIRCUIT_1957.int_memory_1.div_1.A6 _0533_ _0514_ vssd1 vssd1 vccd1 vccd1 _0091_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[3\] _0525_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0048_ sky130_fd_sc_hd__a21o_1
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0826_ _0358_ _0360_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__nor2_1
X_0688_ CIRCUIT_1957.int_memory_1.div_1.B2 _0209_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__and2_1
X_0757_ _0116_ _0295_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__or2_2
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0542_ CIRCUIT_1957.MEMORY_62.s_currentState _0105_ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d
+ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__mux2_1
X_0611_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1
+ sky130_fd_sc_hd__inv_2
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1025_ CIRCUIT_1957.int_memory_1.GATES_5.input2\[0\] _0512_ _0520_ vssd1 vssd1 vccd1
+ vccd1 _0033_ sky130_fd_sc_hd__a21o_1
X_0809_ CIRCUIT_1957.int_memory_1.mul2_1.A3 _0305_ _0306_ vssd1 vssd1 vccd1 vccd1
+ _0348_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0980__A clknet_1_0__leaf__0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result
+ sky130_fd_sc_hd__clkbuf_16
X_1008_ CIRCUIT_1957.MEMORY_67.s_currentState vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__inv_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0784__B _0322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0885__A CIRCUIT_1957.MEMORY_66.s_currentState vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0790_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[3\] _0327_ _0328_ CIRCUIT_1957.int_memory_1.GATES_6.input2\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__a22o_1
X_0988_ _0296_ clknet_1_0__leaf__0502_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_26.result
+ sky130_fd_sc_hd__nor2_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1068__3 clknet_1_0__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__inv_2
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0956__C _0149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0842_ _0180_ _0271_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__xnor2_1
X_0911_ _0443_ _0444_ _0445_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__a21oi_1
X_0773_ _0302_ _0311_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__xor2_1
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1187_ clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result _0061_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_51.input2\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__1112__B1 _0517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0792__B _0326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ CIRCUIT_1957.int_memory_1.div_1.A5 _0533_ _0522_ vssd1 vssd1 vccd1 vccd1 _0090_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__1103__B1 _0517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ CIRCUIT_1957.int_memory_1.GATES_8.input2\[2\] _0525_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0047_ sky130_fd_sc_hd__a21o_1
XFILLER_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0825_ _0358_ _0360_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__and2_1
XFILLER_9_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0687_ _0224_ _0208_ _0225_ _0207_ _0180_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__o311a_1
X_0756_ CIRCUIT_1957.MEMORY_68.s_currentState CIRCUIT_1957.MEMORY_69.s_currentState
+ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__or2_1
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0541_ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d sky130_fd_sc_hd__clkinv_2
X_0610_ CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 _0153_ _0155_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 sky130_fd_sc_hd__a21o_1
X_1024_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[3\] _0512_ _0518_ vssd1 vssd1 vccd1
+ vccd1 _0032_ sky130_fd_sc_hd__a21o_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0808_ _0117_ _0319_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__or2_1
X_0739_ _0256_ _0258_ _0259_ _0267_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__o211ai_1
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0980__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__buf_2
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result CIRCUIT_1957.int_memory_1.GATES_26.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result sky130_fd_sc_hd__clkbuf_16
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0795__B _0326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0987_ _0347_ clknet_1_0__leaf__0502_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_25.result
+ sky130_fd_sc_hd__nor2_2
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0772_ _0309_ _0310_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__or2_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0841_ _0161_ _0379_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__nand2_1
X_0910_ CIRCUIT_1957.MEMORY_64.s_currentState _0102_ _0448_ vssd1 vssd1 vccd1 vccd1
+ _0449_ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1186_ net47 _0060_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__dfxtp_1
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1070__5 clknet_1_0__leaf__0143_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__inv_2
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1040_ _0511_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__buf_2
XFILLER_9_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0824_ _0362_ _0361_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__xnor2_1
X_0755_ _0167_ _0290_ _0287_ _0293_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__a31o_1
X_0686_ _0199_ CIRCUIT_1957.int_memory_1.div_1.A4 vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__and2b_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1169_ CIRCUIT_1957.GATES_38.result CIRCUIT_1957.GATES_35.result _0013_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_71.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1030__B1 _0520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0540_ CIRCUIT_1957.MEMORY_75.s_currentState CIRCUIT_1957.MEMORY_83.s_currentState
+ _0104_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__mux2_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1088__B1 _0523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0994__A clknet_1_0__leaf__0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1023_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[2\] _0512_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0031_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result
+ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result
+ sky130_fd_sc_hd__clkbuf_16
X_0807_ _0317_ _0318_ _0321_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__a31o_1
X_0738_ _0271_ _0275_ _0276_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__a21oi_1
X_0669_ CIRCUIT_1957.int_memory_1.div_1.B1 _0206_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__nor2_1
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ _0121_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result CIRCUIT_1957.int_memory_1.GATES_32.result
+ vssd1 vssd1 vccd1 vccd1 clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result sky130_fd_sc_hd__clkbuf_16
XFILLER_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0986__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0986_ clknet_1_1__leaf__0142_ _0496_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__nand2_2
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0771_ _0305_ _0308_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__nor2_1
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0840_ _0099_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1185_ net46 _0059_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0969_ _0492_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.GATES_28.result sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1112__A2 _0533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0823_ _0351_ _0357_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__nand2_1
X_0685_ CIRCUIT_1957.int_memory_1.div_1.A4 _0199_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__and2b_1
X_0754_ _0167_ _0292_ _0290_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1099_ CIRCUIT_1957.int_memory_1.mul2_1.A3 _0532_ _0517_ vssd1 vssd1 vccd1 vccd1
+ _0080_ sky130_fd_sc_hd__a21o_1
X_1168_ CIRCUIT_1957.GATES_41.result CIRCUIT_1957.GATES_27.result _0012_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_1957.MEMORY_72.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0994__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1022_ CIRCUIT_1957.int_memory_1.GATES_4.input2\[1\] _0512_ _0523_ vssd1 vssd1 vccd1
+ vccd1 _0030_ sky130_fd_sc_hd__a21o_1
X_0668_ _0162_ _0206_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__nand2_1
X_0806_ _0330_ _0336_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__or3_1
X_0737_ _0231_ _0273_ _0274_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__and3_1
X_0599_ _0147_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.D2 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0989__B _0496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1005_ _0510_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_1957.int_memory_1.GATES_53.result sky130_fd_sc_hd__buf_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

