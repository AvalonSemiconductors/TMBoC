magic
tech sky130B
magscale 1 2
timestamp 1674825766
<< viali >>
rect 2605 26537 2639 26571
rect 5181 26537 5215 26571
rect 9321 26537 9355 26571
rect 20361 26537 20395 26571
rect 23673 26537 23707 26571
rect 26525 26537 26559 26571
rect 15301 26401 15335 26435
rect 1685 26333 1719 26367
rect 2789 26333 2823 26367
rect 4997 26333 5031 26367
rect 5825 26333 5859 26367
rect 6561 26333 6595 26367
rect 6745 26333 6779 26367
rect 9137 26333 9171 26367
rect 9873 26333 9907 26367
rect 10057 26333 10091 26367
rect 11805 26333 11839 26367
rect 12357 26333 12391 26367
rect 14289 26333 14323 26367
rect 16865 26333 16899 26367
rect 19533 26333 19567 26367
rect 20177 26333 20211 26367
rect 23489 26333 23523 26367
rect 26341 26333 26375 26367
rect 2053 26265 2087 26299
rect 5733 26265 5767 26299
rect 13369 26265 13403 26299
rect 16129 26265 16163 26299
rect 19441 26265 19475 26299
rect 6561 26197 6595 26231
rect 9965 26197 9999 26231
rect 14473 26197 14507 26231
rect 17049 26197 17083 26231
rect 1685 25993 1719 26027
rect 4537 25993 4571 26027
rect 5089 25993 5123 26027
rect 8677 25993 8711 26027
rect 10149 25993 10183 26027
rect 2605 25857 2639 25891
rect 4445 25857 4479 25891
rect 4629 25857 4663 25891
rect 5457 25857 5491 25891
rect 6745 25857 6779 25891
rect 8309 25857 8343 25891
rect 9781 25857 9815 25891
rect 10793 25857 10827 25891
rect 12081 25857 12115 25891
rect 12725 25857 12759 25891
rect 15485 25857 15519 25891
rect 17141 25857 17175 25891
rect 18797 25857 18831 25891
rect 2513 25789 2547 25823
rect 5365 25789 5399 25823
rect 8217 25789 8251 25823
rect 9873 25789 9907 25823
rect 10701 25789 10735 25823
rect 12817 25789 12851 25823
rect 13277 25789 13311 25823
rect 13553 25789 13587 25823
rect 15025 25789 15059 25823
rect 16221 25789 16255 25823
rect 19809 25789 19843 25823
rect 20637 25789 20671 25823
rect 11161 25721 11195 25755
rect 2237 25653 2271 25687
rect 6745 25653 6779 25687
rect 11897 25653 11931 25687
rect 15485 25653 15519 25687
rect 17141 25653 17175 25687
rect 18613 25653 18647 25687
rect 4813 25449 4847 25483
rect 13645 25449 13679 25483
rect 3433 25381 3467 25415
rect 4353 25381 4387 25415
rect 5733 25381 5767 25415
rect 7389 25381 7423 25415
rect 7481 25381 7515 25415
rect 9413 25381 9447 25415
rect 11069 25381 11103 25415
rect 6009 25313 6043 25347
rect 7021 25313 7055 25347
rect 8217 25313 8251 25347
rect 11897 25313 11931 25347
rect 19441 25313 19475 25347
rect 19717 25313 19751 25347
rect 21189 25313 21223 25347
rect 2053 25245 2087 25279
rect 4353 25245 4387 25279
rect 5089 25245 5123 25279
rect 5217 25245 5251 25279
rect 5917 25245 5951 25279
rect 8028 25245 8062 25279
rect 9229 25245 9263 25279
rect 9321 25245 9355 25279
rect 9505 25245 9539 25279
rect 9689 25245 9723 25279
rect 10609 25245 10643 25279
rect 10885 25245 10919 25279
rect 15209 25245 15243 25279
rect 17417 25245 17451 25279
rect 18153 25245 18187 25279
rect 18889 25245 18923 25279
rect 2298 25177 2332 25211
rect 4813 25177 4847 25211
rect 4997 25177 5031 25211
rect 8125 25177 8159 25211
rect 8217 25177 8251 25211
rect 8401 25177 8435 25211
rect 12173 25177 12207 25211
rect 14933 25177 14967 25211
rect 17141 25177 17175 25211
rect 18613 25177 18647 25211
rect 6377 25109 6411 25143
rect 10701 25109 10735 25143
rect 14289 25109 14323 25143
rect 15669 25109 15703 25143
rect 17969 25109 18003 25143
rect 2237 24905 2271 24939
rect 5457 24905 5491 24939
rect 5733 24905 5767 24939
rect 9137 24905 9171 24939
rect 9873 24905 9907 24939
rect 11161 24905 11195 24939
rect 20729 24905 20763 24939
rect 4721 24837 4755 24871
rect 9229 24837 9263 24871
rect 9413 24837 9447 24871
rect 14841 24837 14875 24871
rect 17141 24837 17175 24871
rect 17601 24837 17635 24871
rect 18613 24837 18647 24871
rect 3361 24769 3395 24803
rect 4445 24769 4479 24803
rect 4629 24769 4663 24803
rect 4813 24769 4847 24803
rect 5641 24769 5675 24803
rect 5825 24769 5859 24803
rect 7021 24769 7055 24803
rect 7277 24769 7311 24803
rect 9045 24769 9079 24803
rect 10793 24769 10827 24803
rect 10977 24769 11011 24803
rect 12081 24769 12115 24803
rect 13093 24769 13127 24803
rect 14105 24769 14139 24803
rect 16865 24769 16899 24803
rect 17693 24769 17727 24803
rect 18337 24769 18371 24803
rect 20913 24769 20947 24803
rect 3617 24701 3651 24735
rect 10333 24701 10367 24735
rect 14565 24701 14599 24735
rect 16313 24701 16347 24735
rect 6009 24633 6043 24667
rect 8861 24633 8895 24667
rect 9965 24633 9999 24667
rect 4997 24565 5031 24599
rect 8401 24565 8435 24599
rect 12081 24565 12115 24599
rect 20085 24565 20119 24599
rect 3985 24361 4019 24395
rect 7297 24361 7331 24395
rect 8585 24361 8619 24395
rect 10977 24361 11011 24395
rect 13369 24361 13403 24395
rect 14381 24361 14415 24395
rect 15117 24361 15151 24395
rect 6745 24293 6779 24327
rect 4261 24225 4295 24259
rect 5365 24225 5399 24259
rect 9137 24225 9171 24259
rect 11897 24225 11931 24259
rect 16589 24225 16623 24259
rect 17141 24225 17175 24259
rect 17417 24225 17451 24259
rect 20269 24225 20303 24259
rect 1961 24157 1995 24191
rect 2228 24157 2262 24191
rect 4353 24157 4387 24191
rect 7205 24157 7239 24191
rect 7408 24157 7442 24191
rect 7573 24157 7607 24191
rect 8033 24157 8067 24191
rect 8401 24157 8435 24191
rect 10977 24157 11011 24191
rect 11161 24157 11195 24191
rect 11621 24157 11655 24191
rect 14565 24157 14599 24191
rect 15669 24157 15703 24191
rect 21005 24157 21039 24191
rect 5632 24089 5666 24123
rect 8217 24089 8251 24123
rect 8309 24089 8343 24123
rect 9404 24089 9438 24123
rect 19717 24089 19751 24123
rect 21281 24089 21315 24123
rect 3341 24021 3375 24055
rect 7297 24021 7331 24055
rect 10517 24021 10551 24055
rect 18889 24021 18923 24055
rect 1685 23817 1719 23851
rect 5825 23817 5859 23851
rect 6929 23817 6963 23851
rect 7757 23817 7791 23851
rect 8677 23817 8711 23851
rect 8861 23817 8895 23851
rect 9413 23817 9447 23851
rect 13461 23817 13495 23851
rect 18153 23817 18187 23851
rect 20361 23817 20395 23851
rect 8493 23749 8527 23783
rect 8585 23749 8619 23783
rect 14749 23749 14783 23783
rect 19073 23749 19107 23783
rect 2809 23681 2843 23715
rect 3525 23681 3559 23715
rect 4712 23681 4746 23715
rect 7113 23681 7147 23715
rect 7573 23681 7607 23715
rect 9597 23681 9631 23715
rect 12081 23681 12115 23715
rect 16865 23681 16899 23715
rect 3065 23613 3099 23647
rect 4445 23613 4479 23647
rect 11989 23613 12023 23647
rect 8309 23545 8343 23579
rect 3709 23477 3743 23511
rect 10517 23477 10551 23511
rect 11161 23477 11195 23511
rect 12449 23477 12483 23511
rect 5641 23273 5675 23307
rect 7757 23273 7791 23307
rect 9505 23273 9539 23307
rect 16865 23273 16899 23307
rect 21207 23273 21241 23307
rect 21925 23273 21959 23307
rect 10701 23205 10735 23239
rect 4261 23137 4295 23171
rect 11345 23137 11379 23171
rect 13185 23137 13219 23171
rect 14749 23137 14783 23171
rect 15025 23137 15059 23171
rect 18521 23137 18555 23171
rect 21465 23137 21499 23171
rect 3085 23069 3119 23103
rect 3341 23069 3375 23103
rect 6377 23069 6411 23103
rect 8217 23069 8251 23103
rect 10241 23069 10275 23103
rect 11161 23069 11195 23103
rect 12173 23069 12207 23103
rect 14657 23069 14691 23103
rect 16773 23069 16807 23103
rect 16865 23069 16899 23103
rect 17601 23069 17635 23103
rect 21925 23069 21959 23103
rect 4528 23001 4562 23035
rect 6622 23001 6656 23035
rect 11069 23001 11103 23035
rect 16589 23001 16623 23035
rect 1961 22933 1995 22967
rect 8401 22933 8435 22967
rect 10057 22933 10091 22967
rect 13737 22933 13771 22967
rect 17049 22933 17083 22967
rect 19717 22933 19751 22967
rect 3433 22729 3467 22763
rect 8309 22729 8343 22763
rect 11161 22729 11195 22763
rect 11805 22729 11839 22763
rect 15025 22729 15059 22763
rect 10048 22661 10082 22695
rect 13369 22661 13403 22695
rect 14933 22661 14967 22695
rect 20821 22661 20855 22695
rect 2145 22593 2179 22627
rect 6929 22593 6963 22627
rect 7196 22593 7230 22627
rect 11897 22593 11931 22627
rect 12541 22593 12575 22627
rect 13461 22593 13495 22627
rect 15945 22593 15979 22627
rect 17601 22593 17635 22627
rect 19080 22593 19114 22627
rect 19809 22593 19843 22627
rect 2053 22525 2087 22559
rect 9321 22525 9355 22559
rect 9781 22525 9815 22559
rect 12449 22525 12483 22559
rect 12909 22525 12943 22559
rect 15117 22525 15151 22559
rect 15853 22525 15887 22559
rect 16313 22525 16347 22559
rect 17233 22525 17267 22559
rect 17509 22525 17543 22559
rect 18705 22525 18739 22559
rect 18981 22525 19015 22559
rect 1777 22389 1811 22423
rect 4353 22389 4387 22423
rect 5181 22389 5215 22423
rect 14565 22389 14599 22423
rect 21373 22389 21407 22423
rect 22017 22389 22051 22423
rect 5733 22185 5767 22219
rect 7205 22185 7239 22219
rect 13737 22185 13771 22219
rect 15669 22185 15703 22219
rect 11437 22117 11471 22151
rect 4261 22049 4295 22083
rect 12449 22049 12483 22083
rect 20085 22049 20119 22083
rect 20361 22049 20395 22083
rect 3985 21981 4019 22015
rect 8318 21981 8352 22015
rect 8585 21981 8619 22015
rect 9413 21981 9447 22015
rect 10057 21981 10091 22015
rect 13553 21981 13587 22015
rect 14289 21981 14323 22015
rect 14545 21981 14579 22015
rect 16221 21981 16255 22015
rect 16865 21981 16899 22015
rect 20453 21981 20487 22015
rect 21097 21981 21131 22015
rect 21741 21981 21775 22015
rect 22008 21981 22042 22015
rect 10302 21913 10336 21947
rect 12357 21913 12391 21947
rect 17110 21913 17144 21947
rect 1685 21845 1719 21879
rect 2605 21845 2639 21879
rect 3249 21845 3283 21879
rect 6653 21845 6687 21879
rect 9597 21845 9631 21879
rect 11897 21845 11931 21879
rect 12265 21845 12299 21879
rect 16405 21845 16439 21879
rect 18245 21845 18279 21879
rect 18705 21845 18739 21879
rect 19533 21845 19567 21879
rect 21281 21845 21315 21879
rect 23121 21845 23155 21879
rect 4123 21641 4157 21675
rect 5365 21641 5399 21675
rect 14933 21641 14967 21675
rect 16957 21641 16991 21675
rect 17417 21641 17451 21675
rect 19533 21641 19567 21675
rect 23397 21641 23431 21675
rect 17325 21573 17359 21607
rect 22262 21573 22296 21607
rect 4813 21505 4847 21539
rect 5365 21505 5399 21539
rect 5549 21505 5583 21539
rect 10048 21505 10082 21539
rect 12173 21505 12207 21539
rect 13809 21505 13843 21539
rect 15393 21505 15427 21539
rect 15669 21505 15703 21539
rect 18153 21505 18187 21539
rect 18889 21505 18923 21539
rect 20657 21505 20691 21539
rect 22017 21505 22051 21539
rect 2329 21437 2363 21471
rect 2697 21437 2731 21471
rect 4629 21437 4663 21471
rect 6561 21437 6595 21471
rect 6837 21437 6871 21471
rect 9781 21437 9815 21471
rect 12081 21437 12115 21471
rect 12541 21437 12575 21471
rect 13553 21437 13587 21471
rect 15485 21437 15519 21471
rect 17509 21437 17543 21471
rect 20913 21437 20947 21471
rect 11161 21369 11195 21403
rect 13001 21369 13035 21403
rect 1593 21301 1627 21335
rect 8309 21301 8343 21335
rect 9229 21301 9263 21335
rect 15393 21301 15427 21335
rect 15853 21301 15887 21335
rect 18337 21301 18371 21335
rect 19073 21301 19107 21335
rect 21373 21301 21407 21335
rect 1639 21097 1673 21131
rect 6883 21097 6917 21131
rect 7481 21097 7515 21131
rect 10149 21097 10183 21131
rect 13093 21097 13127 21131
rect 16865 21097 16899 21131
rect 20913 21097 20947 21131
rect 21373 21097 21407 21131
rect 10793 21029 10827 21063
rect 14289 21029 14323 21063
rect 3433 20961 3467 20995
rect 11253 20961 11287 20995
rect 11437 20961 11471 20995
rect 14933 20961 14967 20995
rect 15853 20961 15887 20995
rect 18337 20961 18371 20995
rect 3065 20893 3099 20927
rect 4445 20893 4479 20927
rect 4629 20893 4663 20927
rect 5089 20893 5123 20927
rect 5457 20893 5491 20927
rect 7389 20893 7423 20927
rect 7573 20893 7607 20927
rect 10333 20893 10367 20927
rect 12357 20893 12391 20927
rect 12909 20893 12943 20927
rect 13553 20893 13587 20927
rect 14749 20893 14783 20927
rect 16037 20893 16071 20927
rect 16129 20893 16163 20927
rect 18613 20893 18647 20927
rect 19533 20893 19567 20927
rect 19789 20893 19823 20927
rect 21557 20893 21591 20927
rect 22201 20893 22235 20927
rect 14657 20825 14691 20859
rect 22468 20825 22502 20859
rect 4629 20757 4663 20791
rect 8033 20757 8067 20791
rect 9689 20757 9723 20791
rect 11161 20757 11195 20791
rect 13737 20757 13771 20791
rect 16129 20757 16163 20791
rect 23581 20757 23615 20791
rect 2789 20553 2823 20587
rect 3433 20553 3467 20587
rect 5733 20553 5767 20587
rect 6561 20553 6595 20587
rect 11069 20553 11103 20587
rect 12725 20553 12759 20587
rect 14289 20553 14323 20587
rect 16313 20553 16347 20587
rect 20085 20553 20119 20587
rect 20545 20553 20579 20587
rect 23489 20553 23523 20587
rect 11805 20485 11839 20519
rect 14657 20485 14691 20519
rect 15945 20485 15979 20519
rect 17325 20485 17359 20519
rect 22569 20485 22603 20519
rect 1685 20417 1719 20451
rect 2697 20417 2731 20451
rect 2881 20417 2915 20451
rect 3341 20417 3375 20451
rect 3525 20417 3559 20451
rect 3985 20417 4019 20451
rect 6561 20417 6595 20451
rect 6745 20417 6779 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 10149 20417 10183 20451
rect 10277 20417 10311 20451
rect 13461 20417 13495 20451
rect 14749 20417 14783 20451
rect 15669 20417 15703 20451
rect 15817 20417 15851 20451
rect 16037 20417 16071 20451
rect 16175 20417 16209 20451
rect 18337 20417 18371 20451
rect 20177 20417 20211 20451
rect 21005 20417 21039 20451
rect 22661 20417 22695 20451
rect 23673 20417 23707 20451
rect 4261 20349 4295 20383
rect 9965 20349 9999 20383
rect 13369 20349 13403 20383
rect 14933 20349 14967 20383
rect 19901 20349 19935 20383
rect 22385 20349 22419 20383
rect 9321 20281 9355 20315
rect 13829 20281 13863 20315
rect 21189 20281 21223 20315
rect 23029 20281 23063 20315
rect 1777 20213 1811 20247
rect 7573 20213 7607 20247
rect 8309 20213 8343 20247
rect 8861 20213 8895 20247
rect 11897 20213 11931 20247
rect 18889 20213 18923 20247
rect 24133 20213 24167 20247
rect 24685 20213 24719 20247
rect 10609 20009 10643 20043
rect 13645 20009 13679 20043
rect 15669 20009 15703 20043
rect 16129 20009 16163 20043
rect 16957 20009 16991 20043
rect 17877 20009 17911 20043
rect 18521 20009 18555 20043
rect 19809 20009 19843 20043
rect 25145 20009 25179 20043
rect 6101 19941 6135 19975
rect 1593 19873 1627 19907
rect 6745 19873 6779 19907
rect 12357 19873 12391 19907
rect 20361 19873 20395 19907
rect 24685 19873 24719 19907
rect 1860 19805 1894 19839
rect 7389 19805 7423 19839
rect 7573 19805 7607 19839
rect 9321 19805 9355 19839
rect 10425 19805 10459 19839
rect 11069 19805 11103 19839
rect 12265 19805 12299 19839
rect 13553 19805 13587 19839
rect 14289 19805 14323 19839
rect 16497 19805 16531 19839
rect 17785 19805 17819 19839
rect 17969 19805 18003 19839
rect 18429 19805 18463 19839
rect 18613 19805 18647 19839
rect 20269 19805 20303 19839
rect 22937 19805 22971 19839
rect 23581 19805 23615 19839
rect 24777 19805 24811 19839
rect 26341 19805 26375 19839
rect 5549 19737 5583 19771
rect 6561 19737 6595 19771
rect 10057 19737 10091 19771
rect 11345 19737 11379 19771
rect 12173 19737 12207 19771
rect 14534 19737 14568 19771
rect 16313 19737 16347 19771
rect 17141 19737 17175 19771
rect 17325 19737 17359 19771
rect 22692 19737 22726 19771
rect 2973 19669 3007 19703
rect 4445 19669 4479 19703
rect 5089 19669 5123 19703
rect 6469 19669 6503 19703
rect 7573 19669 7607 19703
rect 8585 19669 8619 19703
rect 9137 19669 9171 19703
rect 10241 19669 10275 19703
rect 10333 19669 10367 19703
rect 11805 19669 11839 19703
rect 13093 19669 13127 19703
rect 20177 19669 20211 19703
rect 21005 19669 21039 19703
rect 21557 19669 21591 19703
rect 23397 19669 23431 19703
rect 26525 19669 26559 19703
rect 1593 19465 1627 19499
rect 3985 19465 4019 19499
rect 5917 19465 5951 19499
rect 7113 19465 7147 19499
rect 9597 19465 9631 19499
rect 10057 19465 10091 19499
rect 11713 19465 11747 19499
rect 12541 19465 12575 19499
rect 18613 19465 18647 19499
rect 20637 19465 20671 19499
rect 22293 19465 22327 19499
rect 22753 19465 22787 19499
rect 25881 19465 25915 19499
rect 2728 19397 2762 19431
rect 10517 19397 10551 19431
rect 15853 19397 15887 19431
rect 15945 19397 15979 19431
rect 19533 19397 19567 19431
rect 22385 19397 22419 19431
rect 4169 19329 4203 19363
rect 5273 19329 5307 19363
rect 7021 19329 7055 19363
rect 10425 19329 10459 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 12357 19329 12391 19363
rect 13001 19329 13035 19363
rect 17049 19329 17083 19363
rect 18429 19329 18463 19363
rect 19441 19329 19475 19363
rect 20453 19329 20487 19363
rect 21097 19329 21131 19363
rect 23489 19329 23523 19363
rect 23673 19329 23707 19363
rect 24133 19329 24167 19363
rect 26341 19329 26375 19363
rect 2973 19261 3007 19295
rect 7297 19261 7331 19295
rect 7849 19261 7883 19295
rect 8125 19261 8159 19295
rect 10701 19261 10735 19295
rect 15669 19261 15703 19295
rect 18245 19261 18279 19295
rect 19717 19261 19751 19295
rect 20269 19261 20303 19295
rect 22109 19261 22143 19295
rect 24409 19261 24443 19295
rect 14289 19193 14323 19227
rect 16313 19193 16347 19227
rect 4721 19125 4755 19159
rect 5457 19125 5491 19159
rect 6653 19125 6687 19159
rect 16865 19125 16899 19159
rect 17509 19125 17543 19159
rect 19073 19125 19107 19159
rect 21281 19125 21315 19159
rect 26525 19125 26559 19159
rect 4997 18921 5031 18955
rect 9873 18921 9907 18955
rect 13093 18921 13127 18955
rect 15577 18921 15611 18955
rect 20821 18921 20855 18955
rect 23765 18853 23799 18887
rect 6745 18785 6779 18819
rect 8493 18785 8527 18819
rect 11713 18785 11747 18819
rect 14657 18785 14691 18819
rect 19441 18785 19475 18819
rect 21557 18785 21591 18819
rect 21833 18785 21867 18819
rect 25605 18785 25639 18819
rect 4261 18717 4295 18751
rect 4445 18717 4479 18751
rect 7205 18717 7239 18751
rect 8217 18717 8251 18751
rect 9413 18717 9447 18751
rect 11253 18717 11287 18751
rect 13737 18717 13771 18751
rect 14381 18717 14415 18751
rect 14473 18717 14507 18751
rect 16701 18717 16735 18751
rect 16957 18717 16991 18751
rect 17877 18717 17911 18751
rect 18705 18717 18739 18751
rect 23765 18717 23799 18751
rect 24685 18717 24719 18751
rect 26433 18717 26467 18751
rect 26893 18717 26927 18751
rect 4353 18649 4387 18683
rect 6469 18649 6503 18683
rect 8309 18649 8343 18683
rect 11008 18649 11042 18683
rect 11958 18649 11992 18683
rect 19686 18649 19720 18683
rect 26157 18649 26191 18683
rect 27169 18649 27203 18683
rect 1777 18581 1811 18615
rect 2329 18581 2363 18615
rect 2881 18581 2915 18615
rect 3433 18581 3467 18615
rect 7389 18581 7423 18615
rect 7849 18581 7883 18615
rect 9229 18581 9263 18615
rect 13645 18581 13679 18615
rect 18061 18581 18095 18615
rect 18889 18581 18923 18615
rect 23305 18581 23339 18615
rect 4261 18377 4295 18411
rect 6561 18377 6595 18411
rect 9137 18377 9171 18411
rect 10977 18377 11011 18411
rect 12541 18377 12575 18411
rect 14473 18377 14507 18411
rect 20177 18377 20211 18411
rect 23581 18377 23615 18411
rect 24133 18377 24167 18411
rect 5733 18309 5767 18343
rect 7665 18309 7699 18343
rect 9842 18309 9876 18343
rect 11989 18309 12023 18343
rect 13185 18309 13219 18343
rect 22845 18309 22879 18343
rect 3341 18241 3375 18275
rect 6745 18241 6779 18275
rect 12173 18241 12207 18275
rect 12725 18241 12759 18275
rect 15669 18241 15703 18275
rect 16129 18241 16163 18275
rect 17141 18241 17175 18275
rect 17693 18241 17727 18275
rect 18429 18241 18463 18275
rect 20913 18241 20947 18275
rect 22109 18241 22143 18275
rect 3709 18173 3743 18207
rect 6009 18173 6043 18207
rect 7389 18173 7423 18207
rect 9597 18173 9631 18207
rect 12432 18173 12466 18207
rect 12633 18173 12667 18207
rect 18705 18173 18739 18207
rect 20637 18173 20671 18207
rect 25053 18173 25087 18207
rect 25789 18173 25823 18207
rect 26525 18173 26559 18207
rect 16221 18105 16255 18139
rect 1915 18037 1949 18071
rect 15485 18037 15519 18071
rect 16957 18037 16991 18071
rect 17693 18037 17727 18071
rect 21373 18037 21407 18071
rect 5779 17833 5813 17867
rect 7481 17833 7515 17867
rect 8585 17833 8619 17867
rect 10701 17833 10735 17867
rect 15393 17833 15427 17867
rect 18797 17833 18831 17867
rect 25605 17833 25639 17867
rect 1685 17697 1719 17731
rect 1961 17697 1995 17731
rect 3433 17697 3467 17731
rect 4353 17697 4387 17731
rect 9505 17697 9539 17731
rect 11713 17697 11747 17731
rect 12909 17697 12943 17731
rect 15945 17697 15979 17731
rect 22201 17697 22235 17731
rect 22477 17697 22511 17731
rect 27077 17697 27111 17731
rect 27353 17697 27387 17731
rect 3985 17629 4019 17663
rect 7389 17629 7423 17663
rect 7573 17629 7607 17663
rect 9229 17629 9263 17663
rect 10517 17629 10551 17663
rect 11529 17629 11563 17663
rect 14473 17629 14507 17663
rect 14841 17629 14875 17663
rect 15301 17629 15335 17663
rect 15485 17629 15519 17663
rect 18705 17629 18739 17663
rect 18889 17629 18923 17663
rect 19625 17629 19659 17663
rect 20453 17629 20487 17663
rect 20637 17629 20671 17663
rect 21189 17629 21223 17663
rect 22109 17629 22143 17663
rect 23121 17629 23155 17663
rect 23673 17629 23707 17663
rect 24685 17629 24719 17663
rect 6377 17561 6411 17595
rect 13461 17561 13495 17595
rect 14565 17561 14599 17595
rect 14657 17561 14691 17595
rect 16221 17561 16255 17595
rect 19809 17561 19843 17595
rect 6929 17493 6963 17527
rect 11161 17493 11195 17527
rect 11621 17493 11655 17527
rect 14289 17493 14323 17527
rect 17693 17493 17727 17527
rect 18153 17493 18187 17527
rect 19993 17493 20027 17527
rect 20545 17493 20579 17527
rect 21281 17493 21315 17527
rect 22937 17493 22971 17527
rect 23857 17493 23891 17527
rect 24685 17493 24719 17527
rect 2513 17289 2547 17323
rect 3065 17289 3099 17323
rect 4077 17289 4111 17323
rect 4629 17289 4663 17323
rect 6561 17289 6595 17323
rect 10977 17289 11011 17323
rect 14289 17289 14323 17323
rect 25697 17289 25731 17323
rect 9873 17221 9907 17255
rect 10885 17221 10919 17255
rect 11713 17221 11747 17255
rect 19349 17221 19383 17255
rect 20453 17221 20487 17255
rect 24225 17221 24259 17255
rect 1593 17153 1627 17187
rect 3065 17153 3099 17187
rect 3249 17153 3283 17187
rect 3893 17153 3927 17187
rect 4077 17153 4111 17187
rect 4537 17153 4571 17187
rect 4721 17153 4755 17187
rect 5641 17153 5675 17187
rect 7674 17153 7708 17187
rect 9781 17153 9815 17187
rect 10793 17153 10827 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 14841 17153 14875 17187
rect 16865 17153 16899 17187
rect 17693 17153 17727 17187
rect 20085 17153 20119 17187
rect 20178 17153 20212 17187
rect 20361 17153 20395 17187
rect 20550 17153 20584 17187
rect 21189 17153 21223 17187
rect 23949 17153 23983 17187
rect 26433 17153 26467 17187
rect 7941 17085 7975 17119
rect 9965 17085 9999 17119
rect 11161 17085 11195 17119
rect 12541 17085 12575 17119
rect 12817 17085 12851 17119
rect 15761 17085 15795 17119
rect 17601 17085 17635 17119
rect 18061 17085 18095 17119
rect 18797 17085 18831 17119
rect 21465 17085 21499 17119
rect 22477 17085 22511 17119
rect 23305 17085 23339 17119
rect 1777 17017 1811 17051
rect 9413 17017 9447 17051
rect 10609 17017 10643 17051
rect 17049 17017 17083 17051
rect 21281 17017 21315 17051
rect 5733 16949 5767 16983
rect 8861 16949 8895 16983
rect 20729 16949 20763 16983
rect 21373 16949 21407 16983
rect 26341 16949 26375 16983
rect 4169 16745 4203 16779
rect 6745 16745 6779 16779
rect 10701 16745 10735 16779
rect 23397 16745 23431 16779
rect 4997 16609 5031 16643
rect 8033 16609 8067 16643
rect 9965 16609 9999 16643
rect 14289 16609 14323 16643
rect 17601 16609 17635 16643
rect 18429 16609 18463 16643
rect 23489 16609 23523 16643
rect 24869 16609 24903 16643
rect 26433 16609 26467 16643
rect 2237 16541 2271 16575
rect 2973 16541 3007 16575
rect 3985 16541 4019 16575
rect 5733 16541 5767 16575
rect 6653 16541 6687 16575
rect 9781 16541 9815 16575
rect 13737 16541 13771 16575
rect 14657 16541 14691 16575
rect 19625 16541 19659 16575
rect 20453 16541 20487 16575
rect 21189 16541 21223 16575
rect 23673 16541 23707 16575
rect 7757 16473 7791 16507
rect 9873 16473 9907 16507
rect 11253 16473 11287 16507
rect 14565 16473 14599 16507
rect 14774 16473 14808 16507
rect 15393 16473 15427 16507
rect 23397 16473 23431 16507
rect 25697 16473 25731 16507
rect 26985 16473 27019 16507
rect 2053 16405 2087 16439
rect 2789 16405 2823 16439
rect 5549 16405 5583 16439
rect 9413 16405 9447 16439
rect 12541 16405 12575 16439
rect 13553 16405 13587 16439
rect 14933 16405 14967 16439
rect 16681 16405 16715 16439
rect 22477 16405 22511 16439
rect 23857 16405 23891 16439
rect 3617 16201 3651 16235
rect 4261 16201 4295 16235
rect 8217 16201 8251 16235
rect 10057 16201 10091 16235
rect 12449 16201 12483 16235
rect 15945 16201 15979 16235
rect 17325 16201 17359 16235
rect 17417 16201 17451 16235
rect 18705 16201 18739 16235
rect 21281 16201 21315 16235
rect 27169 16201 27203 16235
rect 2145 16133 2179 16167
rect 8922 16133 8956 16167
rect 10885 16133 10919 16167
rect 13737 16133 13771 16167
rect 14473 16133 14507 16167
rect 19993 16133 20027 16167
rect 24225 16133 24259 16167
rect 26525 16133 26559 16167
rect 6009 16065 6043 16099
rect 6561 16065 6595 16099
rect 7389 16065 7423 16099
rect 8033 16065 8067 16099
rect 10793 16065 10827 16099
rect 11161 16065 11195 16099
rect 20913 16065 20947 16099
rect 22017 16065 22051 16099
rect 26433 16065 26467 16099
rect 1869 15997 1903 16031
rect 5733 15997 5767 16031
rect 8677 15997 8711 16031
rect 10676 15997 10710 16031
rect 14197 15997 14231 16031
rect 17233 15997 17267 16031
rect 20637 15997 20671 16031
rect 20821 15997 20855 16031
rect 22293 15997 22327 16031
rect 6561 15929 6595 15963
rect 23765 15929 23799 15963
rect 7573 15861 7607 15895
rect 10517 15861 10551 15895
rect 17785 15861 17819 15895
rect 25513 15861 25547 15895
rect 4169 15657 4203 15691
rect 9229 15657 9263 15691
rect 13277 15657 13311 15691
rect 14841 15657 14875 15691
rect 16957 15657 16991 15691
rect 18889 15657 18923 15691
rect 20085 15657 20119 15691
rect 22477 15657 22511 15691
rect 24869 15657 24903 15691
rect 7757 15589 7791 15623
rect 11529 15589 11563 15623
rect 24593 15589 24627 15623
rect 10701 15521 10735 15555
rect 18429 15521 18463 15555
rect 22017 15521 22051 15555
rect 23397 15521 23431 15555
rect 23673 15521 23707 15555
rect 25513 15521 25547 15555
rect 25789 15521 25823 15555
rect 1685 15453 1719 15487
rect 4905 15453 4939 15487
rect 5549 15453 5583 15487
rect 7757 15453 7791 15487
rect 9137 15453 9171 15487
rect 10609 15453 10643 15487
rect 10977 15453 11011 15487
rect 11253 15453 11287 15487
rect 14289 15453 14323 15487
rect 14565 15453 14599 15487
rect 14709 15453 14743 15487
rect 15669 15453 15703 15487
rect 18521 15453 18555 15487
rect 19625 15453 19659 15487
rect 21465 15453 21499 15487
rect 22109 15453 22143 15487
rect 23305 15453 23339 15487
rect 24777 15453 24811 15487
rect 24869 15453 24903 15487
rect 1961 15385 1995 15419
rect 4077 15385 4111 15419
rect 5825 15385 5859 15419
rect 11989 15385 12023 15419
rect 14473 15385 14507 15419
rect 21220 15385 21254 15419
rect 25053 15385 25087 15419
rect 3433 15317 3467 15351
rect 4997 15317 5031 15351
rect 7297 15317 7331 15351
rect 8493 15317 8527 15351
rect 9597 15317 9631 15351
rect 19441 15317 19475 15351
rect 27261 15317 27295 15351
rect 3709 15113 3743 15147
rect 6653 15113 6687 15147
rect 8033 15113 8067 15147
rect 10517 15113 10551 15147
rect 12081 15113 12115 15147
rect 13461 15113 13495 15147
rect 17509 15113 17543 15147
rect 19717 15113 19751 15147
rect 27169 15113 27203 15147
rect 2145 15045 2179 15079
rect 2881 15045 2915 15079
rect 14749 15045 14783 15079
rect 15853 15045 15887 15079
rect 18644 15045 18678 15079
rect 19533 15045 19567 15079
rect 22477 15045 22511 15079
rect 2237 14977 2271 15011
rect 3157 14977 3191 15011
rect 3801 14977 3835 15011
rect 6745 14977 6779 15011
rect 7297 14977 7331 15011
rect 8493 14977 8527 15011
rect 9393 14977 9427 15011
rect 10977 14977 11011 15011
rect 15945 14977 15979 15011
rect 17049 14977 17083 15011
rect 18889 14977 18923 15011
rect 19349 14977 19383 15011
rect 20453 14977 20487 15011
rect 22385 14977 22419 15011
rect 23397 14977 23431 15011
rect 24409 14977 24443 15011
rect 25513 14977 25547 15011
rect 4261 14909 4295 14943
rect 4537 14909 4571 14943
rect 9137 14909 9171 14943
rect 12173 14909 12207 14943
rect 12265 14909 12299 14943
rect 15761 14909 15795 14943
rect 20177 14909 20211 14943
rect 22569 14909 22603 14943
rect 23305 14909 23339 14943
rect 24317 14909 24351 14943
rect 24777 14909 24811 14943
rect 26525 14909 26559 14943
rect 6009 14841 6043 14875
rect 16313 14841 16347 14875
rect 23765 14841 23799 14875
rect 1685 14773 1719 14807
rect 7389 14773 7423 14807
rect 8585 14773 8619 14807
rect 11161 14773 11195 14807
rect 11713 14773 11747 14807
rect 16865 14773 16899 14807
rect 22017 14773 22051 14807
rect 4261 14569 4295 14603
rect 4997 14569 5031 14603
rect 5641 14569 5675 14603
rect 13737 14569 13771 14603
rect 17601 14569 17635 14603
rect 19533 14569 19567 14603
rect 22477 14569 22511 14603
rect 24593 14569 24627 14603
rect 8585 14501 8619 14535
rect 15025 14501 15059 14535
rect 18889 14501 18923 14535
rect 20085 14501 20119 14535
rect 7021 14433 7055 14467
rect 15117 14433 15151 14467
rect 18337 14433 18371 14467
rect 23029 14433 23063 14467
rect 3433 14365 3467 14399
rect 4445 14365 4479 14399
rect 4905 14365 4939 14399
rect 5825 14365 5859 14399
rect 6561 14365 6595 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 9873 14365 9907 14399
rect 10129 14365 10163 14399
rect 11713 14365 11747 14399
rect 11969 14365 12003 14399
rect 14565 14365 14599 14399
rect 15025 14365 15059 14399
rect 15393 14365 15427 14399
rect 16221 14365 16255 14399
rect 16488 14365 16522 14399
rect 18429 14365 18463 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 20269 14365 20303 14399
rect 21097 14365 21131 14399
rect 23305 14365 23339 14399
rect 25329 14365 25363 14399
rect 26893 14365 26927 14399
rect 3157 14297 3191 14331
rect 9229 14297 9263 14331
rect 21364 14297 21398 14331
rect 26341 14297 26375 14331
rect 26801 14297 26835 14331
rect 1685 14229 1719 14263
rect 6377 14229 6411 14263
rect 7757 14229 7791 14263
rect 9321 14229 9355 14263
rect 11253 14229 11287 14263
rect 13093 14229 13127 14263
rect 18521 14229 18555 14263
rect 23213 14229 23247 14263
rect 23673 14229 23707 14263
rect 1685 14025 1719 14059
rect 2237 14025 2271 14059
rect 3065 14025 3099 14059
rect 3709 14025 3743 14059
rect 6009 14025 6043 14059
rect 9229 14025 9263 14059
rect 12173 14025 12207 14059
rect 18889 14025 18923 14059
rect 21465 14025 21499 14059
rect 27169 14025 27203 14059
rect 7757 13957 7791 13991
rect 17776 13957 17810 13991
rect 22262 13957 22296 13991
rect 2421 13889 2455 13923
rect 2881 13889 2915 13923
rect 3801 13889 3835 13923
rect 4445 13889 4479 13923
rect 5181 13889 5215 13923
rect 5825 13889 5859 13923
rect 6561 13889 6595 13923
rect 7481 13889 7515 13923
rect 10057 13889 10091 13923
rect 10333 13889 10367 13923
rect 10793 13889 10827 13923
rect 11069 13889 11103 13923
rect 11161 13889 11195 13923
rect 12081 13889 12115 13923
rect 12265 13889 12299 13923
rect 12449 13889 12483 13923
rect 13001 13889 13035 13923
rect 15209 13889 15243 13923
rect 15669 13889 15703 13923
rect 16865 13889 16899 13923
rect 17509 13889 17543 13923
rect 19349 13889 19383 13923
rect 19616 13889 19650 13923
rect 21281 13889 21315 13923
rect 24041 13889 24075 13923
rect 4353 13821 4387 13855
rect 5273 13821 5307 13855
rect 9965 13821 9999 13855
rect 14749 13821 14783 13855
rect 15393 13821 15427 13855
rect 15485 13821 15519 13855
rect 15577 13821 15611 13855
rect 22017 13821 22051 13855
rect 24317 13821 24351 13855
rect 24777 13821 24811 13855
rect 26525 13821 26559 13855
rect 11897 13753 11931 13787
rect 6561 13685 6595 13719
rect 15853 13685 15887 13719
rect 16957 13685 16991 13719
rect 20729 13685 20763 13719
rect 23397 13685 23431 13719
rect 25034 13685 25068 13719
rect 9137 13481 9171 13515
rect 11713 13481 11747 13515
rect 12541 13481 12575 13515
rect 16865 13481 16899 13515
rect 18153 13481 18187 13515
rect 21189 13481 21223 13515
rect 23397 13481 23431 13515
rect 24777 13481 24811 13515
rect 27077 13481 27111 13515
rect 13737 13413 13771 13447
rect 4813 13345 4847 13379
rect 6009 13345 6043 13379
rect 6285 13345 6319 13379
rect 10517 13345 10551 13379
rect 11529 13345 11563 13379
rect 12725 13345 12759 13379
rect 14289 13345 14323 13379
rect 14565 13345 14599 13379
rect 20085 13345 20119 13379
rect 20729 13345 20763 13379
rect 22017 13345 22051 13379
rect 25605 13345 25639 13379
rect 1961 13277 1995 13311
rect 2513 13277 2547 13311
rect 3249 13277 3283 13311
rect 4077 13277 4111 13311
rect 4905 13277 4939 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 8309 13277 8343 13311
rect 10250 13277 10284 13311
rect 11069 13277 11103 13311
rect 11989 13277 12023 13311
rect 16773 13277 16807 13311
rect 16865 13277 16899 13311
rect 17417 13277 17451 13311
rect 17601 13277 17635 13311
rect 18061 13277 18095 13311
rect 18245 13277 18279 13311
rect 18705 13277 18739 13311
rect 18889 13277 18923 13311
rect 19809 13277 19843 13311
rect 19901 13277 19935 13311
rect 20821 13277 20855 13311
rect 24041 13277 24075 13311
rect 24593 13277 24627 13311
rect 25329 13277 25363 13311
rect 1869 13209 1903 13243
rect 8585 13209 8619 13243
rect 12909 13209 12943 13243
rect 13185 13209 13219 13243
rect 17509 13209 17543 13243
rect 22284 13209 22318 13243
rect 2513 13141 2547 13175
rect 3433 13141 3467 13175
rect 4261 13141 4295 13175
rect 5549 13141 5583 13175
rect 7757 13141 7791 13175
rect 11897 13141 11931 13175
rect 12817 13141 12851 13175
rect 16037 13141 16071 13175
rect 18705 13141 18739 13175
rect 19441 13141 19475 13175
rect 23857 13141 23891 13175
rect 1685 12937 1719 12971
rect 3985 12937 4019 12971
rect 6561 12937 6595 12971
rect 10333 12937 10367 12971
rect 11897 12937 11931 12971
rect 12909 12937 12943 12971
rect 13737 12937 13771 12971
rect 17233 12937 17267 12971
rect 18245 12937 18279 12971
rect 19533 12937 19567 12971
rect 21281 12937 21315 12971
rect 22017 12937 22051 12971
rect 22477 12937 22511 12971
rect 25421 12937 25455 12971
rect 2513 12869 2547 12903
rect 4874 12869 4908 12903
rect 7849 12869 7883 12903
rect 13829 12869 13863 12903
rect 14105 12869 14139 12903
rect 16313 12869 16347 12903
rect 18521 12869 18555 12903
rect 18613 12869 18647 12903
rect 23305 12869 23339 12903
rect 1777 12801 1811 12835
rect 2237 12801 2271 12835
rect 4629 12801 4663 12835
rect 6929 12801 6963 12835
rect 9597 12801 9631 12835
rect 10333 12801 10367 12835
rect 12817 12801 12851 12835
rect 13553 12801 13587 12835
rect 13921 12801 13955 12835
rect 18424 12801 18458 12835
rect 18741 12801 18775 12835
rect 18889 12801 18923 12835
rect 19349 12801 19383 12835
rect 19993 12801 20027 12835
rect 20177 12801 20211 12835
rect 20637 12801 20671 12835
rect 20821 12801 20855 12835
rect 21465 12801 21499 12835
rect 22385 12801 22419 12835
rect 25421 12801 25455 12835
rect 7021 12733 7055 12767
rect 7205 12733 7239 12767
rect 10149 12733 10183 12767
rect 10701 12733 10735 12767
rect 12265 12733 12299 12767
rect 14565 12733 14599 12767
rect 17325 12733 17359 12767
rect 17417 12733 17451 12767
rect 22661 12733 22695 12767
rect 11713 12665 11747 12699
rect 6009 12597 6043 12631
rect 11897 12597 11931 12631
rect 16865 12597 16899 12631
rect 20085 12597 20119 12631
rect 20729 12597 20763 12631
rect 23765 12597 23799 12631
rect 1961 12393 1995 12427
rect 6561 12393 6595 12427
rect 7021 12393 7055 12427
rect 17233 12393 17267 12427
rect 19809 12393 19843 12427
rect 22845 12393 22879 12427
rect 2605 12257 2639 12291
rect 4629 12257 4663 12291
rect 7481 12257 7515 12291
rect 7665 12257 7699 12291
rect 12173 12257 12207 12291
rect 13369 12257 13403 12291
rect 14749 12257 14783 12291
rect 15301 12257 15335 12291
rect 18613 12257 18647 12291
rect 23121 12257 23155 12291
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 4353 12189 4387 12223
rect 5181 12189 5215 12223
rect 9137 12189 9171 12223
rect 11989 12189 12023 12223
rect 14565 12189 14599 12223
rect 15853 12189 15887 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 20637 12189 20671 12223
rect 21741 12189 21775 12223
rect 23213 12189 23247 12223
rect 1685 12121 1719 12155
rect 3433 12121 3467 12155
rect 5448 12121 5482 12155
rect 7389 12121 7423 12155
rect 8401 12121 8435 12155
rect 8585 12121 8619 12155
rect 9413 12121 9447 12155
rect 12081 12121 12115 12155
rect 16120 12121 16154 12155
rect 18429 12121 18463 12155
rect 23857 12121 23891 12155
rect 3985 12053 4019 12087
rect 4445 12053 4479 12087
rect 8217 12053 8251 12087
rect 10885 12053 10919 12087
rect 11621 12053 11655 12087
rect 12817 12053 12851 12087
rect 13185 12053 13219 12087
rect 13277 12053 13311 12087
rect 18061 12053 18095 12087
rect 18521 12053 18555 12087
rect 20821 12053 20855 12087
rect 21925 12053 21959 12087
rect 2237 11849 2271 11883
rect 4077 11849 4111 11883
rect 10425 11849 10459 11883
rect 13093 11849 13127 11883
rect 14473 11849 14507 11883
rect 15209 11849 15243 11883
rect 16037 11849 16071 11883
rect 18981 11849 19015 11883
rect 19809 11849 19843 11883
rect 20269 11849 20303 11883
rect 2942 11781 2976 11815
rect 8033 11781 8067 11815
rect 8861 11781 8895 11815
rect 14565 11781 14599 11815
rect 17846 11781 17880 11815
rect 19441 11781 19475 11815
rect 22262 11781 22296 11815
rect 2053 11713 2087 11747
rect 4905 11713 4939 11747
rect 5825 11713 5859 11747
rect 6009 11713 6043 11747
rect 6745 11713 6779 11747
rect 7665 11713 7699 11747
rect 7758 11713 7792 11747
rect 7941 11713 7975 11747
rect 8130 11713 8164 11747
rect 9781 11713 9815 11747
rect 10977 11713 11011 11747
rect 11161 11713 11195 11747
rect 11980 11713 12014 11747
rect 13553 11713 13587 11747
rect 13829 11713 13863 11747
rect 15393 11713 15427 11747
rect 16221 11713 16255 11747
rect 16865 11713 16899 11747
rect 19625 11713 19659 11747
rect 24409 11713 24443 11747
rect 2697 11645 2731 11679
rect 4997 11645 5031 11679
rect 5181 11645 5215 11679
rect 6837 11645 6871 11679
rect 7113 11645 7147 11679
rect 9689 11645 9723 11679
rect 11713 11645 11747 11679
rect 13921 11645 13955 11679
rect 17601 11645 17635 11679
rect 22017 11645 22051 11679
rect 5917 11577 5951 11611
rect 11069 11577 11103 11611
rect 21373 11577 21407 11611
rect 4537 11509 4571 11543
rect 8309 11509 8343 11543
rect 17049 11509 17083 11543
rect 20821 11509 20855 11543
rect 23397 11509 23431 11543
rect 24409 11509 24443 11543
rect 3433 11305 3467 11339
rect 7297 11305 7331 11339
rect 9321 11305 9355 11339
rect 17141 11305 17175 11339
rect 17877 11305 17911 11339
rect 18705 11305 18739 11339
rect 19993 11305 20027 11339
rect 21741 11305 21775 11339
rect 22937 11305 22971 11339
rect 23489 11305 23523 11339
rect 26341 11305 26375 11339
rect 4721 11237 4755 11271
rect 6285 11237 6319 11271
rect 7849 11237 7883 11271
rect 9229 11237 9263 11271
rect 16497 11237 16531 11271
rect 4169 11169 4203 11203
rect 8493 11169 8527 11203
rect 12265 11169 12299 11203
rect 20729 11169 20763 11203
rect 22201 11169 22235 11203
rect 22385 11169 22419 11203
rect 24869 11169 24903 11203
rect 2053 11101 2087 11135
rect 4353 11101 4387 11135
rect 5825 11101 5859 11135
rect 6469 11101 6503 11135
rect 7113 11101 7147 11135
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 9137 11101 9171 11135
rect 10057 11101 10091 11135
rect 15781 11101 15815 11135
rect 16037 11101 16071 11135
rect 16681 11101 16715 11135
rect 18061 11101 18095 11135
rect 18613 11101 18647 11135
rect 18797 11101 18831 11135
rect 20821 11101 20855 11135
rect 24593 11101 24627 11135
rect 2298 11033 2332 11067
rect 4261 11033 4295 11067
rect 6929 11033 6963 11067
rect 9413 11033 9447 11067
rect 12532 11033 12566 11067
rect 19533 11033 19567 11067
rect 20913 11033 20947 11067
rect 5641 10965 5675 10999
rect 11345 10965 11379 10999
rect 13645 10965 13679 10999
rect 14657 10965 14691 10999
rect 21281 10965 21315 10999
rect 22109 10965 22143 10999
rect 2145 10761 2179 10795
rect 8309 10761 8343 10795
rect 11897 10761 11931 10795
rect 12357 10761 12391 10795
rect 13921 10761 13955 10795
rect 15853 10761 15887 10795
rect 20453 10761 20487 10795
rect 24961 10761 24995 10795
rect 2872 10693 2906 10727
rect 9597 10693 9631 10727
rect 14473 10693 14507 10727
rect 18337 10693 18371 10727
rect 22262 10693 22296 10727
rect 25421 10693 25455 10727
rect 1961 10625 1995 10659
rect 5181 10625 5215 10659
rect 6745 10625 6779 10659
rect 10425 10625 10459 10659
rect 11713 10625 11747 10659
rect 12541 10625 12575 10659
rect 13185 10625 13219 10659
rect 15393 10625 15427 10659
rect 15485 10625 15519 10659
rect 17325 10625 17359 10659
rect 19533 10625 19567 10659
rect 20269 10625 20303 10659
rect 21097 10625 21131 10659
rect 22017 10625 22051 10659
rect 24133 10625 24167 10659
rect 24593 10625 24627 10659
rect 2605 10557 2639 10591
rect 5089 10557 5123 10591
rect 6653 10557 6687 10591
rect 10149 10557 10183 10591
rect 10333 10557 10367 10591
rect 15301 10557 15335 10591
rect 17509 10557 17543 10591
rect 18429 10557 18463 10591
rect 18521 10557 18555 10591
rect 4537 10489 4571 10523
rect 14657 10489 14691 10523
rect 17969 10489 18003 10523
rect 3985 10421 4019 10455
rect 5549 10421 5583 10455
rect 7113 10421 7147 10455
rect 10793 10421 10827 10455
rect 13001 10421 13035 10455
rect 19349 10421 19383 10455
rect 20913 10421 20947 10455
rect 23397 10421 23431 10455
rect 1685 10217 1719 10251
rect 7389 10217 7423 10251
rect 7849 10217 7883 10251
rect 12725 10217 12759 10251
rect 12909 10217 12943 10251
rect 13737 10217 13771 10251
rect 15117 10217 15151 10251
rect 19441 10217 19475 10251
rect 22569 10217 22603 10251
rect 24777 10217 24811 10251
rect 8585 10149 8619 10183
rect 22109 10149 22143 10183
rect 2881 10081 2915 10115
rect 5457 10081 5491 10115
rect 7481 10081 7515 10115
rect 11989 10081 12023 10115
rect 12265 10081 12299 10115
rect 13001 10081 13035 10115
rect 14841 10081 14875 10115
rect 15761 10081 15795 10115
rect 19993 10081 20027 10115
rect 23121 10081 23155 10115
rect 2697 10013 2731 10047
rect 2973 10013 3007 10047
rect 4537 10013 4571 10047
rect 5181 10013 5215 10047
rect 7665 10013 7699 10047
rect 9597 10013 9631 10047
rect 9873 10013 9907 10047
rect 10793 10013 10827 10047
rect 11897 10013 11931 10047
rect 12909 10013 12943 10047
rect 14749 10013 14783 10047
rect 16773 10013 16807 10047
rect 17417 10013 17451 10047
rect 19809 10013 19843 10047
rect 20729 10013 20763 10047
rect 20996 10013 21030 10047
rect 23765 10013 23799 10047
rect 24593 10013 24627 10047
rect 1961 9945 1995 9979
rect 7389 9945 7423 9979
rect 8401 9945 8435 9979
rect 10701 9945 10735 9979
rect 13185 9945 13219 9979
rect 15945 9945 15979 9979
rect 17662 9945 17696 9979
rect 24041 9945 24075 9979
rect 2513 9877 2547 9911
rect 3985 9877 4019 9911
rect 6929 9877 6963 9911
rect 10241 9877 10275 9911
rect 15853 9877 15887 9911
rect 16313 9877 16347 9911
rect 16957 9877 16991 9911
rect 18797 9877 18831 9911
rect 19901 9877 19935 9911
rect 22937 9877 22971 9911
rect 23029 9877 23063 9911
rect 25329 9877 25363 9911
rect 16313 9673 16347 9707
rect 20545 9673 20579 9707
rect 2320 9605 2354 9639
rect 3985 9605 4019 9639
rect 4169 9605 4203 9639
rect 6561 9605 6595 9639
rect 12817 9605 12851 9639
rect 14473 9605 14507 9639
rect 25237 9605 25271 9639
rect 2053 9537 2087 9571
rect 5273 9537 5307 9571
rect 7021 9537 7055 9571
rect 7389 9537 7423 9571
rect 8309 9537 8343 9571
rect 11713 9537 11747 9571
rect 12725 9537 12759 9571
rect 13737 9537 13771 9571
rect 14933 9537 14967 9571
rect 15200 9537 15234 9571
rect 17233 9537 17267 9571
rect 18245 9537 18279 9571
rect 18521 9537 18555 9571
rect 19432 9537 19466 9571
rect 21189 9537 21223 9571
rect 22385 9537 22419 9571
rect 23213 9537 23247 9571
rect 5181 9469 5215 9503
rect 8401 9469 8435 9503
rect 8861 9469 8895 9503
rect 9137 9469 9171 9503
rect 12909 9469 12943 9503
rect 17325 9469 17359 9503
rect 17417 9469 17451 9503
rect 18337 9469 18371 9503
rect 19165 9469 19199 9503
rect 22293 9469 22327 9503
rect 25513 9469 25547 9503
rect 5641 9401 5675 9435
rect 12357 9401 12391 9435
rect 16865 9401 16899 9435
rect 3433 9333 3467 9367
rect 10609 9333 10643 9367
rect 11897 9333 11931 9367
rect 13553 9333 13587 9367
rect 18521 9333 18555 9367
rect 18705 9333 18739 9367
rect 21005 9333 21039 9367
rect 22017 9333 22051 9367
rect 23305 9333 23339 9367
rect 23765 9333 23799 9367
rect 5089 9129 5123 9163
rect 8033 9129 8067 9163
rect 9137 9129 9171 9163
rect 11621 9129 11655 9163
rect 16589 9129 16623 9163
rect 17601 9129 17635 9163
rect 18429 9129 18463 9163
rect 18889 9129 18923 9163
rect 22845 9129 22879 9163
rect 3249 9061 3283 9095
rect 23857 9061 23891 9095
rect 1869 8993 1903 9027
rect 3985 8993 4019 9027
rect 8493 8993 8527 9027
rect 11345 8993 11379 9027
rect 15209 8993 15243 9027
rect 17141 8993 17175 9027
rect 20821 8993 20855 9027
rect 23121 8993 23155 9027
rect 24685 8993 24719 9027
rect 4169 8925 4203 8959
rect 5089 8925 5123 8959
rect 5549 8925 5583 8959
rect 8401 8925 8435 8959
rect 10517 8925 10551 8959
rect 11253 8925 11287 8959
rect 12081 8925 12115 8959
rect 12337 8925 12371 8959
rect 14565 8925 14599 8959
rect 17233 8925 17267 8959
rect 18613 8925 18647 8959
rect 18705 8925 18739 8959
rect 18889 8925 18923 8959
rect 20565 8925 20599 8959
rect 21557 8925 21591 8959
rect 22017 8925 22051 8959
rect 23213 8925 23247 8959
rect 25145 8925 25179 8959
rect 25329 8925 25363 8959
rect 26157 8925 26191 8959
rect 2136 8857 2170 8891
rect 5825 8857 5859 8891
rect 10272 8857 10306 8891
rect 15454 8857 15488 8891
rect 4353 8789 4387 8823
rect 7297 8789 7331 8823
rect 13461 8789 13495 8823
rect 14749 8789 14783 8823
rect 19441 8789 19475 8823
rect 22385 8789 22419 8823
rect 2697 8585 2731 8619
rect 3709 8585 3743 8619
rect 5641 8585 5675 8619
rect 6561 8585 6595 8619
rect 10977 8585 11011 8619
rect 12541 8585 12575 8619
rect 15945 8585 15979 8619
rect 19257 8585 19291 8619
rect 25053 8585 25087 8619
rect 25697 8585 25731 8619
rect 1961 8517 1995 8551
rect 13001 8517 13035 8551
rect 14749 8517 14783 8551
rect 16957 8517 16991 8551
rect 19717 8517 19751 8551
rect 23581 8517 23615 8551
rect 2145 8449 2179 8483
rect 2237 8449 2271 8483
rect 2881 8449 2915 8483
rect 3157 8449 3191 8483
rect 3893 8449 3927 8483
rect 5089 8449 5123 8483
rect 5825 8449 5859 8483
rect 7021 8449 7055 8483
rect 7205 8449 7239 8483
rect 8125 8449 8159 8483
rect 8309 8449 8343 8483
rect 11161 8449 11195 8483
rect 11989 8449 12023 8483
rect 15393 8449 15427 8483
rect 16129 8449 16163 8483
rect 17877 8449 17911 8483
rect 18061 8449 18095 8483
rect 18889 8449 18923 8483
rect 22385 8449 22419 8483
rect 25513 8449 25547 8483
rect 10241 8381 10275 8415
rect 10517 8381 10551 8415
rect 11713 8381 11747 8415
rect 18613 8381 18647 8415
rect 18797 8381 18831 8415
rect 22293 8381 22327 8415
rect 23305 8381 23339 8415
rect 1961 8313 1995 8347
rect 3065 8313 3099 8347
rect 5089 8313 5123 8347
rect 8125 8313 8159 8347
rect 8769 8313 8803 8347
rect 22017 8313 22051 8347
rect 15301 8245 15335 8279
rect 17969 8245 18003 8279
rect 21005 8245 21039 8279
rect 2053 8041 2087 8075
rect 6009 8041 6043 8075
rect 8033 8041 8067 8075
rect 9137 8041 9171 8075
rect 9873 8041 9907 8075
rect 13369 8041 13403 8075
rect 14289 8041 14323 8075
rect 18521 8041 18555 8075
rect 19533 8041 19567 8075
rect 22109 8041 22143 8075
rect 23029 8041 23063 8075
rect 26157 8041 26191 8075
rect 12173 7905 12207 7939
rect 12725 7905 12759 7939
rect 14565 7905 14599 7939
rect 23305 7905 23339 7939
rect 24685 7905 24719 7939
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 5273 7837 5307 7871
rect 6193 7837 6227 7871
rect 9689 7837 9723 7871
rect 10425 7837 10459 7871
rect 14657 7837 14691 7871
rect 15761 7837 15795 7871
rect 16957 7837 16991 7871
rect 17325 7837 17359 7871
rect 17969 7837 18003 7871
rect 18245 7837 18279 7871
rect 18337 7837 18371 7871
rect 20361 7837 20395 7871
rect 23397 7837 23431 7871
rect 25145 7837 25179 7871
rect 25421 7837 25455 7871
rect 3341 7769 3375 7803
rect 4353 7769 4387 7803
rect 6745 7769 6779 7803
rect 13001 7769 13035 7803
rect 17141 7769 17175 7803
rect 18153 7769 18187 7803
rect 20821 7769 20855 7803
rect 5365 7701 5399 7735
rect 12909 7701 12943 7735
rect 15761 7701 15795 7735
rect 16497 7701 16531 7735
rect 20177 7701 20211 7735
rect 3893 7497 3927 7531
rect 13553 7497 13587 7531
rect 14105 7497 14139 7531
rect 17141 7497 17175 7531
rect 18429 7497 18463 7531
rect 22661 7497 22695 7531
rect 24961 7497 24995 7531
rect 10333 7429 10367 7463
rect 14841 7429 14875 7463
rect 18797 7429 18831 7463
rect 24133 7429 24167 7463
rect 25881 7429 25915 7463
rect 1869 7361 1903 7395
rect 2605 7361 2639 7395
rect 5089 7361 5123 7395
rect 5733 7361 5767 7395
rect 7021 7361 7055 7395
rect 7389 7361 7423 7395
rect 10885 7361 10919 7395
rect 12173 7361 12207 7395
rect 12440 7361 12474 7395
rect 16957 7361 16991 7395
rect 17141 7361 17175 7395
rect 18613 7361 18647 7395
rect 19441 7361 19475 7395
rect 19625 7361 19659 7395
rect 21189 7361 21223 7395
rect 24961 7361 24995 7395
rect 25605 7361 25639 7395
rect 4813 7293 4847 7327
rect 6561 7293 6595 7327
rect 14565 7293 14599 7327
rect 17969 7293 18003 7327
rect 20453 7293 20487 7327
rect 24409 7293 24443 7327
rect 2053 7225 2087 7259
rect 5917 7225 5951 7259
rect 4905 7157 4939 7191
rect 5273 7157 5307 7191
rect 9045 7157 9079 7191
rect 10977 7157 11011 7191
rect 16313 7157 16347 7191
rect 21005 7157 21039 7191
rect 4169 6953 4203 6987
rect 6849 6953 6883 6987
rect 9584 6953 9618 6987
rect 14381 6953 14415 6987
rect 21170 6953 21204 6987
rect 3433 6885 3467 6919
rect 8217 6817 8251 6851
rect 11713 6817 11747 6851
rect 13093 6817 13127 6851
rect 13369 6817 13403 6851
rect 15117 6817 15151 6851
rect 17049 6817 17083 6851
rect 20913 6817 20947 6851
rect 22661 6817 22695 6851
rect 23397 6817 23431 6851
rect 2053 6749 2087 6783
rect 2320 6749 2354 6783
rect 7113 6749 7147 6783
rect 7573 6749 7607 6783
rect 9321 6749 9355 6783
rect 11989 6749 12023 6783
rect 13461 6749 13495 6783
rect 14841 6749 14875 6783
rect 17233 6749 17267 6783
rect 18061 6749 18095 6783
rect 18797 6749 18831 6783
rect 19717 6749 19751 6783
rect 20453 6749 20487 6783
rect 23121 6749 23155 6783
rect 3985 6681 4019 6715
rect 4185 6613 4219 6647
rect 4353 6613 4387 6647
rect 4813 6613 4847 6647
rect 5365 6613 5399 6647
rect 11069 6613 11103 6647
rect 12633 6613 12667 6647
rect 16589 6613 16623 6647
rect 17877 6613 17911 6647
rect 18797 6613 18831 6647
rect 19533 6613 19567 6647
rect 20269 6613 20303 6647
rect 3433 6409 3467 6443
rect 8769 6409 8803 6443
rect 9321 6409 9355 6443
rect 13461 6409 13495 6443
rect 15945 6409 15979 6443
rect 20821 6409 20855 6443
rect 22845 6409 22879 6443
rect 10885 6341 10919 6375
rect 17141 6341 17175 6375
rect 19349 6341 19383 6375
rect 2053 6273 2087 6307
rect 2320 6273 2354 6307
rect 3985 6273 4019 6307
rect 4077 6273 4111 6307
rect 5365 6273 5399 6307
rect 7021 6273 7055 6307
rect 10149 6273 10183 6307
rect 11161 6273 11195 6307
rect 11713 6273 11747 6307
rect 14013 6273 14047 6307
rect 15301 6273 15335 6307
rect 15577 6273 15611 6307
rect 23489 6273 23523 6307
rect 23857 6273 23891 6307
rect 5457 6205 5491 6239
rect 6009 6205 6043 6239
rect 7297 6205 7331 6239
rect 10241 6205 10275 6239
rect 11989 6205 12023 6239
rect 16865 6205 16899 6239
rect 19073 6205 19107 6239
rect 4261 6069 4295 6103
rect 14013 6069 14047 6103
rect 18613 6069 18647 6103
rect 22293 6069 22327 6103
rect 2421 5865 2455 5899
rect 2973 5865 3007 5899
rect 4813 5865 4847 5899
rect 7389 5865 7423 5899
rect 8033 5865 8067 5899
rect 11332 5865 11366 5899
rect 18429 5865 18463 5899
rect 21189 5865 21223 5899
rect 3985 5797 4019 5831
rect 12817 5797 12851 5831
rect 13737 5797 13771 5831
rect 3433 5729 3467 5763
rect 5917 5729 5951 5763
rect 10609 5729 10643 5763
rect 11069 5729 11103 5763
rect 14565 5729 14599 5763
rect 16129 5729 16163 5763
rect 17693 5729 17727 5763
rect 19441 5729 19475 5763
rect 19717 5729 19751 5763
rect 1593 5661 1627 5695
rect 1777 5661 1811 5695
rect 2237 5661 2271 5695
rect 3157 5661 3191 5695
rect 3341 5661 3375 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 4813 5661 4847 5695
rect 4997 5661 5031 5695
rect 5641 5661 5675 5695
rect 8125 5661 8159 5695
rect 9965 5661 9999 5695
rect 10241 5661 10275 5695
rect 13737 5661 13771 5695
rect 15301 5661 15335 5695
rect 15761 5661 15795 5695
rect 16957 5661 16991 5695
rect 17417 5661 17451 5695
rect 18429 5661 18463 5695
rect 1685 5593 1719 5627
rect 4169 5525 4203 5559
rect 2053 5321 2087 5355
rect 5825 5321 5859 5355
rect 6653 5321 6687 5355
rect 8309 5321 8343 5355
rect 11161 5321 11195 5355
rect 12541 5321 12575 5355
rect 14933 5321 14967 5355
rect 18705 5321 18739 5355
rect 4721 5253 4755 5287
rect 9137 5253 9171 5287
rect 11989 5253 12023 5287
rect 16865 5253 16899 5287
rect 19993 5253 20027 5287
rect 1961 5185 1995 5219
rect 2145 5185 2179 5219
rect 2872 5185 2906 5219
rect 4445 5185 4479 5219
rect 5641 5185 5675 5219
rect 6745 5185 6779 5219
rect 7665 5185 7699 5219
rect 8861 5185 8895 5219
rect 10333 5185 10367 5219
rect 10793 5185 10827 5219
rect 11713 5185 11747 5219
rect 12449 5185 12483 5219
rect 17141 5185 17175 5219
rect 2605 5117 2639 5151
rect 7389 5117 7423 5151
rect 4537 5049 4571 5083
rect 3985 4981 4019 5015
rect 4445 4981 4479 5015
rect 3985 4777 4019 4811
rect 5549 4777 5583 4811
rect 9137 4777 9171 4811
rect 11713 4777 11747 4811
rect 2421 4709 2455 4743
rect 4537 4709 4571 4743
rect 3341 4641 3375 4675
rect 8217 4641 8251 4675
rect 2237 4573 2271 4607
rect 2513 4573 2547 4607
rect 3157 4573 3191 4607
rect 3433 4573 3467 4607
rect 4169 4573 4203 4607
rect 4261 4573 4295 4607
rect 7573 4573 7607 4607
rect 10425 4573 10459 4607
rect 7021 4505 7055 4539
rect 2053 4437 2087 4471
rect 2973 4437 3007 4471
rect 4353 4437 4387 4471
rect 9873 4437 9907 4471
rect 4261 4233 4295 4267
rect 4997 4233 5031 4267
rect 3126 4165 3160 4199
rect 5165 4165 5199 4199
rect 5365 4165 5399 4199
rect 1593 4097 1627 4131
rect 2237 4097 2271 4131
rect 2421 4097 2455 4131
rect 7113 4097 7147 4131
rect 7573 4097 7607 4131
rect 8953 4097 8987 4131
rect 18981 4097 19015 4131
rect 19625 4097 19659 4131
rect 2881 4029 2915 4063
rect 18889 4029 18923 4063
rect 5917 3961 5951 3995
rect 1777 3893 1811 3927
rect 2237 3893 2271 3927
rect 5181 3893 5215 3927
rect 8125 3893 8159 3927
rect 3433 3689 3467 3723
rect 4261 3689 4295 3723
rect 4813 3689 4847 3723
rect 5365 3689 5399 3723
rect 5917 3689 5951 3723
rect 6469 3689 6503 3723
rect 2053 3485 2087 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4261 3485 4295 3519
rect 7021 3485 7055 3519
rect 7941 3485 7975 3519
rect 2320 3417 2354 3451
rect 2053 3145 2087 3179
rect 5181 3145 5215 3179
rect 5733 3145 5767 3179
rect 3341 3077 3375 3111
rect 4068 3077 4102 3111
rect 6561 3009 6595 3043
rect 3801 2941 3835 2975
rect 1593 2601 1627 2635
rect 2237 2601 2271 2635
rect 3985 2601 4019 2635
rect 5181 2601 5215 2635
rect 5733 2601 5767 2635
rect 4537 2533 4571 2567
rect 2789 2465 2823 2499
rect 3249 2261 3283 2295
<< metal1 >>
rect 1104 26682 27876 26704
rect 1104 26630 4296 26682
rect 4348 26630 4360 26682
rect 4412 26630 4424 26682
rect 4476 26630 4488 26682
rect 4540 26630 4552 26682
rect 4604 26630 10988 26682
rect 11040 26630 11052 26682
rect 11104 26630 11116 26682
rect 11168 26630 11180 26682
rect 11232 26630 11244 26682
rect 11296 26630 17680 26682
rect 17732 26630 17744 26682
rect 17796 26630 17808 26682
rect 17860 26630 17872 26682
rect 17924 26630 17936 26682
rect 17988 26630 24372 26682
rect 24424 26630 24436 26682
rect 24488 26630 24500 26682
rect 24552 26630 24564 26682
rect 24616 26630 24628 26682
rect 24680 26630 27876 26682
rect 1104 26608 27876 26630
rect 1854 26528 1860 26580
rect 1912 26568 1918 26580
rect 2593 26571 2651 26577
rect 2593 26568 2605 26571
rect 1912 26540 2605 26568
rect 1912 26528 1918 26540
rect 2593 26537 2605 26540
rect 2639 26537 2651 26571
rect 2593 26531 2651 26537
rect 5169 26571 5227 26577
rect 5169 26537 5181 26571
rect 5215 26568 5227 26571
rect 5442 26568 5448 26580
rect 5215 26540 5448 26568
rect 5215 26537 5227 26540
rect 5169 26531 5227 26537
rect 5442 26528 5448 26540
rect 5500 26528 5506 26580
rect 9030 26528 9036 26580
rect 9088 26568 9094 26580
rect 9309 26571 9367 26577
rect 9309 26568 9321 26571
rect 9088 26540 9321 26568
rect 9088 26528 9094 26540
rect 9309 26537 9321 26540
rect 9355 26537 9367 26571
rect 9309 26531 9367 26537
rect 19794 26528 19800 26580
rect 19852 26568 19858 26580
rect 20349 26571 20407 26577
rect 20349 26568 20361 26571
rect 19852 26540 20361 26568
rect 19852 26528 19858 26540
rect 20349 26537 20361 26540
rect 20395 26537 20407 26571
rect 20349 26531 20407 26537
rect 23474 26528 23480 26580
rect 23532 26568 23538 26580
rect 23661 26571 23719 26577
rect 23661 26568 23673 26571
rect 23532 26540 23673 26568
rect 23532 26528 23538 26540
rect 23661 26537 23673 26540
rect 23707 26537 23719 26571
rect 23661 26531 23719 26537
rect 26513 26571 26571 26577
rect 26513 26537 26525 26571
rect 26559 26568 26571 26571
rect 26970 26568 26976 26580
rect 26559 26540 26976 26568
rect 26559 26537 26571 26540
rect 26513 26531 26571 26537
rect 26970 26528 26976 26540
rect 27028 26528 27034 26580
rect 5718 26392 5724 26444
rect 5776 26432 5782 26444
rect 15286 26432 15292 26444
rect 5776 26404 5856 26432
rect 15247 26404 15292 26432
rect 5776 26392 5782 26404
rect 1670 26364 1676 26376
rect 1631 26336 1676 26364
rect 1670 26324 1676 26336
rect 1728 26324 1734 26376
rect 2777 26367 2835 26373
rect 2777 26333 2789 26367
rect 2823 26364 2835 26367
rect 4522 26364 4528 26376
rect 2823 26336 4528 26364
rect 2823 26333 2835 26336
rect 2777 26327 2835 26333
rect 4522 26324 4528 26336
rect 4580 26324 4586 26376
rect 4982 26364 4988 26376
rect 4943 26336 4988 26364
rect 4982 26324 4988 26336
rect 5040 26324 5046 26376
rect 5828 26373 5856 26404
rect 15286 26392 15292 26404
rect 15344 26392 15350 26444
rect 15752 26376 15804 26382
rect 5813 26367 5871 26373
rect 5813 26333 5825 26367
rect 5859 26333 5871 26367
rect 6546 26364 6552 26376
rect 6507 26336 6552 26364
rect 5813 26327 5871 26333
rect 6546 26324 6552 26336
rect 6604 26324 6610 26376
rect 6733 26367 6791 26373
rect 6733 26333 6745 26367
rect 6779 26333 6791 26367
rect 9122 26364 9128 26376
rect 9083 26336 9128 26364
rect 6733 26327 6791 26333
rect 2041 26299 2099 26305
rect 2041 26265 2053 26299
rect 2087 26296 2099 26299
rect 5074 26296 5080 26308
rect 2087 26268 5080 26296
rect 2087 26265 2099 26268
rect 2041 26259 2099 26265
rect 5074 26256 5080 26268
rect 5132 26256 5138 26308
rect 5350 26256 5356 26308
rect 5408 26296 5414 26308
rect 5721 26299 5779 26305
rect 5721 26296 5733 26299
rect 5408 26268 5733 26296
rect 5408 26256 5414 26268
rect 5721 26265 5733 26268
rect 5767 26265 5779 26299
rect 5721 26259 5779 26265
rect 6362 26256 6368 26308
rect 6420 26296 6426 26308
rect 6748 26296 6776 26327
rect 9122 26324 9128 26336
rect 9180 26324 9186 26376
rect 9398 26324 9404 26376
rect 9456 26364 9462 26376
rect 9861 26367 9919 26373
rect 9861 26364 9873 26367
rect 9456 26336 9873 26364
rect 9456 26324 9462 26336
rect 9861 26333 9873 26336
rect 9907 26333 9919 26367
rect 9861 26327 9919 26333
rect 10045 26367 10103 26373
rect 10045 26333 10057 26367
rect 10091 26333 10103 26367
rect 10045 26327 10103 26333
rect 11793 26367 11851 26373
rect 11793 26333 11805 26367
rect 11839 26364 11851 26367
rect 12345 26367 12403 26373
rect 12345 26364 12357 26367
rect 11839 26336 12357 26364
rect 11839 26333 11851 26336
rect 11793 26327 11851 26333
rect 12345 26333 12357 26336
rect 12391 26333 12403 26367
rect 13630 26364 13636 26376
rect 13018 26336 13636 26364
rect 12345 26327 12403 26333
rect 6420 26268 6776 26296
rect 6420 26256 6426 26268
rect 9490 26256 9496 26308
rect 9548 26296 9554 26308
rect 10060 26296 10088 26327
rect 9548 26268 10088 26296
rect 12360 26296 12388 26327
rect 13630 26324 13636 26336
rect 13688 26324 13694 26376
rect 13814 26324 13820 26376
rect 13872 26364 13878 26376
rect 14277 26367 14335 26373
rect 14277 26364 14289 26367
rect 13872 26336 14289 26364
rect 13872 26324 13878 26336
rect 14277 26333 14289 26336
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 16850 26364 16856 26376
rect 16811 26336 16856 26364
rect 16850 26324 16856 26336
rect 16908 26324 16914 26376
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19521 26367 19579 26373
rect 19521 26364 19533 26367
rect 19392 26336 19533 26364
rect 19392 26324 19398 26336
rect 19521 26333 19533 26336
rect 19567 26333 19579 26367
rect 20162 26364 20168 26376
rect 20123 26336 20168 26364
rect 19521 26327 19579 26333
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 23474 26364 23480 26376
rect 23435 26336 23480 26364
rect 23474 26324 23480 26336
rect 23532 26324 23538 26376
rect 26326 26364 26332 26376
rect 26287 26336 26332 26364
rect 26326 26324 26332 26336
rect 26384 26324 26390 26376
rect 15752 26318 15804 26324
rect 12526 26296 12532 26308
rect 12360 26268 12532 26296
rect 9548 26256 9554 26268
rect 12526 26256 12532 26268
rect 12584 26256 12590 26308
rect 13262 26256 13268 26308
rect 13320 26296 13326 26308
rect 13357 26299 13415 26305
rect 13357 26296 13369 26299
rect 13320 26268 13369 26296
rect 13320 26256 13326 26268
rect 13357 26265 13369 26268
rect 13403 26265 13415 26299
rect 16114 26296 16120 26308
rect 16075 26268 16120 26296
rect 13357 26259 13415 26265
rect 16114 26256 16120 26268
rect 16172 26256 16178 26308
rect 19426 26296 19432 26308
rect 19387 26268 19432 26296
rect 19426 26256 19432 26268
rect 19484 26256 19490 26308
rect 5902 26188 5908 26240
rect 5960 26228 5966 26240
rect 6549 26231 6607 26237
rect 6549 26228 6561 26231
rect 5960 26200 6561 26228
rect 5960 26188 5966 26200
rect 6549 26197 6561 26200
rect 6595 26197 6607 26231
rect 6549 26191 6607 26197
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 9953 26231 10011 26237
rect 9953 26228 9965 26231
rect 9916 26200 9965 26228
rect 9916 26188 9922 26200
rect 9953 26197 9965 26200
rect 9999 26197 10011 26231
rect 9953 26191 10011 26197
rect 12618 26188 12624 26240
rect 12676 26228 12682 26240
rect 14461 26231 14519 26237
rect 14461 26228 14473 26231
rect 12676 26200 14473 26228
rect 12676 26188 12682 26200
rect 14461 26197 14473 26200
rect 14507 26197 14519 26231
rect 14461 26191 14519 26197
rect 16206 26188 16212 26240
rect 16264 26228 16270 26240
rect 17037 26231 17095 26237
rect 17037 26228 17049 26231
rect 16264 26200 17049 26228
rect 16264 26188 16270 26200
rect 17037 26197 17049 26200
rect 17083 26197 17095 26231
rect 17037 26191 17095 26197
rect 1104 26138 28032 26160
rect 1104 26086 7642 26138
rect 7694 26086 7706 26138
rect 7758 26086 7770 26138
rect 7822 26086 7834 26138
rect 7886 26086 7898 26138
rect 7950 26086 14334 26138
rect 14386 26086 14398 26138
rect 14450 26086 14462 26138
rect 14514 26086 14526 26138
rect 14578 26086 14590 26138
rect 14642 26086 21026 26138
rect 21078 26086 21090 26138
rect 21142 26086 21154 26138
rect 21206 26086 21218 26138
rect 21270 26086 21282 26138
rect 21334 26086 27718 26138
rect 27770 26086 27782 26138
rect 27834 26086 27846 26138
rect 27898 26086 27910 26138
rect 27962 26086 27974 26138
rect 28026 26086 28032 26138
rect 1104 26064 28032 26086
rect 1670 26024 1676 26036
rect 1631 25996 1676 26024
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 4522 26024 4528 26036
rect 4483 25996 4528 26024
rect 4522 25984 4528 25996
rect 4580 25984 4586 26036
rect 4982 25984 4988 26036
rect 5040 26024 5046 26036
rect 5077 26027 5135 26033
rect 5077 26024 5089 26027
rect 5040 25996 5089 26024
rect 5040 25984 5046 25996
rect 5077 25993 5089 25996
rect 5123 25993 5135 26027
rect 5077 25987 5135 25993
rect 8665 26027 8723 26033
rect 8665 25993 8677 26027
rect 8711 26024 8723 26027
rect 9122 26024 9128 26036
rect 8711 25996 9128 26024
rect 8711 25993 8723 25996
rect 8665 25987 8723 25993
rect 9122 25984 9128 25996
rect 9180 25984 9186 26036
rect 10137 26027 10195 26033
rect 10137 25993 10149 26027
rect 10183 25993 10195 26027
rect 10137 25987 10195 25993
rect 10152 25956 10180 25987
rect 13814 25956 13820 25968
rect 10152 25928 13820 25956
rect 13814 25916 13820 25928
rect 13872 25916 13878 25968
rect 14090 25916 14096 25968
rect 14148 25916 14154 25968
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 2958 25888 2964 25900
rect 2639 25860 2964 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 4433 25891 4491 25897
rect 4433 25857 4445 25891
rect 4479 25857 4491 25891
rect 4433 25851 4491 25857
rect 4617 25891 4675 25897
rect 4617 25857 4629 25891
rect 4663 25888 4675 25891
rect 5442 25888 5448 25900
rect 4663 25860 5448 25888
rect 4663 25857 4675 25860
rect 4617 25851 4675 25857
rect 2498 25820 2504 25832
rect 2459 25792 2504 25820
rect 2498 25780 2504 25792
rect 2556 25780 2562 25832
rect 4448 25820 4476 25851
rect 5442 25848 5448 25860
rect 5500 25848 5506 25900
rect 6730 25888 6736 25900
rect 6691 25860 6736 25888
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25857 8355 25891
rect 9766 25888 9772 25900
rect 9727 25860 9772 25888
rect 8297 25851 8355 25857
rect 4798 25820 4804 25832
rect 4448 25792 4804 25820
rect 4798 25780 4804 25792
rect 4856 25780 4862 25832
rect 5353 25823 5411 25829
rect 5353 25789 5365 25823
rect 5399 25820 5411 25823
rect 5902 25820 5908 25832
rect 5399 25792 5908 25820
rect 5399 25789 5411 25792
rect 5353 25783 5411 25789
rect 5902 25780 5908 25792
rect 5960 25780 5966 25832
rect 7374 25780 7380 25832
rect 7432 25820 7438 25832
rect 8205 25823 8263 25829
rect 8205 25820 8217 25823
rect 7432 25792 8217 25820
rect 7432 25780 7438 25792
rect 8205 25789 8217 25792
rect 8251 25789 8263 25823
rect 8205 25783 8263 25789
rect 2222 25684 2228 25696
rect 2183 25656 2228 25684
rect 2222 25644 2228 25656
rect 2280 25644 2286 25696
rect 6733 25687 6791 25693
rect 6733 25653 6745 25687
rect 6779 25684 6791 25687
rect 7006 25684 7012 25696
rect 6779 25656 7012 25684
rect 6779 25653 6791 25656
rect 6733 25647 6791 25653
rect 7006 25644 7012 25656
rect 7064 25644 7070 25696
rect 7098 25644 7104 25696
rect 7156 25684 7162 25696
rect 8312 25684 8340 25851
rect 9766 25848 9772 25860
rect 9824 25848 9830 25900
rect 10778 25888 10784 25900
rect 10739 25860 10784 25888
rect 10778 25848 10784 25860
rect 10836 25848 10842 25900
rect 12066 25888 12072 25900
rect 12027 25860 12072 25888
rect 12066 25848 12072 25860
rect 12124 25848 12130 25900
rect 12710 25888 12716 25900
rect 12671 25860 12716 25888
rect 12710 25848 12716 25860
rect 12768 25848 12774 25900
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 15028 25860 15485 25888
rect 15028 25832 15056 25860
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25888 17187 25891
rect 17310 25888 17316 25900
rect 17175 25860 17316 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17310 25848 17316 25860
rect 17368 25848 17374 25900
rect 18785 25891 18843 25897
rect 18785 25857 18797 25891
rect 18831 25888 18843 25891
rect 19334 25888 19340 25900
rect 18831 25860 19340 25888
rect 18831 25857 18843 25860
rect 18785 25851 18843 25857
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 19886 25848 19892 25900
rect 19944 25848 19950 25900
rect 9858 25820 9864 25832
rect 9819 25792 9864 25820
rect 9858 25780 9864 25792
rect 9916 25780 9922 25832
rect 10686 25820 10692 25832
rect 10647 25792 10692 25820
rect 10686 25780 10692 25792
rect 10744 25780 10750 25832
rect 12805 25823 12863 25829
rect 12805 25789 12817 25823
rect 12851 25820 12863 25823
rect 13265 25823 13323 25829
rect 13265 25820 13277 25823
rect 12851 25792 13277 25820
rect 12851 25789 12863 25792
rect 12805 25783 12863 25789
rect 13265 25789 13277 25792
rect 13311 25789 13323 25823
rect 13265 25783 13323 25789
rect 13541 25823 13599 25829
rect 13541 25789 13553 25823
rect 13587 25820 13599 25823
rect 14182 25820 14188 25832
rect 13587 25792 14188 25820
rect 13587 25789 13599 25792
rect 13541 25783 13599 25789
rect 14182 25780 14188 25792
rect 14240 25780 14246 25832
rect 15010 25820 15016 25832
rect 14923 25792 15016 25820
rect 15010 25780 15016 25792
rect 15068 25780 15074 25832
rect 15286 25780 15292 25832
rect 15344 25820 15350 25832
rect 16209 25823 16267 25829
rect 16209 25820 16221 25823
rect 15344 25792 16221 25820
rect 15344 25780 15350 25792
rect 16209 25789 16221 25792
rect 16255 25789 16267 25823
rect 16209 25783 16267 25789
rect 19797 25823 19855 25829
rect 19797 25789 19809 25823
rect 19843 25820 19855 25823
rect 20070 25820 20076 25832
rect 19843 25792 20076 25820
rect 19843 25789 19855 25792
rect 19797 25783 19855 25789
rect 20070 25780 20076 25792
rect 20128 25780 20134 25832
rect 20625 25823 20683 25829
rect 20625 25789 20637 25823
rect 20671 25820 20683 25823
rect 20806 25820 20812 25832
rect 20671 25792 20812 25820
rect 20671 25789 20683 25792
rect 20625 25783 20683 25789
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 11149 25755 11207 25761
rect 11149 25721 11161 25755
rect 11195 25752 11207 25755
rect 16850 25752 16856 25764
rect 11195 25724 12434 25752
rect 11195 25721 11207 25724
rect 11149 25715 11207 25721
rect 11330 25684 11336 25696
rect 7156 25656 11336 25684
rect 7156 25644 7162 25656
rect 11330 25644 11336 25656
rect 11388 25644 11394 25696
rect 11882 25684 11888 25696
rect 11843 25656 11888 25684
rect 11882 25644 11888 25656
rect 11940 25644 11946 25696
rect 12406 25684 12434 25724
rect 14568 25724 16856 25752
rect 14568 25684 14596 25724
rect 16850 25712 16856 25724
rect 16908 25712 16914 25764
rect 15470 25684 15476 25696
rect 12406 25656 14596 25684
rect 15431 25656 15476 25684
rect 15470 25644 15476 25656
rect 15528 25644 15534 25696
rect 17126 25684 17132 25696
rect 17087 25656 17132 25684
rect 17126 25644 17132 25656
rect 17184 25644 17190 25696
rect 18598 25684 18604 25696
rect 18559 25656 18604 25684
rect 18598 25644 18604 25656
rect 18656 25644 18662 25696
rect 1104 25594 27876 25616
rect 1104 25542 4296 25594
rect 4348 25542 4360 25594
rect 4412 25542 4424 25594
rect 4476 25542 4488 25594
rect 4540 25542 4552 25594
rect 4604 25542 10988 25594
rect 11040 25542 11052 25594
rect 11104 25542 11116 25594
rect 11168 25542 11180 25594
rect 11232 25542 11244 25594
rect 11296 25542 17680 25594
rect 17732 25542 17744 25594
rect 17796 25542 17808 25594
rect 17860 25542 17872 25594
rect 17924 25542 17936 25594
rect 17988 25542 24372 25594
rect 24424 25542 24436 25594
rect 24488 25542 24500 25594
rect 24552 25542 24564 25594
rect 24616 25542 24628 25594
rect 24680 25542 27876 25594
rect 1104 25520 27876 25542
rect 4798 25480 4804 25492
rect 4759 25452 4804 25480
rect 4798 25440 4804 25452
rect 4856 25440 4862 25492
rect 5276 25452 5488 25480
rect 3421 25415 3479 25421
rect 3421 25381 3433 25415
rect 3467 25412 3479 25415
rect 4154 25412 4160 25424
rect 3467 25384 4160 25412
rect 3467 25381 3479 25384
rect 3421 25375 3479 25381
rect 4154 25372 4160 25384
rect 4212 25372 4218 25424
rect 4341 25415 4399 25421
rect 4341 25381 4353 25415
rect 4387 25412 4399 25415
rect 5276 25412 5304 25452
rect 4387 25384 5304 25412
rect 5460 25412 5488 25452
rect 12710 25440 12716 25492
rect 12768 25480 12774 25492
rect 13633 25483 13691 25489
rect 13633 25480 13645 25483
rect 12768 25452 13645 25480
rect 12768 25440 12774 25452
rect 13633 25449 13645 25452
rect 13679 25449 13691 25483
rect 20162 25480 20168 25492
rect 13633 25443 13691 25449
rect 16132 25452 20168 25480
rect 5534 25412 5540 25424
rect 5460 25384 5540 25412
rect 4387 25381 4399 25384
rect 4341 25375 4399 25381
rect 5534 25372 5540 25384
rect 5592 25372 5598 25424
rect 5721 25415 5779 25421
rect 5721 25381 5733 25415
rect 5767 25412 5779 25415
rect 7374 25412 7380 25424
rect 5767 25384 7380 25412
rect 5767 25381 5779 25384
rect 5721 25375 5779 25381
rect 7374 25372 7380 25384
rect 7432 25372 7438 25424
rect 7469 25415 7527 25421
rect 7469 25381 7481 25415
rect 7515 25412 7527 25415
rect 9398 25412 9404 25424
rect 7515 25384 9404 25412
rect 7515 25381 7527 25384
rect 7469 25375 7527 25381
rect 9398 25372 9404 25384
rect 9456 25372 9462 25424
rect 11057 25415 11115 25421
rect 11057 25381 11069 25415
rect 11103 25412 11115 25415
rect 11103 25384 12020 25412
rect 11103 25381 11115 25384
rect 11057 25375 11115 25381
rect 5442 25304 5448 25356
rect 5500 25344 5506 25356
rect 5997 25347 6055 25353
rect 5997 25344 6009 25347
rect 5500 25316 6009 25344
rect 5500 25304 5506 25316
rect 5997 25313 6009 25316
rect 6043 25313 6055 25347
rect 5997 25307 6055 25313
rect 7009 25347 7067 25353
rect 7009 25313 7021 25347
rect 7055 25344 7067 25347
rect 7098 25344 7104 25356
rect 7055 25316 7104 25344
rect 7055 25313 7067 25316
rect 7009 25307 7067 25313
rect 7098 25304 7104 25316
rect 7156 25304 7162 25356
rect 8205 25347 8263 25353
rect 8205 25313 8217 25347
rect 8251 25344 8263 25347
rect 9582 25344 9588 25356
rect 8251 25316 9588 25344
rect 8251 25313 8263 25316
rect 8205 25307 8263 25313
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 11882 25344 11888 25356
rect 11843 25316 11888 25344
rect 11882 25304 11888 25316
rect 11940 25304 11946 25356
rect 11992 25344 12020 25384
rect 16132 25344 16160 25452
rect 20162 25440 20168 25452
rect 20220 25440 20226 25492
rect 19426 25344 19432 25356
rect 11992 25316 16160 25344
rect 19387 25316 19432 25344
rect 19426 25304 19432 25316
rect 19484 25304 19490 25356
rect 19705 25347 19763 25353
rect 19705 25313 19717 25347
rect 19751 25344 19763 25347
rect 20714 25344 20720 25356
rect 19751 25316 20720 25344
rect 19751 25313 19763 25316
rect 19705 25307 19763 25313
rect 20714 25304 20720 25316
rect 20772 25304 20778 25356
rect 20898 25304 20904 25356
rect 20956 25344 20962 25356
rect 21177 25347 21235 25353
rect 21177 25344 21189 25347
rect 20956 25316 21189 25344
rect 20956 25304 20962 25316
rect 21177 25313 21189 25316
rect 21223 25313 21235 25347
rect 21177 25307 21235 25313
rect 2038 25276 2044 25288
rect 1999 25248 2044 25276
rect 2038 25236 2044 25248
rect 2096 25236 2102 25288
rect 4338 25276 4344 25288
rect 4299 25248 4344 25276
rect 4338 25236 4344 25248
rect 4396 25236 4402 25288
rect 4706 25236 4712 25288
rect 4764 25276 4770 25288
rect 5077 25279 5135 25285
rect 5077 25276 5089 25279
rect 4764 25248 5089 25276
rect 4764 25236 4770 25248
rect 5077 25245 5089 25248
rect 5123 25245 5135 25279
rect 5077 25239 5135 25245
rect 5205 25279 5263 25285
rect 5205 25245 5217 25279
rect 5251 25276 5263 25279
rect 5718 25276 5724 25288
rect 5251 25248 5724 25276
rect 5251 25245 5263 25248
rect 5205 25239 5263 25245
rect 1670 25168 1676 25220
rect 1728 25208 1734 25220
rect 2286 25211 2344 25217
rect 2286 25208 2298 25211
rect 1728 25180 2298 25208
rect 1728 25168 1734 25180
rect 2286 25177 2298 25180
rect 2332 25177 2344 25211
rect 4798 25208 4804 25220
rect 4759 25180 4804 25208
rect 2286 25171 2344 25177
rect 4798 25168 4804 25180
rect 4856 25168 4862 25220
rect 4985 25211 5043 25217
rect 4985 25177 4997 25211
rect 5031 25177 5043 25211
rect 5092 25208 5120 25239
rect 5718 25236 5724 25248
rect 5776 25236 5782 25288
rect 5902 25276 5908 25288
rect 5815 25248 5908 25276
rect 5902 25236 5908 25248
rect 5960 25276 5966 25288
rect 6546 25276 6552 25288
rect 5960 25248 6552 25276
rect 5960 25236 5966 25248
rect 6546 25236 6552 25248
rect 6604 25236 6610 25288
rect 8016 25279 8074 25285
rect 8016 25245 8028 25279
rect 8062 25276 8074 25279
rect 8478 25276 8484 25288
rect 8062 25248 8484 25276
rect 8062 25245 8074 25248
rect 8016 25239 8074 25245
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 9122 25236 9128 25288
rect 9180 25276 9186 25288
rect 9217 25279 9275 25285
rect 9217 25276 9229 25279
rect 9180 25248 9229 25276
rect 9180 25236 9186 25248
rect 9217 25245 9229 25248
rect 9263 25245 9275 25279
rect 9217 25239 9275 25245
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25245 9367 25279
rect 9490 25276 9496 25288
rect 9451 25248 9496 25276
rect 9309 25239 9367 25245
rect 5810 25208 5816 25220
rect 5092 25180 5816 25208
rect 4985 25171 5043 25177
rect 5000 25140 5028 25171
rect 5810 25168 5816 25180
rect 5868 25208 5874 25220
rect 7374 25208 7380 25220
rect 5868 25180 7380 25208
rect 5868 25168 5874 25180
rect 7374 25168 7380 25180
rect 7432 25208 7438 25220
rect 8110 25208 8116 25220
rect 7432 25180 8116 25208
rect 7432 25168 7438 25180
rect 8110 25168 8116 25180
rect 8168 25168 8174 25220
rect 8205 25211 8263 25217
rect 8205 25177 8217 25211
rect 8251 25208 8263 25211
rect 8294 25208 8300 25220
rect 8251 25180 8300 25208
rect 8251 25177 8263 25180
rect 8205 25171 8263 25177
rect 8294 25168 8300 25180
rect 8352 25168 8358 25220
rect 8389 25211 8447 25217
rect 8389 25177 8401 25211
rect 8435 25208 8447 25211
rect 8846 25208 8852 25220
rect 8435 25180 8852 25208
rect 8435 25177 8447 25180
rect 8389 25171 8447 25177
rect 8846 25168 8852 25180
rect 8904 25168 8910 25220
rect 5626 25140 5632 25152
rect 5000 25112 5632 25140
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 6362 25140 6368 25152
rect 6323 25112 6368 25140
rect 6362 25100 6368 25112
rect 6420 25100 6426 25152
rect 9214 25100 9220 25152
rect 9272 25140 9278 25152
rect 9324 25140 9352 25239
rect 9490 25236 9496 25248
rect 9548 25236 9554 25288
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25276 9735 25279
rect 10597 25279 10655 25285
rect 10597 25276 10609 25279
rect 9723 25248 10609 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 10597 25245 10609 25248
rect 10643 25276 10655 25279
rect 10686 25276 10692 25288
rect 10643 25248 10692 25276
rect 10643 25245 10655 25248
rect 10597 25239 10655 25245
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 10870 25276 10876 25288
rect 10831 25248 10876 25276
rect 10870 25236 10876 25248
rect 10928 25236 10934 25288
rect 13262 25236 13268 25288
rect 13320 25236 13326 25288
rect 15197 25279 15255 25285
rect 15197 25245 15209 25279
rect 15243 25276 15255 25279
rect 15562 25276 15568 25288
rect 15243 25248 15568 25276
rect 15243 25245 15255 25248
rect 15197 25239 15255 25245
rect 15562 25236 15568 25248
rect 15620 25236 15626 25288
rect 17402 25236 17408 25288
rect 17460 25276 17466 25288
rect 18141 25279 18199 25285
rect 17460 25248 17505 25276
rect 17460 25236 17466 25248
rect 18141 25245 18153 25279
rect 18187 25276 18199 25279
rect 18874 25276 18880 25288
rect 18187 25248 18880 25276
rect 18187 25245 18199 25248
rect 18141 25239 18199 25245
rect 18874 25236 18880 25248
rect 18932 25236 18938 25288
rect 20806 25236 20812 25288
rect 20864 25236 20870 25288
rect 12161 25211 12219 25217
rect 12161 25177 12173 25211
rect 12207 25208 12219 25211
rect 12434 25208 12440 25220
rect 12207 25180 12440 25208
rect 12207 25177 12219 25180
rect 12161 25171 12219 25177
rect 12434 25168 12440 25180
rect 12492 25168 12498 25220
rect 14918 25208 14924 25220
rect 14879 25180 14924 25208
rect 14918 25168 14924 25180
rect 14976 25168 14982 25220
rect 16574 25168 16580 25220
rect 16632 25168 16638 25220
rect 17129 25211 17187 25217
rect 17129 25177 17141 25211
rect 17175 25208 17187 25211
rect 17586 25208 17592 25220
rect 17175 25180 17592 25208
rect 17175 25177 17187 25180
rect 17129 25171 17187 25177
rect 17586 25168 17592 25180
rect 17644 25168 17650 25220
rect 18322 25168 18328 25220
rect 18380 25208 18386 25220
rect 18601 25211 18659 25217
rect 18601 25208 18613 25211
rect 18380 25180 18613 25208
rect 18380 25168 18386 25180
rect 18601 25177 18613 25180
rect 18647 25177 18659 25211
rect 18601 25171 18659 25177
rect 10686 25140 10692 25152
rect 9272 25112 9352 25140
rect 10647 25112 10692 25140
rect 9272 25100 9278 25112
rect 10686 25100 10692 25112
rect 10744 25100 10750 25152
rect 13998 25100 14004 25152
rect 14056 25140 14062 25152
rect 14277 25143 14335 25149
rect 14277 25140 14289 25143
rect 14056 25112 14289 25140
rect 14056 25100 14062 25112
rect 14277 25109 14289 25112
rect 14323 25140 14335 25143
rect 15102 25140 15108 25152
rect 14323 25112 15108 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 15102 25100 15108 25112
rect 15160 25140 15166 25152
rect 15286 25140 15292 25152
rect 15160 25112 15292 25140
rect 15160 25100 15166 25112
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 15657 25143 15715 25149
rect 15657 25109 15669 25143
rect 15703 25140 15715 25143
rect 17310 25140 17316 25152
rect 15703 25112 17316 25140
rect 15703 25109 15715 25112
rect 15657 25103 15715 25109
rect 17310 25100 17316 25112
rect 17368 25100 17374 25152
rect 17957 25143 18015 25149
rect 17957 25109 17969 25143
rect 18003 25140 18015 25143
rect 18046 25140 18052 25152
rect 18003 25112 18052 25140
rect 18003 25109 18015 25112
rect 17957 25103 18015 25109
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 1104 25050 28032 25072
rect 1104 24998 7642 25050
rect 7694 24998 7706 25050
rect 7758 24998 7770 25050
rect 7822 24998 7834 25050
rect 7886 24998 7898 25050
rect 7950 24998 14334 25050
rect 14386 24998 14398 25050
rect 14450 24998 14462 25050
rect 14514 24998 14526 25050
rect 14578 24998 14590 25050
rect 14642 24998 21026 25050
rect 21078 24998 21090 25050
rect 21142 24998 21154 25050
rect 21206 24998 21218 25050
rect 21270 24998 21282 25050
rect 21334 24998 27718 25050
rect 27770 24998 27782 25050
rect 27834 24998 27846 25050
rect 27898 24998 27910 25050
rect 27962 24998 27974 25050
rect 28026 24998 28032 25050
rect 1104 24976 28032 24998
rect 2225 24939 2283 24945
rect 2225 24905 2237 24939
rect 2271 24936 2283 24939
rect 2498 24936 2504 24948
rect 2271 24908 2504 24936
rect 2271 24905 2283 24908
rect 2225 24899 2283 24905
rect 2498 24896 2504 24908
rect 2556 24896 2562 24948
rect 4338 24896 4344 24948
rect 4396 24936 4402 24948
rect 5442 24936 5448 24948
rect 4396 24908 4844 24936
rect 5403 24908 5448 24936
rect 4396 24896 4402 24908
rect 4706 24868 4712 24880
rect 4667 24840 4712 24868
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 4816 24868 4844 24908
rect 5442 24896 5448 24908
rect 5500 24896 5506 24948
rect 5718 24936 5724 24948
rect 5631 24908 5724 24936
rect 5718 24896 5724 24908
rect 5776 24936 5782 24948
rect 6822 24936 6828 24948
rect 5776 24908 6828 24936
rect 5776 24896 5782 24908
rect 6822 24896 6828 24908
rect 6880 24896 6886 24948
rect 8478 24896 8484 24948
rect 8536 24936 8542 24948
rect 9125 24939 9183 24945
rect 9125 24936 9137 24939
rect 8536 24908 9137 24936
rect 8536 24896 8542 24908
rect 9125 24905 9137 24908
rect 9171 24905 9183 24939
rect 9125 24899 9183 24905
rect 9766 24896 9772 24948
rect 9824 24936 9830 24948
rect 9861 24939 9919 24945
rect 9861 24936 9873 24939
rect 9824 24908 9873 24936
rect 9824 24896 9830 24908
rect 9861 24905 9873 24908
rect 9907 24905 9919 24939
rect 9861 24899 9919 24905
rect 11149 24939 11207 24945
rect 11149 24905 11161 24939
rect 11195 24936 11207 24939
rect 11330 24936 11336 24948
rect 11195 24908 11336 24936
rect 11195 24905 11207 24908
rect 11149 24899 11207 24905
rect 11330 24896 11336 24908
rect 11388 24896 11394 24948
rect 13630 24936 13636 24948
rect 13543 24908 13636 24936
rect 13630 24896 13636 24908
rect 13688 24936 13694 24948
rect 15746 24936 15752 24948
rect 13688 24908 15752 24936
rect 13688 24896 13694 24908
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 20714 24936 20720 24948
rect 20675 24908 20720 24936
rect 20714 24896 20720 24908
rect 20772 24896 20778 24948
rect 6730 24868 6736 24880
rect 4816 24840 6736 24868
rect 3349 24803 3407 24809
rect 3349 24769 3361 24803
rect 3395 24800 3407 24803
rect 3970 24800 3976 24812
rect 3395 24772 3976 24800
rect 3395 24769 3407 24772
rect 3349 24763 3407 24769
rect 3970 24760 3976 24772
rect 4028 24760 4034 24812
rect 4816 24809 4844 24840
rect 6730 24828 6736 24840
rect 6788 24828 6794 24880
rect 8386 24828 8392 24880
rect 8444 24868 8450 24880
rect 9217 24871 9275 24877
rect 9217 24868 9229 24871
rect 8444 24840 9229 24868
rect 8444 24828 8450 24840
rect 9217 24837 9229 24840
rect 9263 24837 9275 24871
rect 9217 24831 9275 24837
rect 9401 24871 9459 24877
rect 9401 24837 9413 24871
rect 9447 24868 9459 24871
rect 9490 24868 9496 24880
rect 9447 24840 9496 24868
rect 9447 24837 9459 24840
rect 9401 24831 9459 24837
rect 9490 24828 9496 24840
rect 9548 24868 9554 24880
rect 9548 24840 10916 24868
rect 9548 24828 9554 24840
rect 4433 24803 4491 24809
rect 4433 24769 4445 24803
rect 4479 24769 4491 24803
rect 4433 24763 4491 24769
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 4801 24803 4859 24809
rect 4801 24769 4813 24803
rect 4847 24769 4859 24803
rect 5626 24800 5632 24812
rect 5587 24772 5632 24800
rect 4801 24763 4859 24769
rect 3602 24732 3608 24744
rect 3563 24704 3608 24732
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 4448 24664 4476 24763
rect 4632 24732 4660 24763
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 5810 24800 5816 24812
rect 5771 24772 5816 24800
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 7006 24800 7012 24812
rect 6967 24772 7012 24800
rect 7006 24760 7012 24772
rect 7064 24760 7070 24812
rect 7098 24760 7104 24812
rect 7156 24800 7162 24812
rect 7265 24803 7323 24809
rect 7265 24800 7277 24803
rect 7156 24772 7277 24800
rect 7156 24760 7162 24772
rect 7265 24769 7277 24772
rect 7311 24769 7323 24803
rect 7265 24763 7323 24769
rect 8110 24760 8116 24812
rect 8168 24800 8174 24812
rect 9033 24803 9091 24809
rect 9033 24800 9045 24803
rect 8168 24772 9045 24800
rect 8168 24760 8174 24772
rect 9033 24769 9045 24772
rect 9079 24769 9091 24803
rect 9033 24763 9091 24769
rect 9582 24760 9588 24812
rect 9640 24800 9646 24812
rect 10781 24803 10839 24809
rect 10781 24800 10793 24803
rect 9640 24772 10793 24800
rect 9640 24760 9646 24772
rect 10781 24769 10793 24772
rect 10827 24769 10839 24803
rect 10888 24800 10916 24840
rect 10965 24803 11023 24809
rect 10965 24800 10977 24803
rect 10888 24772 10977 24800
rect 10781 24763 10839 24769
rect 10965 24769 10977 24772
rect 11011 24769 11023 24803
rect 12066 24800 12072 24812
rect 12027 24772 12072 24800
rect 10965 24763 11023 24769
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 12158 24760 12164 24812
rect 12216 24800 12222 24812
rect 12526 24800 12532 24812
rect 12216 24772 12532 24800
rect 12216 24760 12222 24772
rect 12526 24760 12532 24772
rect 12584 24800 12590 24812
rect 13081 24803 13139 24809
rect 13081 24800 13093 24803
rect 12584 24772 13093 24800
rect 12584 24760 12590 24772
rect 13081 24769 13093 24772
rect 13127 24769 13139 24803
rect 13648 24786 13676 24896
rect 14829 24871 14887 24877
rect 14829 24837 14841 24871
rect 14875 24868 14887 24871
rect 14918 24868 14924 24880
rect 14875 24840 14924 24868
rect 14875 24837 14887 24840
rect 14829 24831 14887 24837
rect 14918 24828 14924 24840
rect 14976 24828 14982 24880
rect 16114 24868 16120 24880
rect 16054 24840 16120 24868
rect 16114 24828 16120 24840
rect 16172 24828 16178 24880
rect 17129 24871 17187 24877
rect 17129 24837 17141 24871
rect 17175 24868 17187 24871
rect 17402 24868 17408 24880
rect 17175 24840 17408 24868
rect 17175 24837 17187 24840
rect 17129 24831 17187 24837
rect 17402 24828 17408 24840
rect 17460 24828 17466 24880
rect 17586 24868 17592 24880
rect 17547 24840 17592 24868
rect 17586 24828 17592 24840
rect 17644 24828 17650 24880
rect 18598 24868 18604 24880
rect 18559 24840 18604 24868
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 14090 24800 14096 24812
rect 14051 24772 14096 24800
rect 13081 24763 13139 24769
rect 5718 24732 5724 24744
rect 4632 24704 5724 24732
rect 5718 24692 5724 24704
rect 5776 24692 5782 24744
rect 10321 24735 10379 24741
rect 10321 24701 10333 24735
rect 10367 24701 10379 24735
rect 10321 24695 10379 24701
rect 4798 24664 4804 24676
rect 4448 24636 4804 24664
rect 4798 24624 4804 24636
rect 4856 24664 4862 24676
rect 5997 24667 6055 24673
rect 5997 24664 6009 24667
rect 4856 24636 6009 24664
rect 4856 24624 4862 24636
rect 5997 24633 6009 24636
rect 6043 24664 6055 24667
rect 6270 24664 6276 24676
rect 6043 24636 6276 24664
rect 6043 24633 6055 24636
rect 5997 24627 6055 24633
rect 6270 24624 6276 24636
rect 6328 24624 6334 24676
rect 8846 24664 8852 24676
rect 8807 24636 8852 24664
rect 8846 24624 8852 24636
rect 8904 24624 8910 24676
rect 9490 24624 9496 24676
rect 9548 24664 9554 24676
rect 9953 24667 10011 24673
rect 9953 24664 9965 24667
rect 9548 24636 9965 24664
rect 9548 24624 9554 24636
rect 9953 24633 9965 24636
rect 9999 24633 10011 24667
rect 9953 24627 10011 24633
rect 4985 24599 5043 24605
rect 4985 24565 4997 24599
rect 5031 24596 5043 24599
rect 5902 24596 5908 24608
rect 5031 24568 5908 24596
rect 5031 24565 5043 24568
rect 4985 24559 5043 24565
rect 5902 24556 5908 24568
rect 5960 24556 5966 24608
rect 8294 24556 8300 24608
rect 8352 24596 8358 24608
rect 8389 24599 8447 24605
rect 8389 24596 8401 24599
rect 8352 24568 8401 24596
rect 8352 24556 8358 24568
rect 8389 24565 8401 24568
rect 8435 24596 8447 24599
rect 8478 24596 8484 24608
rect 8435 24568 8484 24596
rect 8435 24565 8447 24568
rect 8389 24559 8447 24565
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 9214 24556 9220 24608
rect 9272 24596 9278 24608
rect 10336 24596 10364 24695
rect 13096 24664 13124 24763
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 14553 24735 14611 24741
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 15470 24732 15476 24744
rect 14599 24704 15476 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 15470 24692 15476 24704
rect 15528 24692 15534 24744
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 16301 24735 16359 24741
rect 16301 24732 16313 24735
rect 15620 24704 16313 24732
rect 15620 24692 15626 24704
rect 16301 24701 16313 24704
rect 16347 24732 16359 24735
rect 16868 24732 16896 24763
rect 17310 24760 17316 24812
rect 17368 24800 17374 24812
rect 17681 24803 17739 24809
rect 17681 24800 17693 24803
rect 17368 24772 17693 24800
rect 17368 24760 17374 24772
rect 17681 24769 17693 24772
rect 17727 24769 17739 24803
rect 18322 24800 18328 24812
rect 18283 24772 18328 24800
rect 17681 24763 17739 24769
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 19702 24760 19708 24812
rect 19760 24760 19766 24812
rect 20898 24800 20904 24812
rect 20859 24772 20904 24800
rect 20898 24760 20904 24772
rect 20956 24760 20962 24812
rect 16347 24704 16896 24732
rect 16347 24701 16359 24704
rect 16301 24695 16359 24701
rect 13998 24664 14004 24676
rect 13096 24636 14004 24664
rect 13998 24624 14004 24636
rect 14056 24624 14062 24676
rect 9272 24568 10364 24596
rect 9272 24556 9278 24568
rect 11882 24556 11888 24608
rect 11940 24596 11946 24608
rect 12069 24599 12127 24605
rect 12069 24596 12081 24599
rect 11940 24568 12081 24596
rect 11940 24556 11946 24568
rect 12069 24565 12081 24568
rect 12115 24565 12127 24599
rect 12069 24559 12127 24565
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 20073 24599 20131 24605
rect 20073 24596 20085 24599
rect 19392 24568 20085 24596
rect 19392 24556 19398 24568
rect 20073 24565 20085 24568
rect 20119 24565 20131 24599
rect 20073 24559 20131 24565
rect 1104 24506 27876 24528
rect 1104 24454 4296 24506
rect 4348 24454 4360 24506
rect 4412 24454 4424 24506
rect 4476 24454 4488 24506
rect 4540 24454 4552 24506
rect 4604 24454 10988 24506
rect 11040 24454 11052 24506
rect 11104 24454 11116 24506
rect 11168 24454 11180 24506
rect 11232 24454 11244 24506
rect 11296 24454 17680 24506
rect 17732 24454 17744 24506
rect 17796 24454 17808 24506
rect 17860 24454 17872 24506
rect 17924 24454 17936 24506
rect 17988 24454 24372 24506
rect 24424 24454 24436 24506
rect 24488 24454 24500 24506
rect 24552 24454 24564 24506
rect 24616 24454 24628 24506
rect 24680 24454 27876 24506
rect 1104 24432 27876 24454
rect 3970 24392 3976 24404
rect 3931 24364 3976 24392
rect 3970 24352 3976 24364
rect 4028 24352 4034 24404
rect 6362 24352 6368 24404
rect 6420 24392 6426 24404
rect 7285 24395 7343 24401
rect 7285 24392 7297 24395
rect 6420 24364 7297 24392
rect 6420 24352 6426 24364
rect 7285 24361 7297 24364
rect 7331 24361 7343 24395
rect 7285 24355 7343 24361
rect 8573 24395 8631 24401
rect 8573 24361 8585 24395
rect 8619 24392 8631 24395
rect 9122 24392 9128 24404
rect 8619 24364 9128 24392
rect 8619 24361 8631 24364
rect 8573 24355 8631 24361
rect 9122 24352 9128 24364
rect 9180 24392 9186 24404
rect 9490 24392 9496 24404
rect 9180 24364 9496 24392
rect 9180 24352 9186 24364
rect 9490 24352 9496 24364
rect 9548 24352 9554 24404
rect 10686 24352 10692 24404
rect 10744 24392 10750 24404
rect 10965 24395 11023 24401
rect 10965 24392 10977 24395
rect 10744 24364 10977 24392
rect 10744 24352 10750 24364
rect 10965 24361 10977 24364
rect 11011 24361 11023 24395
rect 10965 24355 11023 24361
rect 12066 24352 12072 24404
rect 12124 24392 12130 24404
rect 13357 24395 13415 24401
rect 13357 24392 13369 24395
rect 12124 24364 13369 24392
rect 12124 24352 12130 24364
rect 13357 24361 13369 24364
rect 13403 24361 13415 24395
rect 13357 24355 13415 24361
rect 14182 24352 14188 24404
rect 14240 24392 14246 24404
rect 14369 24395 14427 24401
rect 14369 24392 14381 24395
rect 14240 24364 14381 24392
rect 14240 24352 14246 24364
rect 14369 24361 14381 24364
rect 14415 24361 14427 24395
rect 15102 24392 15108 24404
rect 15063 24364 15108 24392
rect 14369 24355 14427 24361
rect 15102 24352 15108 24364
rect 15160 24352 15166 24404
rect 6730 24324 6736 24336
rect 6691 24296 6736 24324
rect 6730 24284 6736 24296
rect 6788 24284 6794 24336
rect 8846 24324 8852 24336
rect 7116 24296 7604 24324
rect 4154 24216 4160 24268
rect 4212 24256 4218 24268
rect 4249 24259 4307 24265
rect 4249 24256 4261 24259
rect 4212 24228 4261 24256
rect 4212 24216 4218 24228
rect 4249 24225 4261 24228
rect 4295 24225 4307 24259
rect 5350 24256 5356 24268
rect 5311 24228 5356 24256
rect 4249 24219 4307 24225
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 2222 24197 2228 24200
rect 1949 24191 2007 24197
rect 1949 24157 1961 24191
rect 1995 24157 2007 24191
rect 2216 24188 2228 24197
rect 2183 24160 2228 24188
rect 1949 24151 2007 24157
rect 2216 24151 2228 24160
rect 1964 24120 1992 24151
rect 2222 24148 2228 24151
rect 2280 24148 2286 24200
rect 4341 24191 4399 24197
rect 4341 24157 4353 24191
rect 4387 24188 4399 24191
rect 4706 24188 4712 24200
rect 4387 24160 4712 24188
rect 4387 24157 4399 24160
rect 4341 24151 4399 24157
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 6362 24148 6368 24200
rect 6420 24188 6426 24200
rect 7116 24188 7144 24296
rect 6420 24160 7144 24188
rect 7193 24191 7251 24197
rect 6420 24148 6426 24160
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 2038 24120 2044 24132
rect 1951 24092 2044 24120
rect 2038 24080 2044 24092
rect 2096 24120 2102 24132
rect 3050 24120 3056 24132
rect 2096 24092 3056 24120
rect 2096 24080 2102 24092
rect 3050 24080 3056 24092
rect 3108 24120 3114 24132
rect 3602 24120 3608 24132
rect 3108 24092 3608 24120
rect 3108 24080 3114 24092
rect 3602 24080 3608 24092
rect 3660 24080 3666 24132
rect 5620 24123 5678 24129
rect 5620 24089 5632 24123
rect 5666 24089 5678 24123
rect 5620 24083 5678 24089
rect 3234 24012 3240 24064
rect 3292 24052 3298 24064
rect 3329 24055 3387 24061
rect 3329 24052 3341 24055
rect 3292 24024 3341 24052
rect 3292 24012 3298 24024
rect 3329 24021 3341 24024
rect 3375 24021 3387 24055
rect 3329 24015 3387 24021
rect 5534 24012 5540 24064
rect 5592 24052 5598 24064
rect 5644 24052 5672 24083
rect 5718 24080 5724 24132
rect 5776 24120 5782 24132
rect 7208 24120 7236 24151
rect 7374 24148 7380 24200
rect 7432 24197 7438 24200
rect 7576 24197 7604 24296
rect 8036 24296 8852 24324
rect 8036 24197 8064 24296
rect 8846 24284 8852 24296
rect 8904 24284 8910 24336
rect 8110 24216 8116 24268
rect 8168 24256 8174 24268
rect 9125 24259 9183 24265
rect 9125 24256 9137 24259
rect 8168 24228 9137 24256
rect 8168 24216 8174 24228
rect 9125 24225 9137 24228
rect 9171 24225 9183 24259
rect 11882 24256 11888 24268
rect 11843 24228 11888 24256
rect 9125 24219 9183 24225
rect 11882 24216 11888 24228
rect 11940 24216 11946 24268
rect 16574 24256 16580 24268
rect 16535 24228 16580 24256
rect 16574 24216 16580 24228
rect 16632 24216 16638 24268
rect 17126 24256 17132 24268
rect 17087 24228 17132 24256
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 17405 24259 17463 24265
rect 17405 24225 17417 24259
rect 17451 24256 17463 24259
rect 18046 24256 18052 24268
rect 17451 24228 18052 24256
rect 17451 24225 17463 24228
rect 17405 24219 17463 24225
rect 18046 24216 18052 24228
rect 18104 24216 18110 24268
rect 20070 24216 20076 24268
rect 20128 24256 20134 24268
rect 20257 24259 20315 24265
rect 20257 24256 20269 24259
rect 20128 24228 20269 24256
rect 20128 24216 20134 24228
rect 20257 24225 20269 24228
rect 20303 24225 20315 24259
rect 20257 24219 20315 24225
rect 15752 24200 15804 24206
rect 7432 24191 7454 24197
rect 7442 24157 7454 24191
rect 7432 24151 7454 24157
rect 7561 24191 7619 24197
rect 7561 24157 7573 24191
rect 7607 24188 7619 24191
rect 8021 24191 8079 24197
rect 8021 24188 8033 24191
rect 7607 24160 8033 24188
rect 7607 24157 7619 24160
rect 7561 24151 7619 24157
rect 8021 24157 8033 24160
rect 8067 24157 8079 24191
rect 8021 24151 8079 24157
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24188 8447 24191
rect 8435 24160 9076 24188
rect 8435 24157 8447 24160
rect 8389 24151 8447 24157
rect 7432 24148 7438 24151
rect 8202 24120 8208 24132
rect 5776 24092 7236 24120
rect 8163 24092 8208 24120
rect 5776 24080 5782 24092
rect 8202 24080 8208 24092
rect 8260 24080 8266 24132
rect 8297 24123 8355 24129
rect 8297 24089 8309 24123
rect 8343 24089 8355 24123
rect 8297 24083 8355 24089
rect 5592 24024 5672 24052
rect 5592 24012 5598 24024
rect 6730 24012 6736 24064
rect 6788 24052 6794 24064
rect 7285 24055 7343 24061
rect 7285 24052 7297 24055
rect 6788 24024 7297 24052
rect 6788 24012 6794 24024
rect 7285 24021 7297 24024
rect 7331 24021 7343 24055
rect 7285 24015 7343 24021
rect 7466 24012 7472 24064
rect 7524 24052 7530 24064
rect 8018 24052 8024 24064
rect 7524 24024 8024 24052
rect 7524 24012 7530 24024
rect 8018 24012 8024 24024
rect 8076 24052 8082 24064
rect 8312 24052 8340 24083
rect 8076 24024 8340 24052
rect 9048 24052 9076 24160
rect 10594 24148 10600 24200
rect 10652 24188 10658 24200
rect 10870 24188 10876 24200
rect 10652 24160 10876 24188
rect 10652 24148 10658 24160
rect 10870 24148 10876 24160
rect 10928 24188 10934 24200
rect 10965 24191 11023 24197
rect 10965 24188 10977 24191
rect 10928 24160 10977 24188
rect 10928 24148 10934 24160
rect 10965 24157 10977 24160
rect 11011 24157 11023 24191
rect 10965 24151 11023 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24157 11207 24191
rect 11606 24188 11612 24200
rect 11567 24160 11612 24188
rect 11149 24151 11207 24157
rect 9398 24129 9404 24132
rect 9392 24120 9404 24129
rect 9359 24092 9404 24120
rect 9392 24083 9404 24092
rect 9398 24080 9404 24083
rect 9456 24080 9462 24132
rect 11164 24120 11192 24151
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24188 14611 24191
rect 15010 24188 15016 24200
rect 14599 24160 15016 24188
rect 14599 24157 14611 24160
rect 14553 24151 14611 24157
rect 15010 24148 15016 24160
rect 15068 24148 15074 24200
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 15657 24191 15715 24197
rect 15657 24188 15669 24191
rect 15160 24160 15669 24188
rect 15160 24148 15166 24160
rect 15657 24157 15669 24160
rect 15703 24157 15715 24191
rect 15657 24151 15715 24157
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 19886 24148 19892 24200
rect 19944 24148 19950 24200
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 20993 24191 21051 24197
rect 20993 24188 21005 24191
rect 20956 24160 21005 24188
rect 20956 24148 20962 24160
rect 20993 24157 21005 24160
rect 21039 24157 21051 24191
rect 20993 24151 21051 24157
rect 15752 24142 15804 24148
rect 11514 24120 11520 24132
rect 11164 24092 11520 24120
rect 11514 24080 11520 24092
rect 11572 24080 11578 24132
rect 13170 24120 13176 24132
rect 13110 24092 13176 24120
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 19702 24120 19708 24132
rect 19663 24092 19708 24120
rect 19702 24080 19708 24092
rect 19760 24080 19766 24132
rect 21269 24123 21327 24129
rect 21269 24089 21281 24123
rect 21315 24120 21327 24123
rect 21450 24120 21456 24132
rect 21315 24092 21456 24120
rect 21315 24089 21327 24092
rect 21269 24083 21327 24089
rect 21450 24080 21456 24092
rect 21508 24080 21514 24132
rect 9582 24052 9588 24064
rect 9048 24024 9588 24052
rect 8076 24012 8082 24024
rect 9582 24012 9588 24024
rect 9640 24052 9646 24064
rect 10505 24055 10563 24061
rect 10505 24052 10517 24055
rect 9640 24024 10517 24052
rect 9640 24012 9646 24024
rect 10505 24021 10517 24024
rect 10551 24021 10563 24055
rect 18874 24052 18880 24064
rect 18835 24024 18880 24052
rect 10505 24015 10563 24021
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 1104 23962 28032 23984
rect 1104 23910 7642 23962
rect 7694 23910 7706 23962
rect 7758 23910 7770 23962
rect 7822 23910 7834 23962
rect 7886 23910 7898 23962
rect 7950 23910 14334 23962
rect 14386 23910 14398 23962
rect 14450 23910 14462 23962
rect 14514 23910 14526 23962
rect 14578 23910 14590 23962
rect 14642 23910 21026 23962
rect 21078 23910 21090 23962
rect 21142 23910 21154 23962
rect 21206 23910 21218 23962
rect 21270 23910 21282 23962
rect 21334 23910 27718 23962
rect 27770 23910 27782 23962
rect 27834 23910 27846 23962
rect 27898 23910 27910 23962
rect 27962 23910 27974 23962
rect 28026 23910 28032 23962
rect 1104 23888 28032 23910
rect 1670 23848 1676 23860
rect 1631 23820 1676 23848
rect 1670 23808 1676 23820
rect 1728 23808 1734 23860
rect 5626 23808 5632 23860
rect 5684 23848 5690 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 5684 23820 5825 23848
rect 5684 23808 5690 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 5813 23811 5871 23817
rect 6917 23851 6975 23857
rect 6917 23817 6929 23851
rect 6963 23848 6975 23851
rect 7098 23848 7104 23860
rect 6963 23820 7104 23848
rect 6963 23817 6975 23820
rect 6917 23811 6975 23817
rect 7098 23808 7104 23820
rect 7156 23808 7162 23860
rect 7745 23851 7803 23857
rect 7745 23817 7757 23851
rect 7791 23848 7803 23851
rect 8110 23848 8116 23860
rect 7791 23820 8116 23848
rect 7791 23817 7803 23820
rect 7745 23811 7803 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 8202 23808 8208 23860
rect 8260 23848 8266 23860
rect 8665 23851 8723 23857
rect 8665 23848 8677 23851
rect 8260 23820 8677 23848
rect 8260 23808 8266 23820
rect 8665 23817 8677 23820
rect 8711 23817 8723 23851
rect 8665 23811 8723 23817
rect 8849 23851 8907 23857
rect 8849 23817 8861 23851
rect 8895 23848 8907 23851
rect 9214 23848 9220 23860
rect 8895 23820 9220 23848
rect 8895 23817 8907 23820
rect 8849 23811 8907 23817
rect 9214 23808 9220 23820
rect 9272 23808 9278 23860
rect 9398 23848 9404 23860
rect 9359 23820 9404 23848
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 13449 23851 13507 23857
rect 13449 23817 13461 23851
rect 13495 23848 13507 23851
rect 13630 23848 13636 23860
rect 13495 23820 13636 23848
rect 13495 23817 13507 23820
rect 13449 23811 13507 23817
rect 13630 23808 13636 23820
rect 13688 23808 13694 23860
rect 18141 23851 18199 23857
rect 18141 23817 18153 23851
rect 18187 23817 18199 23851
rect 18141 23811 18199 23817
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 8481 23783 8539 23789
rect 8481 23780 8493 23783
rect 8076 23752 8493 23780
rect 8076 23740 8082 23752
rect 8481 23749 8493 23752
rect 8527 23749 8539 23783
rect 8481 23743 8539 23749
rect 8573 23783 8631 23789
rect 8573 23749 8585 23783
rect 8619 23780 8631 23783
rect 14737 23783 14795 23789
rect 8619 23752 9628 23780
rect 8619 23749 8631 23752
rect 8573 23743 8631 23749
rect 9600 23724 9628 23752
rect 14737 23749 14749 23783
rect 14783 23780 14795 23783
rect 18156 23780 18184 23811
rect 19886 23808 19892 23860
rect 19944 23848 19950 23860
rect 20162 23848 20168 23860
rect 19944 23820 20168 23848
rect 19944 23808 19950 23820
rect 20162 23808 20168 23820
rect 20220 23848 20226 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 20220 23820 20361 23848
rect 20220 23808 20226 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 20349 23811 20407 23817
rect 19061 23783 19119 23789
rect 19061 23780 19073 23783
rect 14783 23752 19073 23780
rect 14783 23749 14795 23752
rect 14737 23743 14795 23749
rect 19061 23749 19073 23752
rect 19107 23749 19119 23783
rect 19061 23743 19119 23749
rect 2797 23715 2855 23721
rect 2797 23681 2809 23715
rect 2843 23712 2855 23715
rect 2958 23712 2964 23724
rect 2843 23684 2964 23712
rect 2843 23681 2855 23684
rect 2797 23675 2855 23681
rect 2958 23672 2964 23684
rect 3016 23672 3022 23724
rect 3510 23712 3516 23724
rect 3471 23684 3516 23712
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 4706 23721 4712 23724
rect 4700 23712 4712 23721
rect 4667 23684 4712 23712
rect 4700 23675 4712 23684
rect 4706 23672 4712 23675
rect 4764 23672 4770 23724
rect 7101 23715 7159 23721
rect 7101 23681 7113 23715
rect 7147 23712 7159 23715
rect 7561 23715 7619 23721
rect 7561 23712 7573 23715
rect 7147 23684 7573 23712
rect 7147 23681 7159 23684
rect 7101 23675 7159 23681
rect 7561 23681 7573 23684
rect 7607 23712 7619 23715
rect 8294 23712 8300 23724
rect 7607 23684 8300 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 8294 23672 8300 23684
rect 8352 23672 8358 23724
rect 9582 23712 9588 23724
rect 9543 23684 9588 23712
rect 9582 23672 9588 23684
rect 9640 23672 9646 23724
rect 12066 23712 12072 23724
rect 12027 23684 12072 23712
rect 12066 23672 12072 23684
rect 12124 23672 12130 23724
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 3050 23604 3056 23656
rect 3108 23644 3114 23656
rect 3326 23644 3332 23656
rect 3108 23616 3332 23644
rect 3108 23604 3114 23616
rect 3326 23604 3332 23616
rect 3384 23604 3390 23656
rect 4154 23604 4160 23656
rect 4212 23644 4218 23656
rect 4433 23647 4491 23653
rect 4433 23644 4445 23647
rect 4212 23616 4445 23644
rect 4212 23604 4218 23616
rect 4433 23613 4445 23616
rect 4479 23613 4491 23647
rect 11974 23644 11980 23656
rect 11935 23616 11980 23644
rect 4433 23607 4491 23613
rect 11974 23604 11980 23616
rect 12032 23604 12038 23656
rect 6270 23536 6276 23588
rect 6328 23576 6334 23588
rect 8297 23579 8355 23585
rect 8297 23576 8309 23579
rect 6328 23548 8309 23576
rect 6328 23536 6334 23548
rect 8297 23545 8309 23548
rect 8343 23545 8355 23579
rect 12158 23576 12164 23588
rect 8297 23539 8355 23545
rect 10520 23548 12164 23576
rect 3697 23511 3755 23517
rect 3697 23477 3709 23511
rect 3743 23508 3755 23511
rect 8478 23508 8484 23520
rect 3743 23480 8484 23508
rect 3743 23477 3755 23480
rect 3697 23471 3755 23477
rect 8478 23468 8484 23480
rect 8536 23508 8542 23520
rect 9490 23508 9496 23520
rect 8536 23480 9496 23508
rect 8536 23468 8542 23480
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 9766 23468 9772 23520
rect 9824 23508 9830 23520
rect 10520 23517 10548 23548
rect 12158 23536 12164 23548
rect 12216 23536 12222 23588
rect 10505 23511 10563 23517
rect 10505 23508 10517 23511
rect 9824 23480 10517 23508
rect 9824 23468 9830 23480
rect 10505 23477 10517 23480
rect 10551 23477 10563 23511
rect 10505 23471 10563 23477
rect 11149 23511 11207 23517
rect 11149 23477 11161 23511
rect 11195 23508 11207 23511
rect 12250 23508 12256 23520
rect 11195 23480 12256 23508
rect 11195 23477 11207 23480
rect 11149 23471 11207 23477
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 12437 23511 12495 23517
rect 12437 23477 12449 23511
rect 12483 23508 12495 23511
rect 15378 23508 15384 23520
rect 12483 23480 15384 23508
rect 12483 23477 12495 23480
rect 12437 23471 12495 23477
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 1104 23418 27876 23440
rect 1104 23366 4296 23418
rect 4348 23366 4360 23418
rect 4412 23366 4424 23418
rect 4476 23366 4488 23418
rect 4540 23366 4552 23418
rect 4604 23366 10988 23418
rect 11040 23366 11052 23418
rect 11104 23366 11116 23418
rect 11168 23366 11180 23418
rect 11232 23366 11244 23418
rect 11296 23366 17680 23418
rect 17732 23366 17744 23418
rect 17796 23366 17808 23418
rect 17860 23366 17872 23418
rect 17924 23366 17936 23418
rect 17988 23366 24372 23418
rect 24424 23366 24436 23418
rect 24488 23366 24500 23418
rect 24552 23366 24564 23418
rect 24616 23366 24628 23418
rect 24680 23366 27876 23418
rect 1104 23344 27876 23366
rect 5629 23307 5687 23313
rect 5629 23273 5641 23307
rect 5675 23304 5687 23307
rect 5718 23304 5724 23316
rect 5675 23276 5724 23304
rect 5675 23273 5687 23276
rect 5629 23267 5687 23273
rect 5718 23264 5724 23276
rect 5776 23264 5782 23316
rect 7745 23307 7803 23313
rect 7745 23273 7757 23307
rect 7791 23304 7803 23307
rect 8202 23304 8208 23316
rect 7791 23276 8208 23304
rect 7791 23273 7803 23276
rect 7745 23267 7803 23273
rect 8202 23264 8208 23276
rect 8260 23264 8266 23316
rect 9490 23304 9496 23316
rect 9451 23276 9496 23304
rect 9490 23264 9496 23276
rect 9548 23264 9554 23316
rect 16853 23307 16911 23313
rect 16853 23273 16865 23307
rect 16899 23273 16911 23307
rect 16853 23267 16911 23273
rect 21195 23307 21253 23313
rect 21195 23273 21207 23307
rect 21241 23304 21253 23307
rect 21913 23307 21971 23313
rect 21913 23304 21925 23307
rect 21241 23276 21925 23304
rect 21241 23273 21253 23276
rect 21195 23267 21253 23273
rect 21913 23273 21925 23276
rect 21959 23273 21971 23307
rect 21913 23267 21971 23273
rect 10689 23239 10747 23245
rect 10689 23205 10701 23239
rect 10735 23205 10747 23239
rect 16868 23236 16896 23267
rect 18690 23236 18696 23248
rect 16868 23208 18696 23236
rect 10689 23199 10747 23205
rect 4154 23128 4160 23180
rect 4212 23168 4218 23180
rect 4249 23171 4307 23177
rect 4249 23168 4261 23171
rect 4212 23140 4261 23168
rect 4212 23128 4218 23140
rect 4249 23137 4261 23140
rect 4295 23137 4307 23171
rect 4249 23131 4307 23137
rect 3073 23103 3131 23109
rect 3073 23069 3085 23103
rect 3119 23100 3131 23103
rect 3234 23100 3240 23112
rect 3119 23072 3240 23100
rect 3119 23069 3131 23072
rect 3073 23063 3131 23069
rect 3234 23060 3240 23072
rect 3292 23060 3298 23112
rect 3326 23060 3332 23112
rect 3384 23100 3390 23112
rect 3878 23100 3884 23112
rect 3384 23072 3884 23100
rect 3384 23060 3390 23072
rect 3878 23060 3884 23072
rect 3936 23060 3942 23112
rect 4264 23100 4292 23131
rect 6362 23100 6368 23112
rect 4264 23072 6368 23100
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 8205 23103 8263 23109
rect 8205 23100 8217 23103
rect 6840 23072 8217 23100
rect 6840 23044 6868 23072
rect 8205 23069 8217 23072
rect 8251 23069 8263 23103
rect 8205 23063 8263 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23100 10287 23103
rect 10704 23100 10732 23199
rect 18690 23196 18696 23208
rect 18748 23196 18754 23248
rect 11333 23171 11391 23177
rect 11333 23137 11345 23171
rect 11379 23168 11391 23171
rect 11422 23168 11428 23180
rect 11379 23140 11428 23168
rect 11379 23137 11391 23140
rect 11333 23131 11391 23137
rect 11422 23128 11428 23140
rect 11480 23128 11486 23180
rect 13170 23168 13176 23180
rect 13131 23140 13176 23168
rect 13170 23128 13176 23140
rect 13228 23128 13234 23180
rect 14737 23171 14795 23177
rect 14737 23137 14749 23171
rect 14783 23137 14795 23171
rect 14737 23131 14795 23137
rect 15013 23171 15071 23177
rect 15013 23137 15025 23171
rect 15059 23168 15071 23171
rect 15470 23168 15476 23180
rect 15059 23140 15476 23168
rect 15059 23137 15071 23140
rect 15013 23131 15071 23137
rect 11146 23100 11152 23112
rect 10275 23072 10732 23100
rect 11059 23072 11152 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 11146 23060 11152 23072
rect 11204 23100 11210 23112
rect 11974 23100 11980 23112
rect 11204 23072 11980 23100
rect 11204 23060 11210 23072
rect 11974 23060 11980 23072
rect 12032 23060 12038 23112
rect 12158 23100 12164 23112
rect 12119 23072 12164 23100
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 13630 23100 13636 23112
rect 12834 23072 13636 23100
rect 13630 23060 13636 23072
rect 13688 23060 13694 23112
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23069 14703 23103
rect 14752 23100 14780 23131
rect 15470 23128 15476 23140
rect 15528 23128 15534 23180
rect 18506 23168 18512 23180
rect 18467 23140 18512 23168
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 20162 23168 20168 23180
rect 18892 23140 20168 23168
rect 18236 23112 18288 23118
rect 15194 23100 15200 23112
rect 14752 23072 15200 23100
rect 14645 23063 14703 23069
rect 4516 23035 4574 23041
rect 4516 23001 4528 23035
rect 4562 23032 4574 23035
rect 4614 23032 4620 23044
rect 4562 23004 4620 23032
rect 4562 23001 4574 23004
rect 4516 22995 4574 23001
rect 4614 22992 4620 23004
rect 4672 22992 4678 23044
rect 5718 22992 5724 23044
rect 5776 23032 5782 23044
rect 6610 23035 6668 23041
rect 6610 23032 6622 23035
rect 5776 23004 6622 23032
rect 5776 22992 5782 23004
rect 6610 23001 6622 23004
rect 6656 23001 6668 23035
rect 6610 22995 6668 23001
rect 6822 22992 6828 23044
rect 6880 22992 6886 23044
rect 9490 22992 9496 23044
rect 9548 23032 9554 23044
rect 11057 23035 11115 23041
rect 11057 23032 11069 23035
rect 9548 23004 11069 23032
rect 9548 22992 9554 23004
rect 11057 23001 11069 23004
rect 11103 23032 11115 23035
rect 12618 23032 12624 23044
rect 11103 23004 12624 23032
rect 11103 23001 11115 23004
rect 11057 22995 11115 23001
rect 12618 22992 12624 23004
rect 12676 22992 12682 23044
rect 14660 23032 14688 23063
rect 15194 23060 15200 23072
rect 15252 23060 15258 23112
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 16761 23103 16819 23109
rect 16761 23100 16773 23103
rect 15344 23072 16773 23100
rect 15344 23060 15350 23072
rect 16761 23069 16773 23072
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 16853 23103 16911 23109
rect 16853 23069 16865 23103
rect 16899 23100 16911 23103
rect 17218 23100 17224 23112
rect 16899 23072 17224 23100
rect 16899 23069 16911 23072
rect 16853 23063 16911 23069
rect 17218 23060 17224 23072
rect 17276 23060 17282 23112
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 15010 23032 15016 23044
rect 14660 23004 15016 23032
rect 15010 22992 15016 23004
rect 15068 22992 15074 23044
rect 16298 22992 16304 23044
rect 16356 23032 16362 23044
rect 16577 23035 16635 23041
rect 16577 23032 16589 23035
rect 16356 23004 16589 23032
rect 16356 22992 16362 23004
rect 16577 23001 16589 23004
rect 16623 23001 16635 23035
rect 16577 22995 16635 23001
rect 1949 22967 2007 22973
rect 1949 22933 1961 22967
rect 1995 22964 2007 22967
rect 2038 22964 2044 22976
rect 1995 22936 2044 22964
rect 1995 22933 2007 22936
rect 1949 22927 2007 22933
rect 2038 22924 2044 22936
rect 2096 22924 2102 22976
rect 8294 22924 8300 22976
rect 8352 22964 8358 22976
rect 8389 22967 8447 22973
rect 8389 22964 8401 22967
rect 8352 22936 8401 22964
rect 8352 22924 8358 22936
rect 8389 22933 8401 22936
rect 8435 22933 8447 22967
rect 10042 22964 10048 22976
rect 10003 22936 10048 22964
rect 8389 22927 8447 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 13722 22964 13728 22976
rect 13683 22936 13728 22964
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 17034 22964 17040 22976
rect 16995 22936 17040 22964
rect 17034 22924 17040 22936
rect 17092 22924 17098 22976
rect 17604 22964 17632 23063
rect 18892 23100 18920 23140
rect 20162 23128 20168 23140
rect 20220 23128 20226 23180
rect 21450 23168 21456 23180
rect 21411 23140 21456 23168
rect 21450 23128 21456 23140
rect 21508 23128 21514 23180
rect 18288 23072 18920 23100
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23069 21971 23103
rect 21913 23063 21971 23069
rect 18236 23054 18288 23060
rect 20714 22992 20720 23044
rect 20772 22992 20778 23044
rect 18414 22964 18420 22976
rect 17604 22936 18420 22964
rect 18414 22924 18420 22936
rect 18472 22964 18478 22976
rect 19242 22964 19248 22976
rect 18472 22936 19248 22964
rect 18472 22924 18478 22936
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 19705 22967 19763 22973
rect 19705 22933 19717 22967
rect 19751 22964 19763 22967
rect 20438 22964 20444 22976
rect 19751 22936 20444 22964
rect 19751 22933 19763 22936
rect 19705 22927 19763 22933
rect 20438 22924 20444 22936
rect 20496 22964 20502 22976
rect 21928 22964 21956 23063
rect 20496 22936 21956 22964
rect 20496 22924 20502 22936
rect 1104 22874 28032 22896
rect 1104 22822 7642 22874
rect 7694 22822 7706 22874
rect 7758 22822 7770 22874
rect 7822 22822 7834 22874
rect 7886 22822 7898 22874
rect 7950 22822 14334 22874
rect 14386 22822 14398 22874
rect 14450 22822 14462 22874
rect 14514 22822 14526 22874
rect 14578 22822 14590 22874
rect 14642 22822 21026 22874
rect 21078 22822 21090 22874
rect 21142 22822 21154 22874
rect 21206 22822 21218 22874
rect 21270 22822 21282 22874
rect 21334 22822 27718 22874
rect 27770 22822 27782 22874
rect 27834 22822 27846 22874
rect 27898 22822 27910 22874
rect 27962 22822 27974 22874
rect 28026 22822 28032 22874
rect 1104 22800 28032 22822
rect 3421 22763 3479 22769
rect 3421 22729 3433 22763
rect 3467 22760 3479 22763
rect 3510 22760 3516 22772
rect 3467 22732 3516 22760
rect 3467 22729 3479 22732
rect 3421 22723 3479 22729
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 8297 22763 8355 22769
rect 8297 22729 8309 22763
rect 8343 22760 8355 22763
rect 8386 22760 8392 22772
rect 8343 22732 8392 22760
rect 8343 22729 8355 22732
rect 8297 22723 8355 22729
rect 8386 22720 8392 22732
rect 8444 22720 8450 22772
rect 11146 22760 11152 22772
rect 11107 22732 11152 22760
rect 11146 22720 11152 22732
rect 11204 22720 11210 22772
rect 11606 22720 11612 22772
rect 11664 22760 11670 22772
rect 11793 22763 11851 22769
rect 11793 22760 11805 22763
rect 11664 22732 11805 22760
rect 11664 22720 11670 22732
rect 11793 22729 11805 22732
rect 11839 22729 11851 22763
rect 11793 22723 11851 22729
rect 15013 22763 15071 22769
rect 15013 22729 15025 22763
rect 15059 22760 15071 22763
rect 15194 22760 15200 22772
rect 15059 22732 15200 22760
rect 15059 22729 15071 22732
rect 15013 22723 15071 22729
rect 15194 22720 15200 22732
rect 15252 22720 15258 22772
rect 20898 22760 20904 22772
rect 19168 22732 20904 22760
rect 10042 22701 10048 22704
rect 10036 22692 10048 22701
rect 10003 22664 10048 22692
rect 10036 22655 10048 22664
rect 10042 22652 10048 22655
rect 10100 22652 10106 22704
rect 12434 22652 12440 22704
rect 12492 22692 12498 22704
rect 13357 22695 13415 22701
rect 13357 22692 13369 22695
rect 12492 22664 13369 22692
rect 12492 22652 12498 22664
rect 13357 22661 13369 22664
rect 13403 22661 13415 22695
rect 13357 22655 13415 22661
rect 13722 22652 13728 22704
rect 13780 22692 13786 22704
rect 14921 22695 14979 22701
rect 14921 22692 14933 22695
rect 13780 22664 14933 22692
rect 13780 22652 13786 22664
rect 14921 22661 14933 22664
rect 14967 22692 14979 22695
rect 18966 22692 18972 22704
rect 14967 22664 18972 22692
rect 14967 22661 14979 22664
rect 14921 22655 14979 22661
rect 18966 22652 18972 22664
rect 19024 22652 19030 22704
rect 2133 22627 2191 22633
rect 2133 22593 2145 22627
rect 2179 22624 2191 22627
rect 2958 22624 2964 22636
rect 2179 22596 2964 22624
rect 2179 22593 2191 22596
rect 2133 22587 2191 22593
rect 2958 22584 2964 22596
rect 3016 22624 3022 22636
rect 4706 22624 4712 22636
rect 3016 22596 4712 22624
rect 3016 22584 3022 22596
rect 4706 22584 4712 22596
rect 4764 22584 4770 22636
rect 6362 22584 6368 22636
rect 6420 22624 6426 22636
rect 6638 22624 6644 22636
rect 6420 22596 6644 22624
rect 6420 22584 6426 22596
rect 6638 22584 6644 22596
rect 6696 22624 6702 22636
rect 6917 22627 6975 22633
rect 6917 22624 6929 22627
rect 6696 22596 6929 22624
rect 6696 22584 6702 22596
rect 6917 22593 6929 22596
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7184 22627 7242 22633
rect 7184 22593 7196 22627
rect 7230 22624 7242 22627
rect 8202 22624 8208 22636
rect 7230 22596 8208 22624
rect 7230 22593 7242 22596
rect 7184 22587 7242 22593
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22624 11943 22627
rect 12158 22624 12164 22636
rect 11931 22596 12164 22624
rect 11931 22593 11943 22596
rect 11885 22587 11943 22593
rect 12158 22584 12164 22596
rect 12216 22584 12222 22636
rect 12529 22627 12587 22633
rect 12529 22593 12541 22627
rect 12575 22624 12587 22627
rect 12710 22624 12716 22636
rect 12575 22596 12716 22624
rect 12575 22593 12587 22596
rect 12529 22587 12587 22593
rect 12710 22584 12716 22596
rect 12768 22624 12774 22636
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 12768 22596 13461 22624
rect 12768 22584 12774 22596
rect 13449 22593 13461 22596
rect 13495 22593 13507 22627
rect 15286 22624 15292 22636
rect 13449 22587 13507 22593
rect 15028 22596 15292 22624
rect 2038 22556 2044 22568
rect 1999 22528 2044 22556
rect 2038 22516 2044 22528
rect 2096 22516 2102 22568
rect 9214 22516 9220 22568
rect 9272 22556 9278 22568
rect 9309 22559 9367 22565
rect 9309 22556 9321 22559
rect 9272 22528 9321 22556
rect 9272 22516 9278 22528
rect 9309 22525 9321 22528
rect 9355 22556 9367 22559
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9355 22528 9781 22556
rect 9355 22525 9367 22528
rect 9309 22519 9367 22525
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 9769 22519 9827 22525
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 12897 22559 12955 22565
rect 12492 22528 12537 22556
rect 12492 22516 12498 22528
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 15028 22556 15056 22596
rect 15286 22584 15292 22596
rect 15344 22584 15350 22636
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 15933 22627 15991 22633
rect 15933 22624 15945 22627
rect 15620 22596 15945 22624
rect 15620 22584 15626 22596
rect 15933 22593 15945 22596
rect 15979 22593 15991 22627
rect 15933 22587 15991 22593
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22624 17647 22627
rect 18874 22624 18880 22636
rect 17635 22596 18880 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 19068 22627 19126 22633
rect 19068 22593 19080 22627
rect 19114 22624 19126 22627
rect 19168 22624 19196 22732
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 19242 22652 19248 22704
rect 19300 22652 19306 22704
rect 20714 22652 20720 22704
rect 20772 22692 20778 22704
rect 20809 22695 20867 22701
rect 20809 22692 20821 22695
rect 20772 22664 20821 22692
rect 20772 22652 20778 22664
rect 20809 22661 20821 22664
rect 20855 22661 20867 22695
rect 20809 22655 20867 22661
rect 19114 22596 19196 22624
rect 19260 22624 19288 22652
rect 19794 22624 19800 22636
rect 19260 22596 19800 22624
rect 19114 22593 19126 22596
rect 19068 22587 19126 22593
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 20162 22584 20168 22636
rect 20220 22584 20226 22636
rect 12943 22528 15056 22556
rect 15105 22559 15163 22565
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 15105 22525 15117 22559
rect 15151 22525 15163 22559
rect 15838 22556 15844 22568
rect 15799 22528 15844 22556
rect 15105 22519 15163 22525
rect 14918 22448 14924 22500
rect 14976 22488 14982 22500
rect 15120 22488 15148 22519
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 16298 22556 16304 22568
rect 16259 22528 16304 22556
rect 16298 22516 16304 22528
rect 16356 22516 16362 22568
rect 17218 22556 17224 22568
rect 17179 22528 17224 22556
rect 17218 22516 17224 22528
rect 17276 22516 17282 22568
rect 17494 22556 17500 22568
rect 17455 22528 17500 22556
rect 17494 22516 17500 22528
rect 17552 22516 17558 22568
rect 18690 22556 18696 22568
rect 18651 22528 18696 22556
rect 18690 22516 18696 22528
rect 18748 22516 18754 22568
rect 18969 22559 19027 22565
rect 18969 22525 18981 22559
rect 19015 22525 19027 22559
rect 18969 22519 19027 22525
rect 14976 22460 15148 22488
rect 18984 22488 19012 22519
rect 19242 22516 19248 22568
rect 19300 22556 19306 22568
rect 19300 22528 20024 22556
rect 19300 22516 19306 22528
rect 19426 22488 19432 22500
rect 18984 22460 19432 22488
rect 14976 22448 14982 22460
rect 19426 22448 19432 22460
rect 19484 22448 19490 22500
rect 1765 22423 1823 22429
rect 1765 22389 1777 22423
rect 1811 22420 1823 22423
rect 1854 22420 1860 22432
rect 1811 22392 1860 22420
rect 1811 22389 1823 22392
rect 1765 22383 1823 22389
rect 1854 22380 1860 22392
rect 1912 22380 1918 22432
rect 3510 22380 3516 22432
rect 3568 22420 3574 22432
rect 4341 22423 4399 22429
rect 4341 22420 4353 22423
rect 3568 22392 4353 22420
rect 3568 22380 3574 22392
rect 4341 22389 4353 22392
rect 4387 22420 4399 22423
rect 5169 22423 5227 22429
rect 5169 22420 5181 22423
rect 4387 22392 5181 22420
rect 4387 22389 4399 22392
rect 4341 22383 4399 22389
rect 5169 22389 5181 22392
rect 5215 22389 5227 22423
rect 5169 22383 5227 22389
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 14553 22423 14611 22429
rect 14553 22420 14565 22423
rect 13872 22392 14565 22420
rect 13872 22380 13878 22392
rect 14553 22389 14565 22392
rect 14599 22389 14611 22423
rect 19996 22420 20024 22528
rect 21361 22423 21419 22429
rect 21361 22420 21373 22423
rect 19996 22392 21373 22420
rect 14553 22383 14611 22389
rect 21361 22389 21373 22392
rect 21407 22420 21419 22423
rect 22002 22420 22008 22432
rect 21407 22392 22008 22420
rect 21407 22389 21419 22392
rect 21361 22383 21419 22389
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 1104 22330 27876 22352
rect 1104 22278 4296 22330
rect 4348 22278 4360 22330
rect 4412 22278 4424 22330
rect 4476 22278 4488 22330
rect 4540 22278 4552 22330
rect 4604 22278 10988 22330
rect 11040 22278 11052 22330
rect 11104 22278 11116 22330
rect 11168 22278 11180 22330
rect 11232 22278 11244 22330
rect 11296 22278 17680 22330
rect 17732 22278 17744 22330
rect 17796 22278 17808 22330
rect 17860 22278 17872 22330
rect 17924 22278 17936 22330
rect 17988 22278 24372 22330
rect 24424 22278 24436 22330
rect 24488 22278 24500 22330
rect 24552 22278 24564 22330
rect 24616 22278 24628 22330
rect 24680 22278 27876 22330
rect 1104 22256 27876 22278
rect 4706 22176 4712 22228
rect 4764 22216 4770 22228
rect 5721 22219 5779 22225
rect 5721 22216 5733 22219
rect 4764 22188 5733 22216
rect 4764 22176 4770 22188
rect 5721 22185 5733 22188
rect 5767 22185 5779 22219
rect 5721 22179 5779 22185
rect 6822 22176 6828 22228
rect 6880 22216 6886 22228
rect 7193 22219 7251 22225
rect 7193 22216 7205 22219
rect 6880 22188 7205 22216
rect 6880 22176 6886 22188
rect 7193 22185 7205 22188
rect 7239 22185 7251 22219
rect 7193 22179 7251 22185
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 13725 22219 13783 22225
rect 11388 22188 12434 22216
rect 11388 22176 11394 22188
rect 11425 22151 11483 22157
rect 11425 22117 11437 22151
rect 11471 22148 11483 22151
rect 12406 22148 12434 22188
rect 13725 22185 13737 22219
rect 13771 22185 13783 22219
rect 13725 22179 13783 22185
rect 11471 22120 11505 22148
rect 12406 22120 12480 22148
rect 11471 22117 11483 22120
rect 11425 22111 11483 22117
rect 4249 22083 4307 22089
rect 4249 22049 4261 22083
rect 4295 22080 4307 22083
rect 4614 22080 4620 22092
rect 4295 22052 4620 22080
rect 4295 22049 4307 22052
rect 4249 22043 4307 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 11440 22080 11468 22111
rect 12452 22089 12480 22120
rect 12437 22083 12495 22089
rect 9416 22052 10180 22080
rect 11440 22052 12112 22080
rect 3878 21972 3884 22024
rect 3936 22012 3942 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3936 21984 3985 22012
rect 3936 21972 3942 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 8294 22012 8300 22024
rect 8352 22021 8358 22024
rect 8264 21984 8300 22012
rect 8294 21972 8300 21984
rect 8352 21975 8364 22021
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 9306 22012 9312 22024
rect 8619 21984 9312 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 8352 21972 8358 21975
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 9416 22021 9444 22052
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 21981 9459 22015
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 9401 21975 9459 21981
rect 9508 21984 10057 22012
rect 9214 21904 9220 21956
rect 9272 21944 9278 21956
rect 9508 21944 9536 21984
rect 10045 21981 10057 21984
rect 10091 21981 10103 22015
rect 10152 22012 10180 22052
rect 10152 21984 11928 22012
rect 10045 21975 10103 21981
rect 10290 21947 10348 21953
rect 10290 21944 10302 21947
rect 9272 21916 9536 21944
rect 9600 21916 10302 21944
rect 9272 21904 9278 21916
rect 1670 21876 1676 21888
rect 1631 21848 1676 21876
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 2593 21879 2651 21885
rect 2593 21845 2605 21879
rect 2639 21876 2651 21879
rect 3237 21879 3295 21885
rect 3237 21876 3249 21879
rect 2639 21848 3249 21876
rect 2639 21845 2651 21848
rect 2593 21839 2651 21845
rect 3237 21845 3249 21848
rect 3283 21876 3295 21879
rect 3510 21876 3516 21888
rect 3283 21848 3516 21876
rect 3283 21845 3295 21848
rect 3237 21839 3295 21845
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 9600 21885 9628 21916
rect 10290 21913 10302 21916
rect 10336 21913 10348 21947
rect 10290 21907 10348 21913
rect 11900 21885 11928 21984
rect 12084 21944 12112 22052
rect 12437 22049 12449 22083
rect 12483 22049 12495 22083
rect 13740 22080 13768 22179
rect 15194 22176 15200 22228
rect 15252 22216 15258 22228
rect 15657 22219 15715 22225
rect 15657 22216 15669 22219
rect 15252 22188 15669 22216
rect 15252 22176 15258 22188
rect 15657 22185 15669 22188
rect 15703 22185 15715 22219
rect 15657 22179 15715 22185
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 20806 22216 20812 22228
rect 19484 22188 20812 22216
rect 19484 22176 19490 22188
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 20073 22083 20131 22089
rect 13740 22052 14412 22080
rect 12437 22043 12495 22049
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 13814 22012 13820 22024
rect 13587 21984 13820 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 21981 14335 22015
rect 14384 22012 14412 22052
rect 20073 22049 20085 22083
rect 20119 22049 20131 22083
rect 20346 22080 20352 22092
rect 20307 22052 20352 22080
rect 20073 22043 20131 22049
rect 14533 22015 14591 22021
rect 14533 22012 14545 22015
rect 14384 21984 14545 22012
rect 14277 21975 14335 21981
rect 14533 21981 14545 21984
rect 14579 21981 14591 22015
rect 16206 22012 16212 22024
rect 16167 21984 16212 22012
rect 14533 21975 14591 21981
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12084 21916 12357 21944
rect 12345 21913 12357 21916
rect 12391 21944 12403 21947
rect 12434 21944 12440 21956
rect 12391 21916 12440 21944
rect 12391 21913 12403 21916
rect 12345 21907 12403 21913
rect 12434 21904 12440 21916
rect 12492 21904 12498 21956
rect 13722 21904 13728 21956
rect 13780 21944 13786 21956
rect 14292 21944 14320 21975
rect 16206 21972 16212 21984
rect 16264 21972 16270 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16316 21984 16865 22012
rect 16316 21944 16344 21984
rect 16853 21981 16865 21984
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 17402 21972 17408 22024
rect 17460 22012 17466 22024
rect 20088 22012 20116 22043
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20438 22012 20444 22024
rect 17460 21984 20116 22012
rect 20399 21984 20444 22012
rect 17460 21972 17466 21984
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 20898 21972 20904 22024
rect 20956 22012 20962 22024
rect 21085 22015 21143 22021
rect 21085 22012 21097 22015
rect 20956 21984 21097 22012
rect 20956 21972 20962 21984
rect 21085 21981 21097 21984
rect 21131 21981 21143 22015
rect 21726 22012 21732 22024
rect 21687 21984 21732 22012
rect 21085 21975 21143 21981
rect 21726 21972 21732 21984
rect 21784 21972 21790 22024
rect 22002 22021 22008 22024
rect 21996 22012 22008 22021
rect 21963 21984 22008 22012
rect 21996 21975 22008 21984
rect 22002 21972 22008 21975
rect 22060 21972 22066 22024
rect 17098 21947 17156 21953
rect 17098 21944 17110 21947
rect 13780 21916 16344 21944
rect 16408 21916 17110 21944
rect 13780 21904 13786 21916
rect 6641 21879 6699 21885
rect 6641 21876 6653 21879
rect 6604 21848 6653 21876
rect 6604 21836 6610 21848
rect 6641 21845 6653 21848
rect 6687 21845 6699 21879
rect 6641 21839 6699 21845
rect 9585 21879 9643 21885
rect 9585 21845 9597 21879
rect 9631 21845 9643 21879
rect 9585 21839 9643 21845
rect 11885 21879 11943 21885
rect 11885 21845 11897 21879
rect 11931 21845 11943 21879
rect 12250 21876 12256 21888
rect 12211 21848 12256 21876
rect 11885 21839 11943 21845
rect 12250 21836 12256 21848
rect 12308 21876 12314 21888
rect 16298 21876 16304 21888
rect 12308 21848 16304 21876
rect 12308 21836 12314 21848
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 16408 21885 16436 21916
rect 17098 21913 17110 21916
rect 17144 21913 17156 21947
rect 17098 21907 17156 21913
rect 16393 21879 16451 21885
rect 16393 21845 16405 21879
rect 16439 21845 16451 21879
rect 16393 21839 16451 21845
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 18233 21879 18291 21885
rect 18233 21876 18245 21879
rect 17552 21848 18245 21876
rect 17552 21836 17558 21848
rect 18233 21845 18245 21848
rect 18279 21845 18291 21879
rect 18690 21876 18696 21888
rect 18651 21848 18696 21876
rect 18233 21839 18291 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19518 21876 19524 21888
rect 19479 21848 19524 21876
rect 19518 21836 19524 21848
rect 19576 21836 19582 21888
rect 21269 21879 21327 21885
rect 21269 21845 21281 21879
rect 21315 21876 21327 21879
rect 21358 21876 21364 21888
rect 21315 21848 21364 21876
rect 21315 21845 21327 21848
rect 21269 21839 21327 21845
rect 21358 21836 21364 21848
rect 21416 21836 21422 21888
rect 23109 21879 23167 21885
rect 23109 21845 23121 21879
rect 23155 21876 23167 21879
rect 23474 21876 23480 21888
rect 23155 21848 23480 21876
rect 23155 21845 23167 21848
rect 23109 21839 23167 21845
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 1104 21786 28032 21808
rect 1104 21734 7642 21786
rect 7694 21734 7706 21786
rect 7758 21734 7770 21786
rect 7822 21734 7834 21786
rect 7886 21734 7898 21786
rect 7950 21734 14334 21786
rect 14386 21734 14398 21786
rect 14450 21734 14462 21786
rect 14514 21734 14526 21786
rect 14578 21734 14590 21786
rect 14642 21734 21026 21786
rect 21078 21734 21090 21786
rect 21142 21734 21154 21786
rect 21206 21734 21218 21786
rect 21270 21734 21282 21786
rect 21334 21734 27718 21786
rect 27770 21734 27782 21786
rect 27834 21734 27846 21786
rect 27898 21734 27910 21786
rect 27962 21734 27974 21786
rect 28026 21734 28032 21786
rect 1104 21712 28032 21734
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 4111 21675 4169 21681
rect 3568 21644 4016 21672
rect 3568 21632 3574 21644
rect 3418 21564 3424 21616
rect 3476 21564 3482 21616
rect 3988 21604 4016 21644
rect 4111 21641 4123 21675
rect 4157 21672 4169 21675
rect 4614 21672 4620 21684
rect 4157 21644 4620 21672
rect 4157 21641 4169 21644
rect 4111 21635 4169 21641
rect 4614 21632 4620 21644
rect 4672 21632 4678 21684
rect 5350 21672 5356 21684
rect 5311 21644 5356 21672
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 14921 21675 14979 21681
rect 14921 21641 14933 21675
rect 14967 21672 14979 21675
rect 15194 21672 15200 21684
rect 14967 21644 15200 21672
rect 14967 21641 14979 21644
rect 14921 21635 14979 21641
rect 15194 21632 15200 21644
rect 15252 21672 15258 21684
rect 15838 21672 15844 21684
rect 15252 21644 15844 21672
rect 15252 21632 15258 21644
rect 15838 21632 15844 21644
rect 15896 21632 15902 21684
rect 16206 21632 16212 21684
rect 16264 21672 16270 21684
rect 16945 21675 17003 21681
rect 16945 21672 16957 21675
rect 16264 21644 16957 21672
rect 16264 21632 16270 21644
rect 16945 21641 16957 21644
rect 16991 21641 17003 21675
rect 16945 21635 17003 21641
rect 17405 21675 17463 21681
rect 17405 21641 17417 21675
rect 17451 21672 17463 21675
rect 17494 21672 17500 21684
rect 17451 21644 17500 21672
rect 17451 21641 17463 21644
rect 17405 21635 17463 21641
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 19521 21675 19579 21681
rect 19521 21641 19533 21675
rect 19567 21672 19579 21675
rect 20346 21672 20352 21684
rect 19567 21644 20352 21672
rect 19567 21641 19579 21644
rect 19521 21635 19579 21641
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 22002 21632 22008 21684
rect 22060 21672 22066 21684
rect 23385 21675 23443 21681
rect 22060 21632 22094 21672
rect 23385 21641 23397 21675
rect 23431 21672 23443 21675
rect 26326 21672 26332 21684
rect 23431 21644 26332 21672
rect 23431 21641 23443 21644
rect 23385 21635 23443 21641
rect 26326 21632 26332 21644
rect 26384 21632 26390 21684
rect 6546 21604 6552 21616
rect 3988 21576 6552 21604
rect 3970 21496 3976 21548
rect 4028 21536 4034 21548
rect 4801 21539 4859 21545
rect 4801 21536 4813 21539
rect 4028 21508 4813 21536
rect 4028 21496 4034 21508
rect 4801 21505 4813 21508
rect 4847 21536 4859 21539
rect 4982 21536 4988 21548
rect 4847 21508 4988 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 5350 21536 5356 21548
rect 5311 21508 5356 21536
rect 5350 21496 5356 21508
rect 5408 21496 5414 21548
rect 5552 21545 5580 21576
rect 6546 21564 6552 21576
rect 6604 21564 6610 21616
rect 7466 21564 7472 21616
rect 7524 21564 7530 21616
rect 13004 21576 15700 21604
rect 10042 21545 10048 21548
rect 5537 21539 5595 21545
rect 5537 21505 5549 21539
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 10036 21499 10048 21545
rect 10100 21536 10106 21548
rect 12158 21536 12164 21548
rect 10100 21508 10136 21536
rect 12119 21508 12164 21536
rect 10042 21496 10048 21499
rect 10100 21496 10106 21508
rect 12158 21496 12164 21508
rect 12216 21496 12222 21548
rect 1486 21428 1492 21480
rect 1544 21468 1550 21480
rect 2317 21471 2375 21477
rect 2317 21468 2329 21471
rect 1544 21440 2329 21468
rect 1544 21428 1550 21440
rect 2317 21437 2329 21440
rect 2363 21437 2375 21471
rect 2682 21468 2688 21480
rect 2643 21440 2688 21468
rect 2317 21431 2375 21437
rect 2682 21428 2688 21440
rect 2740 21428 2746 21480
rect 3878 21428 3884 21480
rect 3936 21468 3942 21480
rect 4617 21471 4675 21477
rect 4617 21468 4629 21471
rect 3936 21440 4629 21468
rect 3936 21428 3942 21440
rect 4617 21437 4629 21440
rect 4663 21437 4675 21471
rect 5000 21468 5028 21496
rect 6549 21471 6607 21477
rect 6549 21468 6561 21471
rect 5000 21440 6561 21468
rect 4617 21431 4675 21437
rect 6549 21437 6561 21440
rect 6595 21437 6607 21471
rect 6822 21468 6828 21480
rect 6783 21440 6828 21468
rect 6549 21431 6607 21437
rect 6822 21428 6828 21440
rect 6880 21428 6886 21480
rect 7374 21428 7380 21480
rect 7432 21468 7438 21480
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 7432 21440 9781 21468
rect 7432 21428 7438 21440
rect 9769 21437 9781 21440
rect 9815 21437 9827 21471
rect 11330 21468 11336 21480
rect 9769 21431 9827 21437
rect 11164 21440 11336 21468
rect 11164 21409 11192 21440
rect 11330 21428 11336 21440
rect 11388 21468 11394 21480
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 11388 21440 12081 21468
rect 11388 21428 11394 21440
rect 12069 21437 12081 21440
rect 12115 21437 12127 21471
rect 12069 21431 12127 21437
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 13004 21468 13032 21576
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 15672 21545 15700 21576
rect 16298 21564 16304 21616
rect 16356 21604 16362 21616
rect 17313 21607 17371 21613
rect 17313 21604 17325 21607
rect 16356 21576 17325 21604
rect 16356 21564 16362 21576
rect 17313 21573 17325 21576
rect 17359 21604 17371 21607
rect 18690 21604 18696 21616
rect 17359 21576 18696 21604
rect 17359 21573 17371 21576
rect 17313 21567 17371 21573
rect 18690 21564 18696 21576
rect 18748 21564 18754 21616
rect 22066 21604 22094 21632
rect 22250 21607 22308 21613
rect 22250 21604 22262 21607
rect 22066 21576 22262 21604
rect 22250 21573 22262 21576
rect 22296 21573 22308 21607
rect 22250 21567 22308 21573
rect 13797 21539 13855 21545
rect 13797 21536 13809 21539
rect 13136 21508 13809 21536
rect 13136 21496 13142 21508
rect 13797 21505 13809 21508
rect 13843 21505 13855 21539
rect 13797 21499 13855 21505
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21536 15439 21539
rect 15657 21539 15715 21545
rect 15427 21508 15608 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 12575 21440 13032 21468
rect 13541 21471 13599 21477
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 13541 21437 13553 21471
rect 13587 21437 13599 21471
rect 15470 21468 15476 21480
rect 15431 21440 15476 21468
rect 13541 21431 13599 21437
rect 11149 21403 11207 21409
rect 11149 21369 11161 21403
rect 11195 21369 11207 21403
rect 11149 21363 11207 21369
rect 12342 21360 12348 21412
rect 12400 21400 12406 21412
rect 12989 21403 13047 21409
rect 12989 21400 13001 21403
rect 12400 21372 13001 21400
rect 12400 21360 12406 21372
rect 12989 21369 13001 21372
rect 13035 21369 13047 21403
rect 12989 21363 13047 21369
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 8297 21335 8355 21341
rect 8297 21332 8309 21335
rect 8260 21304 8309 21332
rect 8260 21292 8266 21304
rect 8297 21301 8309 21304
rect 8343 21301 8355 21335
rect 9214 21332 9220 21344
rect 9175 21304 9220 21332
rect 8297 21295 8355 21301
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 13556 21332 13584 21431
rect 15470 21428 15476 21440
rect 15528 21428 15534 21480
rect 15580 21468 15608 21508
rect 15657 21505 15669 21539
rect 15703 21505 15715 21539
rect 18138 21536 18144 21548
rect 18099 21508 18144 21536
rect 15657 21499 15715 21505
rect 18138 21496 18144 21508
rect 18196 21496 18202 21548
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21536 18935 21539
rect 19794 21536 19800 21548
rect 18923 21508 19800 21536
rect 18923 21505 18935 21508
rect 18877 21499 18935 21505
rect 19794 21496 19800 21508
rect 19852 21496 19858 21548
rect 20645 21539 20703 21545
rect 20645 21505 20657 21539
rect 20691 21536 20703 21539
rect 21266 21536 21272 21548
rect 20691 21508 21272 21536
rect 20691 21505 20703 21508
rect 20645 21499 20703 21505
rect 21266 21496 21272 21508
rect 21324 21496 21330 21548
rect 21358 21496 21364 21548
rect 21416 21536 21422 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21416 21508 22017 21536
rect 21416 21496 21422 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 17402 21468 17408 21480
rect 15580 21440 17408 21468
rect 17402 21428 17408 21440
rect 17460 21428 17466 21480
rect 17497 21471 17555 21477
rect 17497 21437 17509 21471
rect 17543 21437 17555 21471
rect 17497 21431 17555 21437
rect 20901 21471 20959 21477
rect 20901 21437 20913 21471
rect 20947 21468 20959 21471
rect 21910 21468 21916 21480
rect 20947 21440 21916 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 14918 21360 14924 21412
rect 14976 21400 14982 21412
rect 17512 21400 17540 21431
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 14976 21372 17540 21400
rect 14976 21360 14982 21372
rect 13722 21332 13728 21344
rect 13556 21304 13728 21332
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 15378 21332 15384 21344
rect 15339 21304 15384 21332
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15838 21332 15844 21344
rect 15799 21304 15844 21332
rect 15838 21292 15844 21304
rect 15896 21292 15902 21344
rect 18322 21332 18328 21344
rect 18283 21304 18328 21332
rect 18322 21292 18328 21304
rect 18380 21292 18386 21344
rect 19058 21332 19064 21344
rect 19019 21304 19064 21332
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 21358 21332 21364 21344
rect 21319 21304 21364 21332
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 1104 21242 27876 21264
rect 1104 21190 4296 21242
rect 4348 21190 4360 21242
rect 4412 21190 4424 21242
rect 4476 21190 4488 21242
rect 4540 21190 4552 21242
rect 4604 21190 10988 21242
rect 11040 21190 11052 21242
rect 11104 21190 11116 21242
rect 11168 21190 11180 21242
rect 11232 21190 11244 21242
rect 11296 21190 17680 21242
rect 17732 21190 17744 21242
rect 17796 21190 17808 21242
rect 17860 21190 17872 21242
rect 17924 21190 17936 21242
rect 17988 21190 24372 21242
rect 24424 21190 24436 21242
rect 24488 21190 24500 21242
rect 24552 21190 24564 21242
rect 24616 21190 24628 21242
rect 24680 21190 27876 21242
rect 1104 21168 27876 21190
rect 1627 21131 1685 21137
rect 1627 21097 1639 21131
rect 1673 21128 1685 21131
rect 2682 21128 2688 21140
rect 1673 21100 2688 21128
rect 1673 21097 1685 21100
rect 1627 21091 1685 21097
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 6822 21088 6828 21140
rect 6880 21137 6886 21140
rect 6880 21131 6929 21137
rect 6880 21097 6883 21131
rect 6917 21097 6929 21131
rect 7466 21128 7472 21140
rect 7427 21100 7472 21128
rect 6880 21091 6929 21097
rect 6880 21088 6886 21091
rect 7466 21088 7472 21100
rect 7524 21088 7530 21140
rect 10042 21088 10048 21140
rect 10100 21128 10106 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 10100 21100 10149 21128
rect 10100 21088 10106 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 11330 21088 11336 21140
rect 11388 21088 11394 21140
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 16853 21131 16911 21137
rect 16853 21128 16865 21131
rect 14200 21100 16865 21128
rect 10781 21063 10839 21069
rect 10781 21029 10793 21063
rect 10827 21029 10839 21063
rect 11348 21060 11376 21088
rect 10781 21023 10839 21029
rect 11256 21032 11376 21060
rect 1486 20952 1492 21004
rect 1544 20992 1550 21004
rect 3421 20995 3479 21001
rect 3421 20992 3433 20995
rect 1544 20964 3433 20992
rect 1544 20952 1550 20964
rect 3421 20961 3433 20964
rect 3467 20992 3479 20995
rect 3878 20992 3884 21004
rect 3467 20964 3884 20992
rect 3467 20961 3479 20964
rect 3421 20955 3479 20961
rect 3878 20952 3884 20964
rect 3936 20952 3942 21004
rect 8202 20992 8208 21004
rect 4356 20964 8208 20992
rect 3053 20927 3111 20933
rect 3053 20893 3065 20927
rect 3099 20924 3111 20927
rect 4356 20924 4384 20964
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 3099 20896 4384 20924
rect 4433 20927 4491 20933
rect 3099 20893 3111 20896
rect 3053 20887 3111 20893
rect 4433 20893 4445 20927
rect 4479 20893 4491 20927
rect 4433 20887 4491 20893
rect 4617 20927 4675 20933
rect 4617 20893 4629 20927
rect 4663 20924 4675 20927
rect 4798 20924 4804 20936
rect 4663 20896 4804 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 2714 20828 2820 20856
rect 2792 20800 2820 20828
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 4448 20856 4476 20887
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 4982 20884 4988 20936
rect 5040 20924 5046 20936
rect 5077 20927 5135 20933
rect 5077 20924 5089 20927
rect 5040 20896 5089 20924
rect 5040 20884 5046 20896
rect 5077 20893 5089 20896
rect 5123 20893 5135 20927
rect 5077 20887 5135 20893
rect 5445 20927 5503 20933
rect 5445 20893 5457 20927
rect 5491 20924 5503 20927
rect 5534 20924 5540 20936
rect 5491 20896 5540 20924
rect 5491 20893 5503 20896
rect 5445 20887 5503 20893
rect 5534 20884 5540 20896
rect 5592 20884 5598 20936
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 6972 20896 7389 20924
rect 6972 20884 6978 20896
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 7466 20884 7472 20936
rect 7524 20924 7530 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7524 20896 7573 20924
rect 7524 20884 7530 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20924 10379 20927
rect 10796 20924 10824 21023
rect 11256 21001 11284 21032
rect 12158 21020 12164 21072
rect 12216 21060 12222 21072
rect 14200 21060 14228 21100
rect 16853 21097 16865 21100
rect 16899 21128 16911 21131
rect 18138 21128 18144 21140
rect 16899 21100 18144 21128
rect 16899 21097 16911 21100
rect 16853 21091 16911 21097
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 20901 21131 20959 21137
rect 20901 21128 20913 21131
rect 20864 21100 20913 21128
rect 20864 21088 20870 21100
rect 20901 21097 20913 21100
rect 20947 21097 20959 21131
rect 20901 21091 20959 21097
rect 21266 21088 21272 21140
rect 21324 21128 21330 21140
rect 21361 21131 21419 21137
rect 21361 21128 21373 21131
rect 21324 21100 21373 21128
rect 21324 21088 21330 21100
rect 21361 21097 21373 21100
rect 21407 21097 21419 21131
rect 21361 21091 21419 21097
rect 12216 21032 14228 21060
rect 14277 21063 14335 21069
rect 12216 21020 12222 21032
rect 14277 21029 14289 21063
rect 14323 21029 14335 21063
rect 14277 21023 14335 21029
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11422 20992 11428 21004
rect 11383 20964 11428 20992
rect 11241 20955 11299 20961
rect 11422 20952 11428 20964
rect 11480 20952 11486 21004
rect 14292 20992 14320 21023
rect 14918 20992 14924 21004
rect 12912 20964 14320 20992
rect 14879 20964 14924 20992
rect 12342 20924 12348 20936
rect 10367 20896 10824 20924
rect 11808 20896 12348 20924
rect 10367 20893 10379 20896
rect 10321 20887 10379 20893
rect 3568 20828 4476 20856
rect 3568 20816 3574 20828
rect 6454 20816 6460 20868
rect 6512 20816 6518 20868
rect 9214 20816 9220 20868
rect 9272 20856 9278 20868
rect 11054 20856 11060 20868
rect 9272 20828 11060 20856
rect 9272 20816 9278 20828
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 11808 20800 11836 20896
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 12912 20933 12940 20964
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 15838 20992 15844 21004
rect 15799 20964 15844 20992
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 18322 20992 18328 21004
rect 18283 20964 18328 20992
rect 18322 20952 18328 20964
rect 18380 20952 18386 21004
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 19116 20964 19656 20992
rect 19116 20952 19122 20964
rect 12897 20927 12955 20933
rect 12897 20893 12909 20927
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20924 13599 20927
rect 14182 20924 14188 20936
rect 13587 20896 14188 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 15194 20924 15200 20936
rect 14783 20896 15200 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 16022 20924 16028 20936
rect 15983 20896 16028 20924
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20924 16175 20927
rect 17034 20924 17040 20936
rect 16163 20896 17040 20924
rect 16163 20893 16175 20896
rect 16117 20887 16175 20893
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 18598 20884 18604 20936
rect 18656 20924 18662 20936
rect 19521 20927 19579 20933
rect 18656 20896 18701 20924
rect 18656 20884 18662 20896
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19628 20924 19656 20964
rect 19777 20927 19835 20933
rect 19777 20924 19789 20927
rect 19628 20896 19789 20924
rect 19521 20887 19579 20893
rect 19777 20893 19789 20896
rect 19823 20893 19835 20927
rect 21542 20924 21548 20936
rect 21503 20896 21548 20924
rect 19777 20887 19835 20893
rect 12360 20856 12388 20884
rect 14645 20859 14703 20865
rect 14645 20856 14657 20859
rect 12360 20828 14657 20856
rect 14645 20825 14657 20828
rect 14691 20825 14703 20859
rect 14645 20819 14703 20825
rect 17310 20816 17316 20868
rect 17368 20816 17374 20868
rect 19536 20856 19564 20887
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 21910 20884 21916 20936
rect 21968 20924 21974 20936
rect 22189 20927 22247 20933
rect 22189 20924 22201 20927
rect 21968 20896 22201 20924
rect 21968 20884 21974 20896
rect 22189 20893 22201 20896
rect 22235 20893 22247 20927
rect 22189 20887 22247 20893
rect 21928 20856 21956 20884
rect 19536 20828 21956 20856
rect 22456 20859 22514 20865
rect 22456 20825 22468 20859
rect 22502 20856 22514 20859
rect 23474 20856 23480 20868
rect 22502 20828 23480 20856
rect 22502 20825 22514 20828
rect 22456 20819 22514 20825
rect 23474 20816 23480 20828
rect 23532 20816 23538 20868
rect 2774 20748 2780 20800
rect 2832 20748 2838 20800
rect 4617 20791 4675 20797
rect 4617 20757 4629 20791
rect 4663 20788 4675 20791
rect 4706 20788 4712 20800
rect 4663 20760 4712 20788
rect 4663 20757 4675 20760
rect 4617 20751 4675 20757
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 5350 20788 5356 20800
rect 4856 20760 5356 20788
rect 4856 20748 4862 20760
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 7006 20748 7012 20800
rect 7064 20788 7070 20800
rect 8021 20791 8079 20797
rect 8021 20788 8033 20791
rect 7064 20760 8033 20788
rect 7064 20748 7070 20760
rect 8021 20757 8033 20760
rect 8067 20757 8079 20791
rect 9674 20788 9680 20800
rect 9635 20760 9680 20788
rect 8021 20751 8079 20757
rect 9674 20748 9680 20760
rect 9732 20788 9738 20800
rect 11149 20791 11207 20797
rect 11149 20788 11161 20791
rect 9732 20760 11161 20788
rect 9732 20748 9738 20760
rect 11149 20757 11161 20760
rect 11195 20788 11207 20791
rect 11790 20788 11796 20800
rect 11195 20760 11796 20788
rect 11195 20757 11207 20760
rect 11149 20751 11207 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 13725 20791 13783 20797
rect 13725 20757 13737 20791
rect 13771 20788 13783 20791
rect 14090 20788 14096 20800
rect 13771 20760 14096 20788
rect 13771 20757 13783 20760
rect 13725 20751 13783 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 16114 20788 16120 20800
rect 16075 20760 16120 20788
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 23569 20791 23627 20797
rect 23569 20757 23581 20791
rect 23615 20788 23627 20791
rect 23658 20788 23664 20800
rect 23615 20760 23664 20788
rect 23615 20757 23627 20760
rect 23569 20751 23627 20757
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 1104 20698 28032 20720
rect 1104 20646 7642 20698
rect 7694 20646 7706 20698
rect 7758 20646 7770 20698
rect 7822 20646 7834 20698
rect 7886 20646 7898 20698
rect 7950 20646 14334 20698
rect 14386 20646 14398 20698
rect 14450 20646 14462 20698
rect 14514 20646 14526 20698
rect 14578 20646 14590 20698
rect 14642 20646 21026 20698
rect 21078 20646 21090 20698
rect 21142 20646 21154 20698
rect 21206 20646 21218 20698
rect 21270 20646 21282 20698
rect 21334 20646 27718 20698
rect 27770 20646 27782 20698
rect 27834 20646 27846 20698
rect 27898 20646 27910 20698
rect 27962 20646 27974 20698
rect 28026 20646 28032 20698
rect 1104 20624 28032 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 3418 20584 3424 20596
rect 2832 20556 2877 20584
rect 3379 20556 3424 20584
rect 2832 20544 2838 20556
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 4890 20584 4896 20596
rect 3528 20556 4896 20584
rect 3234 20516 3240 20528
rect 2700 20488 3240 20516
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 2700 20457 2728 20488
rect 3234 20476 3240 20488
rect 3292 20476 3298 20528
rect 3528 20516 3556 20556
rect 4890 20544 4896 20556
rect 4948 20544 4954 20596
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 5721 20587 5779 20593
rect 5721 20584 5733 20587
rect 5592 20556 5733 20584
rect 5592 20544 5598 20556
rect 5721 20553 5733 20556
rect 5767 20553 5779 20587
rect 5721 20547 5779 20553
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 6512 20556 6561 20584
rect 6512 20544 6518 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 11054 20584 11060 20596
rect 11015 20556 11060 20584
rect 6549 20547 6607 20553
rect 11054 20544 11060 20556
rect 11112 20584 11118 20596
rect 11698 20584 11704 20596
rect 11112 20556 11704 20584
rect 11112 20544 11118 20556
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 12618 20544 12624 20596
rect 12676 20584 12682 20596
rect 12713 20587 12771 20593
rect 12713 20584 12725 20587
rect 12676 20556 12725 20584
rect 12676 20544 12682 20556
rect 12713 20553 12725 20556
rect 12759 20553 12771 20587
rect 12713 20547 12771 20553
rect 3344 20488 3556 20516
rect 3344 20457 3372 20488
rect 4706 20476 4712 20528
rect 4764 20476 4770 20528
rect 7466 20516 7472 20528
rect 6564 20488 7472 20516
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 2915 20420 3341 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3510 20448 3516 20460
rect 3471 20420 3516 20448
rect 3329 20411 3387 20417
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 6564 20457 6592 20488
rect 7466 20476 7472 20488
rect 7524 20476 7530 20528
rect 11606 20516 11612 20528
rect 9968 20488 11612 20516
rect 3973 20451 4031 20457
rect 3973 20448 3985 20451
rect 3936 20420 3985 20448
rect 3936 20408 3942 20420
rect 3973 20417 3985 20420
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20448 6791 20451
rect 6914 20448 6920 20460
rect 6779 20420 6920 20448
rect 6779 20417 6791 20420
rect 6733 20411 6791 20417
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20380 4307 20383
rect 5534 20380 5540 20392
rect 4295 20352 5540 20380
rect 4295 20349 4307 20352
rect 4249 20343 4307 20349
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 5350 20272 5356 20324
rect 5408 20312 5414 20324
rect 6564 20312 6592 20411
rect 6914 20408 6920 20420
rect 6972 20408 6978 20460
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 9861 20451 9919 20457
rect 9861 20448 9873 20451
rect 9640 20420 9873 20448
rect 9640 20408 9646 20420
rect 9861 20417 9873 20420
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 9674 20380 9680 20392
rect 5408 20284 6592 20312
rect 7484 20352 9680 20380
rect 5408 20272 5414 20284
rect 1765 20247 1823 20253
rect 1765 20213 1777 20247
rect 1811 20244 1823 20247
rect 4890 20244 4896 20256
rect 1811 20216 4896 20244
rect 1811 20213 1823 20216
rect 1765 20207 1823 20213
rect 4890 20204 4896 20216
rect 4948 20244 4954 20256
rect 7484 20244 7512 20352
rect 9674 20340 9680 20352
rect 9732 20340 9738 20392
rect 9968 20389 9996 20488
rect 11606 20476 11612 20488
rect 11664 20476 11670 20528
rect 11790 20516 11796 20528
rect 11751 20488 11796 20516
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 12728 20516 12756 20547
rect 14182 20544 14188 20596
rect 14240 20584 14246 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 14240 20556 14289 20584
rect 14240 20544 14246 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 16301 20587 16359 20593
rect 16301 20584 16313 20587
rect 16080 20556 16313 20584
rect 16080 20544 16086 20556
rect 16301 20553 16313 20556
rect 16347 20553 16359 20587
rect 16301 20547 16359 20553
rect 20073 20587 20131 20593
rect 20073 20553 20085 20587
rect 20119 20584 20131 20587
rect 20346 20584 20352 20596
rect 20119 20556 20352 20584
rect 20119 20553 20131 20556
rect 20073 20547 20131 20553
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 20533 20587 20591 20593
rect 20533 20553 20545 20587
rect 20579 20584 20591 20587
rect 21542 20584 21548 20596
rect 20579 20556 21548 20584
rect 20579 20553 20591 20556
rect 20533 20547 20591 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 23474 20584 23480 20596
rect 23435 20556 23480 20584
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 23658 20544 23664 20596
rect 23716 20544 23722 20596
rect 14645 20519 14703 20525
rect 14645 20516 14657 20519
rect 12728 20488 14657 20516
rect 14645 20485 14657 20488
rect 14691 20485 14703 20519
rect 14645 20479 14703 20485
rect 15933 20519 15991 20525
rect 15933 20485 15945 20519
rect 15979 20516 15991 20519
rect 16942 20516 16948 20528
rect 15979 20488 16948 20516
rect 15979 20485 15991 20488
rect 15933 20479 15991 20485
rect 16942 20476 16948 20488
rect 17000 20476 17006 20528
rect 17310 20516 17316 20528
rect 17271 20488 17316 20516
rect 17310 20476 17316 20488
rect 17368 20476 17374 20528
rect 22557 20519 22615 20525
rect 20180 20488 22232 20516
rect 18236 20460 18288 20466
rect 20180 20460 20208 20488
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 9953 20383 10011 20389
rect 9953 20349 9965 20383
rect 9999 20349 10011 20383
rect 10060 20380 10088 20411
rect 10134 20408 10140 20460
rect 10192 20448 10198 20460
rect 10265 20451 10323 20457
rect 10192 20420 10237 20448
rect 10192 20408 10198 20420
rect 10265 20417 10277 20451
rect 10311 20448 10323 20451
rect 10410 20448 10416 20460
rect 10311 20420 10416 20448
rect 10311 20417 10323 20420
rect 10265 20411 10323 20417
rect 10410 20408 10416 20420
rect 10468 20408 10474 20460
rect 11514 20408 11520 20460
rect 11572 20448 11578 20460
rect 13170 20448 13176 20460
rect 11572 20420 13176 20448
rect 11572 20408 11578 20420
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 13538 20448 13544 20460
rect 13495 20420 13544 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20448 14795 20451
rect 15562 20448 15568 20460
rect 14783 20420 15568 20448
rect 14783 20417 14795 20420
rect 14737 20411 14795 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15805 20451 15863 20457
rect 15805 20417 15817 20451
rect 15851 20448 15863 20451
rect 16022 20448 16028 20460
rect 15851 20417 15884 20448
rect 15983 20420 16028 20448
rect 15805 20411 15884 20417
rect 10060 20352 10364 20380
rect 9953 20343 10011 20349
rect 10336 20324 10364 20352
rect 13078 20340 13084 20392
rect 13136 20380 13142 20392
rect 13357 20383 13415 20389
rect 13357 20380 13369 20383
rect 13136 20352 13369 20380
rect 13136 20340 13142 20352
rect 13357 20349 13369 20352
rect 13403 20349 13415 20383
rect 14918 20380 14924 20392
rect 14879 20352 14924 20380
rect 13357 20343 13415 20349
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 8478 20312 8484 20324
rect 8128 20284 8484 20312
rect 8128 20256 8156 20284
rect 8478 20272 8484 20284
rect 8536 20272 8542 20324
rect 8754 20272 8760 20324
rect 8812 20312 8818 20324
rect 9309 20315 9367 20321
rect 9309 20312 9321 20315
rect 8812 20284 9321 20312
rect 8812 20272 8818 20284
rect 9309 20281 9321 20284
rect 9355 20281 9367 20315
rect 9309 20275 9367 20281
rect 4948 20216 7512 20244
rect 7561 20247 7619 20253
rect 4948 20204 4954 20216
rect 7561 20213 7573 20247
rect 7607 20244 7619 20247
rect 8110 20244 8116 20256
rect 7607 20216 8116 20244
rect 7607 20213 7619 20216
rect 7561 20207 7619 20213
rect 8110 20204 8116 20216
rect 8168 20204 8174 20256
rect 8294 20244 8300 20256
rect 8255 20216 8300 20244
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 8846 20244 8852 20256
rect 8807 20216 8852 20244
rect 8846 20204 8852 20216
rect 8904 20204 8910 20256
rect 9324 20244 9352 20275
rect 10318 20272 10324 20324
rect 10376 20272 10382 20324
rect 12158 20312 12164 20324
rect 11440 20284 12164 20312
rect 11440 20244 11468 20284
rect 12158 20272 12164 20284
rect 12216 20272 12222 20324
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 15672 20312 15700 20411
rect 15856 20380 15884 20411
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 16163 20451 16221 20457
rect 16163 20417 16175 20451
rect 16209 20448 16221 20451
rect 17586 20448 17592 20460
rect 16209 20420 17592 20448
rect 16209 20417 16221 20420
rect 16163 20411 16221 20417
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20448 18383 20451
rect 18414 20448 18420 20460
rect 18371 20420 18420 20448
rect 18371 20417 18383 20420
rect 18325 20411 18383 20417
rect 18414 20408 18420 20420
rect 18472 20448 18478 20460
rect 18782 20448 18788 20460
rect 18472 20420 18788 20448
rect 18472 20408 18478 20420
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 20162 20448 20168 20460
rect 20123 20420 20168 20448
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20680 20420 21005 20448
rect 20680 20408 20686 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 22204 20448 22232 20488
rect 22557 20485 22569 20519
rect 22603 20516 22615 20519
rect 23676 20516 23704 20544
rect 22603 20488 23704 20516
rect 22603 20485 22615 20488
rect 22557 20479 22615 20485
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 22204 20420 22661 20448
rect 20993 20411 21051 20417
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 23661 20451 23719 20457
rect 23661 20448 23673 20451
rect 22649 20411 22707 20417
rect 23032 20420 23673 20448
rect 18236 20402 18288 20408
rect 18046 20380 18052 20392
rect 15856 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 19242 20340 19248 20392
rect 19300 20380 19306 20392
rect 19889 20383 19947 20389
rect 19889 20380 19901 20383
rect 19300 20352 19901 20380
rect 19300 20340 19306 20352
rect 19889 20349 19901 20352
rect 19935 20349 19947 20383
rect 19889 20343 19947 20349
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 22373 20383 22431 20389
rect 22373 20380 22385 20383
rect 22152 20352 22385 20380
rect 22152 20340 22158 20352
rect 22373 20349 22385 20352
rect 22419 20349 22431 20383
rect 22373 20343 22431 20349
rect 18598 20312 18604 20324
rect 13863 20284 15700 20312
rect 15764 20284 18604 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 9324 20216 11468 20244
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 11572 20216 11897 20244
rect 11572 20204 11578 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 13630 20204 13636 20256
rect 13688 20244 13694 20256
rect 15764 20244 15792 20284
rect 18598 20272 18604 20284
rect 18656 20272 18662 20324
rect 21177 20315 21235 20321
rect 21177 20281 21189 20315
rect 21223 20312 21235 20315
rect 21726 20312 21732 20324
rect 21223 20284 21732 20312
rect 21223 20281 21235 20284
rect 21177 20275 21235 20281
rect 21726 20272 21732 20284
rect 21784 20272 21790 20324
rect 13688 20216 15792 20244
rect 13688 20204 13694 20216
rect 15930 20204 15936 20256
rect 15988 20244 15994 20256
rect 18138 20244 18144 20256
rect 15988 20216 18144 20244
rect 15988 20204 15994 20216
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18564 20216 18889 20244
rect 18564 20204 18570 20216
rect 18877 20213 18889 20216
rect 18923 20244 18935 20247
rect 19058 20244 19064 20256
rect 18923 20216 19064 20244
rect 18923 20213 18935 20216
rect 18877 20207 18935 20213
rect 19058 20204 19064 20216
rect 19116 20244 19122 20256
rect 21358 20244 21364 20256
rect 19116 20216 21364 20244
rect 19116 20204 19122 20216
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 22664 20244 22692 20411
rect 23032 20321 23060 20420
rect 23661 20417 23673 20420
rect 23707 20417 23719 20451
rect 23661 20411 23719 20417
rect 23017 20315 23075 20321
rect 23017 20281 23029 20315
rect 23063 20281 23075 20315
rect 23017 20275 23075 20281
rect 24121 20247 24179 20253
rect 24121 20244 24133 20247
rect 22664 20216 24133 20244
rect 24121 20213 24133 20216
rect 24167 20244 24179 20247
rect 24673 20247 24731 20253
rect 24673 20244 24685 20247
rect 24167 20216 24685 20244
rect 24167 20213 24179 20216
rect 24121 20207 24179 20213
rect 24673 20213 24685 20216
rect 24719 20213 24731 20247
rect 24673 20207 24731 20213
rect 1104 20154 27876 20176
rect 1104 20102 4296 20154
rect 4348 20102 4360 20154
rect 4412 20102 4424 20154
rect 4476 20102 4488 20154
rect 4540 20102 4552 20154
rect 4604 20102 10988 20154
rect 11040 20102 11052 20154
rect 11104 20102 11116 20154
rect 11168 20102 11180 20154
rect 11232 20102 11244 20154
rect 11296 20102 17680 20154
rect 17732 20102 17744 20154
rect 17796 20102 17808 20154
rect 17860 20102 17872 20154
rect 17924 20102 17936 20154
rect 17988 20102 24372 20154
rect 24424 20102 24436 20154
rect 24488 20102 24500 20154
rect 24552 20102 24564 20154
rect 24616 20102 24628 20154
rect 24680 20102 27876 20154
rect 1104 20080 27876 20102
rect 10594 20040 10600 20052
rect 10555 20012 10600 20040
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 13630 20040 13636 20052
rect 13591 20012 13636 20040
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 15562 20000 15568 20052
rect 15620 20040 15626 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15620 20012 15669 20040
rect 15620 20000 15626 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 5258 19932 5264 19984
rect 5316 19972 5322 19984
rect 6089 19975 6147 19981
rect 6089 19972 6101 19975
rect 5316 19944 6101 19972
rect 5316 19932 5322 19944
rect 6089 19941 6101 19944
rect 6135 19941 6147 19975
rect 12250 19972 12256 19984
rect 6089 19935 6147 19941
rect 9232 19944 12256 19972
rect 1486 19864 1492 19916
rect 1544 19904 1550 19916
rect 1581 19907 1639 19913
rect 1581 19904 1593 19907
rect 1544 19876 1593 19904
rect 1544 19864 1550 19876
rect 1581 19873 1593 19876
rect 1627 19873 1639 19907
rect 1581 19867 1639 19873
rect 6733 19907 6791 19913
rect 6733 19873 6745 19907
rect 6779 19904 6791 19907
rect 7282 19904 7288 19916
rect 6779 19876 7288 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 1854 19845 1860 19848
rect 1848 19836 1860 19845
rect 1815 19808 1860 19836
rect 1848 19799 1860 19808
rect 1854 19796 1860 19799
rect 1912 19796 1918 19848
rect 6914 19836 6920 19848
rect 5920 19808 6920 19836
rect 5920 19780 5948 19808
rect 6914 19796 6920 19808
rect 6972 19836 6978 19848
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 6972 19808 7389 19836
rect 6972 19796 6978 19808
rect 7377 19805 7389 19808
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 7466 19796 7472 19848
rect 7524 19836 7530 19848
rect 7561 19839 7619 19845
rect 7561 19836 7573 19839
rect 7524 19808 7573 19836
rect 7524 19796 7530 19808
rect 7561 19805 7573 19808
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 5537 19771 5595 19777
rect 5537 19768 5549 19771
rect 4448 19740 5549 19768
rect 2958 19700 2964 19712
rect 2919 19672 2964 19700
rect 2958 19660 2964 19672
rect 3016 19660 3022 19712
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 4448 19709 4476 19740
rect 5537 19737 5549 19740
rect 5583 19768 5595 19771
rect 5902 19768 5908 19780
rect 5583 19740 5908 19768
rect 5583 19737 5595 19740
rect 5537 19731 5595 19737
rect 5902 19728 5908 19740
rect 5960 19728 5966 19780
rect 6012 19740 6316 19768
rect 4433 19703 4491 19709
rect 4433 19700 4445 19703
rect 3568 19672 4445 19700
rect 3568 19660 3574 19672
rect 4433 19669 4445 19672
rect 4479 19669 4491 19703
rect 5074 19700 5080 19712
rect 5035 19672 5080 19700
rect 4433 19663 4491 19669
rect 5074 19660 5080 19672
rect 5132 19700 5138 19712
rect 6012 19700 6040 19740
rect 5132 19672 6040 19700
rect 6288 19700 6316 19740
rect 6362 19728 6368 19780
rect 6420 19768 6426 19780
rect 6549 19771 6607 19777
rect 6549 19768 6561 19771
rect 6420 19740 6561 19768
rect 6420 19728 6426 19740
rect 6549 19737 6561 19740
rect 6595 19737 6607 19771
rect 9232 19768 9260 19944
rect 12250 19932 12256 19944
rect 12308 19932 12314 19984
rect 11422 19864 11428 19916
rect 11480 19904 11486 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 11480 19876 12357 19904
rect 11480 19864 11486 19876
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12345 19867 12403 19873
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 9950 19836 9956 19848
rect 9355 19808 9956 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 10376 19808 10425 19836
rect 10376 19796 10382 19808
rect 10413 19805 10425 19808
rect 10459 19836 10471 19839
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 10459 19808 11069 19836
rect 10459 19805 10471 19808
rect 10413 19799 10471 19805
rect 11057 19805 11069 19808
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19836 12311 19839
rect 13078 19836 13084 19848
rect 12299 19808 13084 19836
rect 12299 19805 12311 19808
rect 12253 19799 12311 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 13722 19796 13728 19848
rect 13780 19836 13786 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 13780 19808 14289 19836
rect 13780 19796 13786 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 15672 19836 15700 20003
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16117 20043 16175 20049
rect 16117 20040 16129 20043
rect 16080 20012 16129 20040
rect 16080 20000 16086 20012
rect 16117 20009 16129 20012
rect 16163 20009 16175 20043
rect 16942 20040 16948 20052
rect 16903 20012 16948 20040
rect 16117 20003 16175 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17586 20000 17592 20052
rect 17644 20040 17650 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 17644 20012 17877 20040
rect 17644 20000 17650 20012
rect 17865 20009 17877 20012
rect 17911 20009 17923 20043
rect 17865 20003 17923 20009
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18104 20012 18521 20040
rect 18104 20000 18110 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 19794 20040 19800 20052
rect 19755 20012 19800 20040
rect 18509 20003 18567 20009
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 24854 20000 24860 20052
rect 24912 20040 24918 20052
rect 25133 20043 25191 20049
rect 25133 20040 25145 20043
rect 24912 20012 25145 20040
rect 24912 20000 24918 20012
rect 25133 20009 25145 20012
rect 25179 20009 25191 20043
rect 25133 20003 25191 20009
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17184 19944 18644 19972
rect 17184 19932 17190 19944
rect 16500 19876 18000 19904
rect 16500 19845 16528 19876
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 15672 19808 16497 19836
rect 14277 19799 14335 19805
rect 16485 19805 16497 19808
rect 16531 19805 16543 19839
rect 17402 19836 17408 19848
rect 16485 19799 16543 19805
rect 17052 19808 17408 19836
rect 6549 19731 6607 19737
rect 7392 19740 9260 19768
rect 10045 19771 10103 19777
rect 6457 19703 6515 19709
rect 6457 19700 6469 19703
rect 6288 19672 6469 19700
rect 5132 19660 5138 19672
rect 6457 19669 6469 19672
rect 6503 19700 6515 19703
rect 7392 19700 7420 19740
rect 10045 19737 10057 19771
rect 10091 19768 10103 19771
rect 10134 19768 10140 19780
rect 10091 19740 10140 19768
rect 10091 19737 10103 19740
rect 10045 19731 10103 19737
rect 10134 19728 10140 19740
rect 10192 19728 10198 19780
rect 11330 19768 11336 19780
rect 11291 19740 11336 19768
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 12158 19768 12164 19780
rect 12071 19740 12164 19768
rect 12158 19728 12164 19740
rect 12216 19768 12222 19780
rect 13446 19768 13452 19780
rect 12216 19740 13452 19768
rect 12216 19728 12222 19740
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 7558 19700 7564 19712
rect 6503 19672 7420 19700
rect 7519 19672 7564 19700
rect 6503 19669 6515 19672
rect 6457 19663 6515 19669
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 8570 19700 8576 19712
rect 8531 19672 8576 19700
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 9122 19700 9128 19712
rect 9083 19672 9128 19700
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 9582 19660 9588 19712
rect 9640 19700 9646 19712
rect 10229 19703 10287 19709
rect 10229 19700 10241 19703
rect 9640 19672 10241 19700
rect 9640 19660 9646 19672
rect 10229 19669 10241 19672
rect 10275 19669 10287 19703
rect 10229 19663 10287 19669
rect 10321 19703 10379 19709
rect 10321 19669 10333 19703
rect 10367 19700 10379 19703
rect 10410 19700 10416 19712
rect 10367 19672 10416 19700
rect 10367 19669 10379 19672
rect 10321 19663 10379 19669
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 11793 19703 11851 19709
rect 11793 19700 11805 19703
rect 10560 19672 11805 19700
rect 10560 19660 10566 19672
rect 11793 19669 11805 19672
rect 11839 19669 11851 19703
rect 11793 19663 11851 19669
rect 13081 19703 13139 19709
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 13262 19700 13268 19712
rect 13127 19672 13268 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 13262 19660 13268 19672
rect 13320 19660 13326 19712
rect 13556 19700 13584 19796
rect 14090 19728 14096 19780
rect 14148 19768 14154 19780
rect 14522 19771 14580 19777
rect 14522 19768 14534 19771
rect 14148 19740 14534 19768
rect 14148 19728 14154 19740
rect 14522 19737 14534 19740
rect 14568 19737 14580 19771
rect 14522 19731 14580 19737
rect 16301 19771 16359 19777
rect 16301 19737 16313 19771
rect 16347 19768 16359 19771
rect 17052 19768 17080 19808
rect 17402 19796 17408 19808
rect 17460 19836 17466 19848
rect 17972 19845 18000 19876
rect 18616 19845 18644 19944
rect 19242 19864 19248 19916
rect 19300 19904 19306 19916
rect 20349 19907 20407 19913
rect 20349 19904 20361 19907
rect 19300 19876 20361 19904
rect 19300 19864 19306 19876
rect 20349 19873 20361 19876
rect 20395 19873 20407 19907
rect 20349 19867 20407 19873
rect 23658 19864 23664 19916
rect 23716 19904 23722 19916
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 23716 19876 24685 19904
rect 23716 19864 23722 19876
rect 24673 19873 24685 19876
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 17460 19808 17785 19836
rect 17460 19796 17466 19808
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 19334 19836 19340 19848
rect 18647 19808 19340 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 16347 19740 17080 19768
rect 16347 19737 16359 19740
rect 16301 19731 16359 19737
rect 17126 19728 17132 19780
rect 17184 19768 17190 19780
rect 17313 19771 17371 19777
rect 17184 19740 17229 19768
rect 17184 19728 17190 19740
rect 17313 19737 17325 19771
rect 17359 19768 17371 19771
rect 18432 19768 18460 19799
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20806 19836 20812 19848
rect 20303 19808 20812 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 21450 19796 21456 19848
rect 21508 19836 21514 19848
rect 21910 19836 21916 19848
rect 21508 19808 21916 19836
rect 21508 19796 21514 19808
rect 21910 19796 21916 19808
rect 21968 19836 21974 19848
rect 22925 19839 22983 19845
rect 22925 19836 22937 19839
rect 21968 19808 22937 19836
rect 21968 19796 21974 19808
rect 22925 19805 22937 19808
rect 22971 19805 22983 19839
rect 23566 19836 23572 19848
rect 23527 19808 23572 19836
rect 22925 19799 22983 19805
rect 23566 19796 23572 19808
rect 23624 19796 23630 19848
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19836 24823 19839
rect 25866 19836 25872 19848
rect 24811 19808 25872 19836
rect 24811 19805 24823 19808
rect 24765 19799 24823 19805
rect 25866 19796 25872 19808
rect 25924 19836 25930 19848
rect 26329 19839 26387 19845
rect 26329 19836 26341 19839
rect 25924 19808 26341 19836
rect 25924 19796 25930 19808
rect 26329 19805 26341 19808
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 17359 19740 18460 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 15194 19700 15200 19712
rect 13556 19672 15200 19700
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 17328 19700 17356 19731
rect 18690 19728 18696 19780
rect 18748 19768 18754 19780
rect 20898 19768 20904 19780
rect 18748 19740 20904 19768
rect 18748 19728 18754 19740
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 22680 19771 22738 19777
rect 22680 19737 22692 19771
rect 22726 19768 22738 19771
rect 22726 19740 23428 19768
rect 22726 19737 22738 19740
rect 22680 19731 22738 19737
rect 15896 19672 17356 19700
rect 15896 19660 15902 19672
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19518 19700 19524 19712
rect 19392 19672 19524 19700
rect 19392 19660 19398 19672
rect 19518 19660 19524 19672
rect 19576 19700 19582 19712
rect 20165 19703 20223 19709
rect 20165 19700 20177 19703
rect 19576 19672 20177 19700
rect 19576 19660 19582 19672
rect 20165 19669 20177 19672
rect 20211 19700 20223 19703
rect 20530 19700 20536 19712
rect 20211 19672 20536 19700
rect 20211 19669 20223 19672
rect 20165 19663 20223 19669
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 20993 19703 21051 19709
rect 20993 19700 21005 19703
rect 20772 19672 21005 19700
rect 20772 19660 20778 19672
rect 20993 19669 21005 19672
rect 21039 19669 21051 19703
rect 20993 19663 21051 19669
rect 21545 19703 21603 19709
rect 21545 19669 21557 19703
rect 21591 19700 21603 19703
rect 22278 19700 22284 19712
rect 21591 19672 22284 19700
rect 21591 19669 21603 19672
rect 21545 19663 21603 19669
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 23400 19709 23428 19740
rect 23385 19703 23443 19709
rect 23385 19669 23397 19703
rect 23431 19669 23443 19703
rect 23385 19663 23443 19669
rect 25406 19660 25412 19712
rect 25464 19700 25470 19712
rect 26513 19703 26571 19709
rect 26513 19700 26525 19703
rect 25464 19672 26525 19700
rect 25464 19660 25470 19672
rect 26513 19669 26525 19672
rect 26559 19669 26571 19703
rect 26513 19663 26571 19669
rect 1104 19610 28032 19632
rect 1104 19558 7642 19610
rect 7694 19558 7706 19610
rect 7758 19558 7770 19610
rect 7822 19558 7834 19610
rect 7886 19558 7898 19610
rect 7950 19558 14334 19610
rect 14386 19558 14398 19610
rect 14450 19558 14462 19610
rect 14514 19558 14526 19610
rect 14578 19558 14590 19610
rect 14642 19558 21026 19610
rect 21078 19558 21090 19610
rect 21142 19558 21154 19610
rect 21206 19558 21218 19610
rect 21270 19558 21282 19610
rect 21334 19558 27718 19610
rect 27770 19558 27782 19610
rect 27834 19558 27846 19610
rect 27898 19558 27910 19610
rect 27962 19558 27974 19610
rect 28026 19558 28032 19610
rect 1104 19536 28032 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 3326 19496 3332 19508
rect 1627 19468 3332 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 3973 19499 4031 19505
rect 3973 19465 3985 19499
rect 4019 19496 4031 19499
rect 4798 19496 4804 19508
rect 4019 19468 4804 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 4798 19456 4804 19468
rect 4856 19456 4862 19508
rect 5902 19496 5908 19508
rect 5863 19468 5908 19496
rect 5902 19456 5908 19468
rect 5960 19456 5966 19508
rect 7098 19496 7104 19508
rect 7059 19468 7104 19496
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 8478 19456 8484 19508
rect 8536 19496 8542 19508
rect 9585 19499 9643 19505
rect 8536 19468 9536 19496
rect 8536 19456 8542 19468
rect 2716 19431 2774 19437
rect 2716 19397 2728 19431
rect 2762 19428 2774 19431
rect 2958 19428 2964 19440
rect 2762 19400 2964 19428
rect 2762 19397 2774 19400
rect 2716 19391 2774 19397
rect 2958 19388 2964 19400
rect 3016 19388 3022 19440
rect 4172 19400 7420 19428
rect 4172 19369 4200 19400
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19329 4215 19363
rect 5258 19360 5264 19372
rect 5219 19332 5264 19360
rect 4157 19323 4215 19329
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 7006 19360 7012 19372
rect 6967 19332 7012 19360
rect 7006 19320 7012 19332
rect 7064 19320 7070 19372
rect 7392 19304 7420 19400
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 7616 19400 8602 19428
rect 7616 19388 7622 19400
rect 9508 19360 9536 19468
rect 9585 19465 9597 19499
rect 9631 19465 9643 19499
rect 9585 19459 9643 19465
rect 9600 19428 9628 19459
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 10045 19499 10103 19505
rect 10045 19496 10057 19499
rect 10008 19468 10057 19496
rect 10008 19456 10014 19468
rect 10045 19465 10057 19468
rect 10091 19465 10103 19499
rect 10045 19459 10103 19465
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11480 19468 11713 19496
rect 11480 19456 11486 19468
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 12529 19499 12587 19505
rect 12529 19465 12541 19499
rect 12575 19496 12587 19499
rect 16850 19496 16856 19508
rect 12575 19468 16856 19496
rect 12575 19465 12587 19468
rect 12529 19459 12587 19465
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 18601 19499 18659 19505
rect 18601 19465 18613 19499
rect 18647 19496 18659 19499
rect 18690 19496 18696 19508
rect 18647 19468 18696 19496
rect 18647 19465 18659 19468
rect 18601 19459 18659 19465
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 20622 19496 20628 19508
rect 20583 19468 20628 19496
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 22278 19496 22284 19508
rect 22239 19468 22284 19496
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 22741 19499 22799 19505
rect 22741 19465 22753 19499
rect 22787 19496 22799 19499
rect 23566 19496 23572 19508
rect 22787 19468 23572 19496
rect 22787 19465 22799 19468
rect 22741 19459 22799 19465
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 25866 19496 25872 19508
rect 25827 19468 25872 19496
rect 25866 19456 25872 19468
rect 25924 19456 25930 19508
rect 10134 19428 10140 19440
rect 9600 19400 10140 19428
rect 10134 19388 10140 19400
rect 10192 19428 10198 19440
rect 10505 19431 10563 19437
rect 10505 19428 10517 19431
rect 10192 19400 10517 19428
rect 10192 19388 10198 19400
rect 10505 19397 10517 19400
rect 10551 19397 10563 19431
rect 12618 19428 12624 19440
rect 10505 19391 10563 19397
rect 11716 19400 12624 19428
rect 10413 19363 10471 19369
rect 10413 19360 10425 19363
rect 9508 19332 10425 19360
rect 10413 19329 10425 19332
rect 10459 19360 10471 19363
rect 11514 19360 11520 19372
rect 10459 19332 11520 19360
rect 10459 19329 10471 19332
rect 10413 19323 10471 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11716 19369 11744 19400
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 15838 19428 15844 19440
rect 13228 19400 15700 19428
rect 15799 19400 15844 19428
rect 13228 19388 13234 19400
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 12066 19360 12072 19372
rect 11931 19332 12072 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19360 13047 19363
rect 14182 19360 14188 19372
rect 13035 19332 14188 19360
rect 13035 19329 13047 19332
rect 12989 19323 13047 19329
rect 2958 19292 2964 19304
rect 2919 19264 2964 19292
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 7282 19292 7288 19304
rect 7243 19264 7288 19292
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 7834 19292 7840 19304
rect 7432 19264 7840 19292
rect 7432 19252 7438 19264
rect 7834 19252 7840 19264
rect 7892 19252 7898 19304
rect 8113 19295 8171 19301
rect 8113 19261 8125 19295
rect 8159 19292 8171 19295
rect 9122 19292 9128 19304
rect 8159 19264 9128 19292
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 11422 19292 11428 19304
rect 10735 19264 11428 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 11422 19252 11428 19264
rect 11480 19252 11486 19304
rect 12360 19224 12388 19323
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 15672 19360 15700 19400
rect 15838 19388 15844 19400
rect 15896 19388 15902 19440
rect 15930 19388 15936 19440
rect 15988 19428 15994 19440
rect 19334 19428 19340 19440
rect 15988 19400 16033 19428
rect 16224 19400 19340 19428
rect 15988 19388 15994 19400
rect 16224 19360 16252 19400
rect 19334 19388 19340 19400
rect 19392 19388 19398 19440
rect 19521 19431 19579 19437
rect 19521 19397 19533 19431
rect 19567 19428 19579 19431
rect 20806 19428 20812 19440
rect 19567 19400 20812 19428
rect 19567 19397 19579 19400
rect 19521 19391 19579 19397
rect 20806 19388 20812 19400
rect 20864 19388 20870 19440
rect 21634 19428 21640 19440
rect 21192 19400 21640 19428
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 15672 19332 16252 19360
rect 16316 19332 17049 19360
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15436 19264 15669 19292
rect 15436 19252 15442 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 15657 19255 15715 19261
rect 14277 19227 14335 19233
rect 14277 19224 14289 19227
rect 4816 19196 7972 19224
rect 12360 19196 14289 19224
rect 4816 19168 4844 19196
rect 4709 19159 4767 19165
rect 4709 19125 4721 19159
rect 4755 19156 4767 19159
rect 4798 19156 4804 19168
rect 4755 19128 4804 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5445 19159 5503 19165
rect 5445 19125 5457 19159
rect 5491 19156 5503 19159
rect 5718 19156 5724 19168
rect 5491 19128 5724 19156
rect 5491 19125 5503 19128
rect 5445 19119 5503 19125
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6730 19156 6736 19168
rect 6687 19128 6736 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 7944 19156 7972 19196
rect 14277 19193 14289 19196
rect 14323 19193 14335 19227
rect 15672 19224 15700 19255
rect 16316 19233 16344 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 17037 19323 17095 19329
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19116 19332 19441 19360
rect 19116 19320 19122 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 20438 19360 20444 19372
rect 19429 19323 19487 19329
rect 19628 19334 19840 19360
rect 19628 19332 19932 19334
rect 20399 19332 20444 19360
rect 18230 19292 18236 19304
rect 18191 19264 18236 19292
rect 18230 19252 18236 19264
rect 18288 19292 18294 19304
rect 19628 19292 19656 19332
rect 19812 19306 19932 19332
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20588 19332 20852 19360
rect 20588 19320 20594 19332
rect 18288 19264 19656 19292
rect 19705 19295 19763 19301
rect 18288 19252 18294 19264
rect 19705 19261 19717 19295
rect 19751 19261 19763 19295
rect 19904 19292 19932 19306
rect 20257 19295 20315 19301
rect 20257 19292 20269 19295
rect 19904 19264 20269 19292
rect 19705 19255 19763 19261
rect 20257 19261 20269 19264
rect 20303 19261 20315 19295
rect 20824 19292 20852 19332
rect 20898 19320 20904 19372
rect 20956 19360 20962 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20956 19332 21097 19360
rect 20956 19320 20962 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 21192 19292 21220 19400
rect 21634 19388 21640 19400
rect 21692 19428 21698 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 21692 19400 22385 19428
rect 21692 19388 21698 19400
rect 22373 19397 22385 19400
rect 22419 19428 22431 19431
rect 22419 19400 23612 19428
rect 22419 19397 22431 19400
rect 22373 19391 22431 19397
rect 23584 19372 23612 19400
rect 23474 19360 23480 19372
rect 23435 19332 23480 19360
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 23566 19320 23572 19372
rect 23624 19320 23630 19372
rect 23661 19363 23719 19369
rect 23661 19329 23673 19363
rect 23707 19360 23719 19363
rect 24121 19363 24179 19369
rect 24121 19360 24133 19363
rect 23707 19332 24133 19360
rect 23707 19329 23719 19332
rect 23661 19323 23719 19329
rect 24121 19329 24133 19332
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 25498 19320 25504 19372
rect 25556 19320 25562 19372
rect 26326 19360 26332 19372
rect 26287 19332 26332 19360
rect 26326 19320 26332 19332
rect 26384 19320 26390 19372
rect 20824 19264 21220 19292
rect 20257 19255 20315 19261
rect 16301 19227 16359 19233
rect 15672 19196 16252 19224
rect 14277 19187 14335 19193
rect 9214 19156 9220 19168
rect 7944 19128 9220 19156
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 16114 19156 16120 19168
rect 12216 19128 16120 19156
rect 12216 19116 12222 19128
rect 16114 19116 16120 19128
rect 16172 19116 16178 19168
rect 16224 19156 16252 19196
rect 16301 19193 16313 19227
rect 16347 19193 16359 19227
rect 19242 19224 19248 19236
rect 16301 19187 16359 19193
rect 16684 19196 19248 19224
rect 16684 19156 16712 19196
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 19610 19184 19616 19236
rect 19668 19224 19674 19236
rect 19720 19224 19748 19255
rect 21818 19252 21824 19304
rect 21876 19292 21882 19304
rect 22094 19292 22100 19304
rect 21876 19264 22100 19292
rect 21876 19252 21882 19264
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 24397 19295 24455 19301
rect 24397 19261 24409 19295
rect 24443 19292 24455 19295
rect 25406 19292 25412 19304
rect 24443 19264 25412 19292
rect 24443 19261 24455 19264
rect 24397 19255 24455 19261
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 19668 19196 19748 19224
rect 19668 19184 19674 19196
rect 16850 19156 16856 19168
rect 16224 19128 16712 19156
rect 16811 19128 16856 19156
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17402 19116 17408 19168
rect 17460 19156 17466 19168
rect 17497 19159 17555 19165
rect 17497 19156 17509 19159
rect 17460 19128 17509 19156
rect 17460 19116 17466 19128
rect 17497 19125 17509 19128
rect 17543 19125 17555 19159
rect 17497 19119 17555 19125
rect 18690 19116 18696 19168
rect 18748 19156 18754 19168
rect 19061 19159 19119 19165
rect 19061 19156 19073 19159
rect 18748 19128 19073 19156
rect 18748 19116 18754 19128
rect 19061 19125 19073 19128
rect 19107 19125 19119 19159
rect 19061 19119 19119 19125
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21542 19156 21548 19168
rect 21315 19128 21548 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 26513 19159 26571 19165
rect 26513 19125 26525 19159
rect 26559 19156 26571 19159
rect 27062 19156 27068 19168
rect 26559 19128 27068 19156
rect 26559 19125 26571 19128
rect 26513 19119 26571 19125
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 1104 19066 27876 19088
rect 1104 19014 4296 19066
rect 4348 19014 4360 19066
rect 4412 19014 4424 19066
rect 4476 19014 4488 19066
rect 4540 19014 4552 19066
rect 4604 19014 10988 19066
rect 11040 19014 11052 19066
rect 11104 19014 11116 19066
rect 11168 19014 11180 19066
rect 11232 19014 11244 19066
rect 11296 19014 17680 19066
rect 17732 19014 17744 19066
rect 17796 19014 17808 19066
rect 17860 19014 17872 19066
rect 17924 19014 17936 19066
rect 17988 19014 24372 19066
rect 24424 19014 24436 19066
rect 24488 19014 24500 19066
rect 24552 19014 24564 19066
rect 24616 19014 24628 19066
rect 24680 19014 27876 19066
rect 1104 18992 27876 19014
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 7098 18952 7104 18964
rect 5031 18924 7104 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 9861 18955 9919 18961
rect 9861 18921 9873 18955
rect 9907 18952 9919 18955
rect 10318 18952 10324 18964
rect 9907 18924 10324 18952
rect 9907 18921 9919 18924
rect 9861 18915 9919 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 13078 18952 13084 18964
rect 13039 18924 13084 18952
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 15565 18955 15623 18961
rect 15565 18921 15577 18955
rect 15611 18952 15623 18955
rect 15838 18952 15844 18964
rect 15611 18924 15844 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 18414 18952 18420 18964
rect 15948 18924 18420 18952
rect 7374 18884 7380 18896
rect 6748 18856 7380 18884
rect 6748 18825 6776 18856
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 15102 18884 15108 18896
rect 14476 18856 15108 18884
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18785 6791 18819
rect 6733 18779 6791 18785
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 7340 18788 8493 18816
rect 7340 18776 7346 18788
rect 8481 18785 8493 18788
rect 8527 18816 8539 18819
rect 11422 18816 11428 18828
rect 8527 18788 9812 18816
rect 8527 18785 8539 18788
rect 8481 18779 8539 18785
rect 4154 18748 4160 18760
rect 2240 18720 4160 18748
rect 2240 18624 2268 18720
rect 4154 18708 4160 18720
rect 4212 18748 4218 18760
rect 4249 18751 4307 18757
rect 4249 18748 4261 18751
rect 4212 18720 4261 18748
rect 4212 18708 4218 18720
rect 4249 18717 4261 18720
rect 4295 18717 4307 18751
rect 4249 18711 4307 18717
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18748 4491 18751
rect 4706 18748 4712 18760
rect 4479 18720 4712 18748
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 8202 18748 8208 18760
rect 7239 18720 7880 18748
rect 8163 18720 8208 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 4341 18683 4399 18689
rect 4341 18649 4353 18683
rect 4387 18680 4399 18683
rect 6457 18683 6515 18689
rect 4387 18652 5290 18680
rect 4387 18649 4399 18652
rect 4341 18643 4399 18649
rect 6457 18649 6469 18683
rect 6503 18680 6515 18683
rect 6546 18680 6552 18692
rect 6503 18652 6552 18680
rect 6503 18649 6515 18652
rect 6457 18643 6515 18649
rect 6546 18640 6552 18652
rect 6604 18640 6610 18692
rect 1765 18615 1823 18621
rect 1765 18581 1777 18615
rect 1811 18612 1823 18615
rect 2222 18612 2228 18624
rect 1811 18584 2228 18612
rect 1811 18581 1823 18584
rect 1765 18575 1823 18581
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 2317 18615 2375 18621
rect 2317 18581 2329 18615
rect 2363 18612 2375 18615
rect 2590 18612 2596 18624
rect 2363 18584 2596 18612
rect 2363 18581 2375 18584
rect 2317 18575 2375 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 2869 18615 2927 18621
rect 2869 18581 2881 18615
rect 2915 18612 2927 18615
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 2915 18584 3433 18612
rect 2915 18581 2927 18584
rect 2869 18575 2927 18581
rect 3421 18581 3433 18584
rect 3467 18612 3479 18615
rect 3510 18612 3516 18624
rect 3467 18584 3516 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 3510 18572 3516 18584
rect 3568 18572 3574 18624
rect 7374 18612 7380 18624
rect 7335 18584 7380 18612
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 7852 18621 7880 18720
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 9674 18748 9680 18760
rect 9447 18720 9680 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 9784 18748 9812 18788
rect 11164 18788 11428 18816
rect 11164 18748 11192 18788
rect 11422 18776 11428 18788
rect 11480 18776 11486 18828
rect 11698 18816 11704 18828
rect 11659 18788 11704 18816
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 14476 18816 14504 18856
rect 15102 18844 15108 18856
rect 15160 18884 15166 18896
rect 15948 18884 15976 18924
rect 18414 18912 18420 18924
rect 18472 18912 18478 18964
rect 20162 18952 20168 18964
rect 19444 18924 20168 18952
rect 15160 18856 15976 18884
rect 15160 18844 15166 18856
rect 17402 18844 17408 18896
rect 17460 18884 17466 18896
rect 19444 18884 19472 18924
rect 20162 18912 20168 18924
rect 20220 18912 20226 18964
rect 20806 18952 20812 18964
rect 20767 18924 20812 18952
rect 20806 18912 20812 18924
rect 20864 18912 20870 18964
rect 17460 18856 19472 18884
rect 23753 18887 23811 18893
rect 17460 18844 17466 18856
rect 23753 18853 23765 18887
rect 23799 18853 23811 18887
rect 23753 18847 23811 18853
rect 14384 18788 14504 18816
rect 14645 18819 14703 18825
rect 9784 18720 11192 18748
rect 11241 18751 11299 18757
rect 11241 18717 11253 18751
rect 11287 18748 11299 18751
rect 13725 18751 13783 18757
rect 11287 18720 11652 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 8297 18683 8355 18689
rect 8297 18649 8309 18683
rect 8343 18680 8355 18683
rect 9582 18680 9588 18692
rect 8343 18652 9588 18680
rect 8343 18649 8355 18652
rect 8297 18643 8355 18649
rect 9582 18640 9588 18652
rect 9640 18640 9646 18692
rect 10996 18683 11054 18689
rect 10996 18649 11008 18683
rect 11042 18680 11054 18683
rect 11330 18680 11336 18692
rect 11042 18652 11336 18680
rect 11042 18649 11054 18652
rect 10996 18643 11054 18649
rect 11330 18640 11336 18652
rect 11388 18640 11394 18692
rect 7837 18615 7895 18621
rect 7837 18581 7849 18615
rect 7883 18581 7895 18615
rect 9214 18612 9220 18624
rect 9175 18584 9220 18612
rect 7837 18575 7895 18581
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 11624 18612 11652 18720
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 13998 18748 14004 18760
rect 13771 18720 14004 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 14384 18757 14412 18788
rect 14645 18785 14657 18819
rect 14691 18816 14703 18819
rect 14918 18816 14924 18828
rect 14691 18788 14924 18816
rect 14691 18785 14703 18788
rect 14645 18779 14703 18785
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 16960 18788 19441 18816
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18717 14427 18751
rect 14369 18711 14427 18717
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 16689 18751 16747 18757
rect 16689 18717 16701 18751
rect 16735 18748 16747 18751
rect 16850 18748 16856 18760
rect 16735 18720 16856 18748
rect 16735 18717 16747 18720
rect 16689 18711 16747 18717
rect 11790 18640 11796 18692
rect 11848 18680 11854 18692
rect 11946 18683 12004 18689
rect 11946 18680 11958 18683
rect 11848 18652 11958 18680
rect 11848 18640 11854 18652
rect 11946 18649 11958 18652
rect 11992 18649 12004 18683
rect 11946 18643 12004 18649
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 14476 18680 14504 18711
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 16960 18757 16988 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 21542 18816 21548 18828
rect 21503 18788 21548 18816
rect 19429 18779 19487 18785
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18816 21879 18819
rect 23768 18816 23796 18847
rect 21867 18788 23796 18816
rect 21867 18785 21879 18788
rect 21821 18779 21879 18785
rect 25498 18776 25504 18828
rect 25556 18816 25562 18828
rect 25593 18819 25651 18825
rect 25593 18816 25605 18819
rect 25556 18788 25605 18816
rect 25556 18776 25562 18788
rect 25593 18785 25605 18788
rect 25639 18785 25651 18819
rect 25593 18779 25651 18785
rect 25320 18760 25372 18766
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 12676 18652 14504 18680
rect 12676 18640 12682 18652
rect 16390 18640 16396 18692
rect 16448 18680 16454 18692
rect 16960 18680 16988 18711
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17552 18720 17877 18748
rect 17552 18708 17558 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 18690 18748 18696 18760
rect 18651 18720 18696 18748
rect 17865 18711 17923 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 23474 18748 23480 18760
rect 23308 18720 23480 18748
rect 19674 18683 19732 18689
rect 19674 18680 19686 18683
rect 16448 18652 16988 18680
rect 18892 18652 19686 18680
rect 16448 18640 16454 18652
rect 12158 18612 12164 18624
rect 11624 18584 12164 18612
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 13630 18612 13636 18624
rect 13591 18584 13636 18612
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 18049 18615 18107 18621
rect 18049 18581 18061 18615
rect 18095 18612 18107 18615
rect 18414 18612 18420 18624
rect 18095 18584 18420 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18892 18621 18920 18652
rect 19674 18649 19686 18652
rect 19720 18649 19732 18683
rect 19674 18643 19732 18649
rect 22830 18640 22836 18692
rect 22888 18640 22894 18692
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18581 18935 18615
rect 18877 18575 18935 18581
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 23308 18621 23336 18720
rect 23474 18708 23480 18720
rect 23532 18748 23538 18760
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23532 18720 23765 18748
rect 23532 18708 23538 18720
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 24670 18748 24676 18760
rect 24631 18720 24676 18748
rect 23753 18711 23811 18717
rect 24670 18708 24676 18720
rect 24728 18708 24734 18760
rect 26421 18751 26479 18757
rect 26421 18717 26433 18751
rect 26467 18748 26479 18751
rect 26602 18748 26608 18760
rect 26467 18720 26608 18748
rect 26467 18717 26479 18720
rect 26421 18711 26479 18717
rect 26602 18708 26608 18720
rect 26660 18748 26666 18760
rect 26881 18751 26939 18757
rect 26881 18748 26893 18751
rect 26660 18720 26893 18748
rect 26660 18708 26666 18720
rect 26881 18717 26893 18720
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 25320 18702 25372 18708
rect 25774 18640 25780 18692
rect 25832 18680 25838 18692
rect 26145 18683 26203 18689
rect 26145 18680 26157 18683
rect 25832 18652 26157 18680
rect 25832 18640 25838 18652
rect 26145 18649 26157 18652
rect 26191 18649 26203 18683
rect 26145 18643 26203 18649
rect 27157 18683 27215 18689
rect 27157 18649 27169 18683
rect 27203 18680 27215 18683
rect 27338 18680 27344 18692
rect 27203 18652 27344 18680
rect 27203 18649 27215 18652
rect 27157 18643 27215 18649
rect 27338 18640 27344 18652
rect 27396 18640 27402 18692
rect 23293 18615 23351 18621
rect 23293 18612 23305 18615
rect 22152 18584 23305 18612
rect 22152 18572 22158 18584
rect 23293 18581 23305 18584
rect 23339 18581 23351 18615
rect 23293 18575 23351 18581
rect 1104 18522 28032 18544
rect 1104 18470 7642 18522
rect 7694 18470 7706 18522
rect 7758 18470 7770 18522
rect 7822 18470 7834 18522
rect 7886 18470 7898 18522
rect 7950 18470 14334 18522
rect 14386 18470 14398 18522
rect 14450 18470 14462 18522
rect 14514 18470 14526 18522
rect 14578 18470 14590 18522
rect 14642 18470 21026 18522
rect 21078 18470 21090 18522
rect 21142 18470 21154 18522
rect 21206 18470 21218 18522
rect 21270 18470 21282 18522
rect 21334 18470 27718 18522
rect 27770 18470 27782 18522
rect 27834 18470 27846 18522
rect 27898 18470 27910 18522
rect 27962 18470 27974 18522
rect 28026 18470 28032 18522
rect 1104 18448 28032 18470
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 6362 18408 6368 18420
rect 4295 18380 6368 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 9125 18411 9183 18417
rect 9125 18377 9137 18411
rect 9171 18408 9183 18411
rect 9582 18408 9588 18420
rect 9171 18380 9588 18408
rect 9171 18377 9183 18380
rect 9125 18371 9183 18377
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10410 18408 10416 18420
rect 9732 18380 10416 18408
rect 9732 18368 9738 18380
rect 10410 18368 10416 18380
rect 10468 18408 10474 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10468 18380 10977 18408
rect 10468 18368 10474 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 10965 18371 11023 18377
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 13722 18408 13728 18420
rect 12575 18380 13728 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 13722 18368 13728 18380
rect 13780 18408 13786 18420
rect 13780 18380 14136 18408
rect 13780 18368 13786 18380
rect 2590 18300 2596 18352
rect 2648 18300 2654 18352
rect 5718 18340 5724 18352
rect 5679 18312 5724 18340
rect 5718 18300 5724 18312
rect 5776 18300 5782 18352
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 7432 18312 7665 18340
rect 7432 18300 7438 18312
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 7653 18303 7711 18309
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 9830 18343 9888 18349
rect 9830 18340 9842 18343
rect 9272 18312 9842 18340
rect 9272 18300 9278 18312
rect 9830 18309 9842 18312
rect 9876 18309 9888 18343
rect 9830 18303 9888 18309
rect 11977 18343 12035 18349
rect 11977 18309 11989 18343
rect 12023 18340 12035 18343
rect 13173 18343 13231 18349
rect 13173 18340 13185 18343
rect 12023 18312 13185 18340
rect 12023 18309 12035 18312
rect 11977 18303 12035 18309
rect 13173 18309 13185 18312
rect 13219 18309 13231 18343
rect 14108 18340 14136 18380
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 14461 18411 14519 18417
rect 14461 18408 14473 18411
rect 14240 18380 14473 18408
rect 14240 18368 14246 18380
rect 14461 18377 14473 18380
rect 14507 18377 14519 18411
rect 14461 18371 14519 18377
rect 20165 18411 20223 18417
rect 20165 18377 20177 18411
rect 20211 18408 20223 18411
rect 20622 18408 20628 18420
rect 20211 18380 20628 18408
rect 20211 18377 20223 18380
rect 20165 18371 20223 18377
rect 20622 18368 20628 18380
rect 20680 18408 20686 18420
rect 20898 18408 20904 18420
rect 20680 18380 20904 18408
rect 20680 18368 20686 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 23566 18408 23572 18420
rect 23527 18380 23572 18408
rect 23566 18368 23572 18380
rect 23624 18408 23630 18420
rect 24121 18411 24179 18417
rect 24121 18408 24133 18411
rect 23624 18380 24133 18408
rect 23624 18368 23630 18380
rect 24121 18377 24133 18380
rect 24167 18377 24179 18411
rect 24121 18371 24179 18377
rect 16390 18340 16396 18352
rect 14108 18312 16396 18340
rect 13173 18303 13231 18309
rect 16390 18300 16396 18312
rect 16448 18300 16454 18352
rect 19334 18300 19340 18352
rect 19392 18300 19398 18352
rect 22830 18340 22836 18352
rect 22791 18312 22836 18340
rect 22830 18300 22836 18312
rect 22888 18300 22894 18352
rect 1946 18077 1952 18080
rect 1903 18071 1952 18077
rect 1903 18037 1915 18071
rect 1949 18037 1952 18071
rect 1903 18031 1952 18037
rect 1946 18028 1952 18031
rect 2004 18028 2010 18080
rect 2608 18068 2636 18300
rect 3326 18272 3332 18284
rect 3287 18244 3332 18272
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 4614 18232 4620 18284
rect 4672 18232 4678 18284
rect 6730 18272 6736 18284
rect 6691 18244 6736 18272
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 12158 18272 12164 18284
rect 12119 18244 12164 18272
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18272 12771 18275
rect 13630 18272 13636 18284
rect 12759 18244 13636 18272
rect 12759 18241 12771 18244
rect 12713 18235 12771 18241
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 15930 18272 15936 18284
rect 15703 18244 15936 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18241 17187 18275
rect 17129 18235 17187 18241
rect 3697 18207 3755 18213
rect 3697 18173 3709 18207
rect 3743 18204 3755 18207
rect 3970 18204 3976 18216
rect 3743 18176 3976 18204
rect 3743 18173 3755 18176
rect 3697 18167 3755 18173
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 5994 18204 6000 18216
rect 5907 18176 6000 18204
rect 5994 18164 6000 18176
rect 6052 18204 6058 18216
rect 7377 18207 7435 18213
rect 7377 18204 7389 18207
rect 6052 18176 7389 18204
rect 6052 18164 6058 18176
rect 7377 18173 7389 18176
rect 7423 18204 7435 18207
rect 8018 18204 8024 18216
rect 7423 18176 8024 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 8018 18164 8024 18176
rect 8076 18204 8082 18216
rect 8662 18204 8668 18216
rect 8076 18176 8668 18204
rect 8076 18164 8082 18176
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 9582 18204 9588 18216
rect 9543 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 12420 18207 12478 18213
rect 12420 18173 12432 18207
rect 12466 18204 12478 18207
rect 12526 18204 12532 18216
rect 12466 18176 12532 18204
rect 12466 18173 12478 18176
rect 12420 18167 12478 18173
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12676 18176 12721 18204
rect 12676 18164 12682 18176
rect 15194 18164 15200 18216
rect 15252 18204 15258 18216
rect 16132 18204 16160 18235
rect 15252 18176 16160 18204
rect 17144 18204 17172 18235
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 17681 18275 17739 18281
rect 17681 18272 17693 18275
rect 17552 18244 17693 18272
rect 17552 18232 17558 18244
rect 17681 18241 17693 18244
rect 17727 18241 17739 18275
rect 18414 18272 18420 18284
rect 18375 18244 18420 18272
rect 17681 18235 17739 18241
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 20898 18272 20904 18284
rect 20859 18244 20904 18272
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 21910 18232 21916 18284
rect 21968 18272 21974 18284
rect 22097 18275 22155 18281
rect 22097 18272 22109 18275
rect 21968 18244 22109 18272
rect 21968 18232 21974 18244
rect 22097 18241 22109 18244
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 25314 18232 25320 18284
rect 25372 18272 25378 18284
rect 25372 18244 25714 18272
rect 25372 18232 25378 18244
rect 17586 18204 17592 18216
rect 17144 18176 17592 18204
rect 15252 18164 15258 18176
rect 17586 18164 17592 18176
rect 17644 18164 17650 18216
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18204 18751 18207
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 18739 18176 20637 18204
rect 18739 18173 18751 18176
rect 18693 18167 18751 18173
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 25041 18207 25099 18213
rect 25041 18173 25053 18207
rect 25087 18204 25099 18207
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25087 18176 25789 18204
rect 25087 18173 25099 18176
rect 25041 18167 25099 18173
rect 25777 18173 25789 18176
rect 25823 18204 25835 18207
rect 26510 18204 26516 18216
rect 25823 18176 26234 18204
rect 26471 18176 26516 18204
rect 25823 18173 25835 18176
rect 25777 18167 25835 18173
rect 26206 18148 26234 18176
rect 26510 18164 26516 18176
rect 26568 18164 26574 18216
rect 13814 18096 13820 18148
rect 13872 18136 13878 18148
rect 16209 18139 16267 18145
rect 16209 18136 16221 18139
rect 13872 18108 16221 18136
rect 13872 18096 13878 18108
rect 16209 18105 16221 18108
rect 16255 18105 16267 18139
rect 26206 18108 26240 18148
rect 16209 18099 16267 18105
rect 26234 18096 26240 18108
rect 26292 18096 26298 18148
rect 9490 18068 9496 18080
rect 2608 18040 9496 18068
rect 9490 18028 9496 18040
rect 9548 18068 9554 18080
rect 9766 18068 9772 18080
rect 9548 18040 9772 18068
rect 9548 18028 9554 18040
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 14792 18040 15485 18068
rect 14792 18028 14798 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 16942 18068 16948 18080
rect 16903 18040 16948 18068
rect 15473 18031 15531 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17034 18028 17040 18080
rect 17092 18068 17098 18080
rect 17681 18071 17739 18077
rect 17681 18068 17693 18071
rect 17092 18040 17693 18068
rect 17092 18028 17098 18040
rect 17681 18037 17693 18040
rect 17727 18037 17739 18071
rect 17681 18031 17739 18037
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21361 18071 21419 18077
rect 21361 18068 21373 18071
rect 20956 18040 21373 18068
rect 20956 18028 20962 18040
rect 21361 18037 21373 18040
rect 21407 18037 21419 18071
rect 21361 18031 21419 18037
rect 1104 17978 27876 18000
rect 1104 17926 4296 17978
rect 4348 17926 4360 17978
rect 4412 17926 4424 17978
rect 4476 17926 4488 17978
rect 4540 17926 4552 17978
rect 4604 17926 10988 17978
rect 11040 17926 11052 17978
rect 11104 17926 11116 17978
rect 11168 17926 11180 17978
rect 11232 17926 11244 17978
rect 11296 17926 17680 17978
rect 17732 17926 17744 17978
rect 17796 17926 17808 17978
rect 17860 17926 17872 17978
rect 17924 17926 17936 17978
rect 17988 17926 24372 17978
rect 24424 17926 24436 17978
rect 24488 17926 24500 17978
rect 24552 17926 24564 17978
rect 24616 17926 24628 17978
rect 24680 17926 27876 17978
rect 1104 17904 27876 17926
rect 2958 17864 2964 17876
rect 1688 17836 2964 17864
rect 1688 17737 1716 17836
rect 2958 17824 2964 17836
rect 3016 17864 3022 17876
rect 3970 17864 3976 17876
rect 3016 17836 3976 17864
rect 3016 17824 3022 17836
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5767 17867 5825 17873
rect 5767 17864 5779 17867
rect 5592 17836 5779 17864
rect 5592 17824 5598 17836
rect 5767 17833 5779 17836
rect 5813 17833 5825 17867
rect 5767 17827 5825 17833
rect 7469 17867 7527 17873
rect 7469 17833 7481 17867
rect 7515 17864 7527 17867
rect 8294 17864 8300 17876
rect 7515 17836 8300 17864
rect 7515 17833 7527 17836
rect 7469 17827 7527 17833
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 8570 17864 8576 17876
rect 8531 17836 8576 17864
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 10689 17867 10747 17873
rect 10689 17833 10701 17867
rect 10735 17864 10747 17867
rect 11790 17864 11796 17876
rect 10735 17836 11796 17864
rect 10735 17833 10747 17836
rect 10689 17827 10747 17833
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 15378 17864 15384 17876
rect 13136 17836 15056 17864
rect 15339 17836 15384 17864
rect 13136 17824 13142 17836
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 9456 17768 12434 17796
rect 9456 17756 9462 17768
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1946 17728 1952 17740
rect 1907 17700 1952 17728
rect 1673 17691 1731 17697
rect 1946 17688 1952 17700
rect 2004 17688 2010 17740
rect 3421 17731 3479 17737
rect 3421 17697 3433 17731
rect 3467 17728 3479 17731
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 3467 17700 4353 17728
rect 3467 17697 3479 17700
rect 3421 17691 3479 17697
rect 4341 17697 4353 17700
rect 4387 17697 4399 17731
rect 9490 17728 9496 17740
rect 9451 17700 9496 17728
rect 4341 17691 4399 17697
rect 9490 17688 9496 17700
rect 9548 17728 9554 17740
rect 9548 17700 9904 17728
rect 9548 17688 9554 17700
rect 3050 17620 3056 17672
rect 3108 17620 3114 17672
rect 3970 17660 3976 17672
rect 3931 17632 3976 17660
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 6972 17632 7389 17660
rect 6972 17620 6978 17632
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 7561 17663 7619 17669
rect 7561 17660 7573 17663
rect 7524 17632 7573 17660
rect 7524 17620 7530 17632
rect 7561 17629 7573 17632
rect 7607 17629 7619 17663
rect 7561 17623 7619 17629
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 8904 17632 9229 17660
rect 8904 17620 8910 17632
rect 9217 17629 9229 17632
rect 9263 17660 9275 17663
rect 9674 17660 9680 17672
rect 9263 17632 9680 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 6365 17595 6423 17601
rect 4632 17564 4738 17592
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4632 17524 4660 17564
rect 6365 17561 6377 17595
rect 6411 17592 6423 17595
rect 9876 17592 9904 17700
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 11701 17731 11759 17737
rect 11701 17728 11713 17731
rect 10008 17700 11713 17728
rect 10008 17688 10014 17700
rect 11701 17697 11713 17700
rect 11747 17697 11759 17731
rect 11701 17691 11759 17697
rect 10502 17660 10508 17672
rect 10463 17632 10508 17660
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 11514 17660 11520 17672
rect 11475 17632 11520 17660
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 11698 17592 11704 17604
rect 6411 17564 8892 17592
rect 9876 17564 11704 17592
rect 6411 17561 6423 17564
rect 6365 17555 6423 17561
rect 8864 17536 8892 17564
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 12406 17592 12434 17768
rect 12710 17756 12716 17808
rect 12768 17796 12774 17808
rect 12768 17768 14964 17796
rect 12768 17756 12774 17768
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 13262 17728 13268 17740
rect 12943 17700 13268 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 13648 17700 14872 17728
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12710 17592 12716 17604
rect 12406 17564 12716 17592
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 13446 17592 13452 17604
rect 13407 17564 13452 17592
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 6914 17524 6920 17536
rect 4120 17496 4660 17524
rect 6875 17496 6920 17524
rect 4120 17484 4126 17496
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 8846 17484 8852 17536
rect 8904 17484 8910 17536
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 10928 17496 11161 17524
rect 10928 17484 10934 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 11609 17527 11667 17533
rect 11609 17493 11621 17527
rect 11655 17524 11667 17527
rect 12342 17524 12348 17536
rect 11655 17496 12348 17524
rect 11655 17493 11667 17496
rect 11609 17487 11667 17493
rect 12342 17484 12348 17496
rect 12400 17524 12406 17536
rect 13648 17524 13676 17700
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 14844 17669 14872 17700
rect 14461 17663 14519 17669
rect 14461 17660 14473 17663
rect 14056 17632 14473 17660
rect 14056 17620 14062 17632
rect 14461 17629 14473 17632
rect 14507 17629 14519 17663
rect 14461 17623 14519 17629
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17629 14887 17663
rect 14936 17660 14964 17768
rect 15028 17728 15056 17836
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 18785 17867 18843 17873
rect 15856 17836 17632 17864
rect 15028 17700 15516 17728
rect 15488 17669 15516 17700
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 14936 17632 15301 17660
rect 14829 17623 14887 17629
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17629 15531 17663
rect 15473 17623 15531 17629
rect 13722 17552 13728 17604
rect 13780 17592 13786 17604
rect 14553 17595 14611 17601
rect 14553 17592 14565 17595
rect 13780 17564 14565 17592
rect 13780 17552 13786 17564
rect 14553 17561 14565 17564
rect 14599 17561 14611 17595
rect 14553 17555 14611 17561
rect 14645 17595 14703 17601
rect 14645 17561 14657 17595
rect 14691 17592 14703 17595
rect 14918 17592 14924 17604
rect 14691 17564 14924 17592
rect 14691 17561 14703 17564
rect 14645 17555 14703 17561
rect 12400 17496 13676 17524
rect 12400 17484 12406 17496
rect 14090 17484 14096 17536
rect 14148 17524 14154 17536
rect 14277 17527 14335 17533
rect 14277 17524 14289 17527
rect 14148 17496 14289 17524
rect 14148 17484 14154 17496
rect 14277 17493 14289 17496
rect 14323 17493 14335 17527
rect 14568 17524 14596 17555
rect 14918 17552 14924 17564
rect 14976 17552 14982 17604
rect 15856 17524 15884 17836
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 16942 17728 16948 17740
rect 15979 17700 16948 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 17604 17728 17632 17836
rect 18785 17833 18797 17867
rect 18831 17864 18843 17867
rect 19610 17864 19616 17876
rect 18831 17836 19616 17864
rect 18831 17833 18843 17836
rect 18785 17827 18843 17833
rect 19610 17824 19616 17836
rect 19668 17864 19674 17876
rect 21818 17864 21824 17876
rect 19668 17836 21824 17864
rect 19668 17824 19674 17836
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 25593 17867 25651 17873
rect 25593 17864 25605 17867
rect 22066 17836 25605 17864
rect 17678 17756 17684 17808
rect 17736 17796 17742 17808
rect 22066 17796 22094 17836
rect 25593 17833 25605 17836
rect 25639 17833 25651 17867
rect 25593 17827 25651 17833
rect 22278 17796 22284 17808
rect 17736 17768 22094 17796
rect 22204 17768 22284 17796
rect 17736 17756 17742 17768
rect 18230 17728 18236 17740
rect 17604 17700 18236 17728
rect 18230 17688 18236 17700
rect 18288 17728 18294 17740
rect 20806 17728 20812 17740
rect 18288 17700 18920 17728
rect 18288 17688 18294 17700
rect 18892 17669 18920 17700
rect 20456 17700 20812 17728
rect 20456 17669 20484 17700
rect 20806 17688 20812 17700
rect 20864 17688 20870 17740
rect 22204 17737 22232 17768
rect 22278 17756 22284 17768
rect 22336 17756 22342 17808
rect 22189 17731 22247 17737
rect 22189 17697 22201 17731
rect 22235 17697 22247 17731
rect 22462 17728 22468 17740
rect 22423 17700 22468 17728
rect 22189 17691 22247 17697
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 20441 17663 20499 17669
rect 20441 17660 20453 17663
rect 19659 17632 20453 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 20441 17629 20453 17632
rect 20487 17629 20499 17663
rect 20622 17660 20628 17672
rect 20583 17632 20628 17660
rect 20441 17623 20499 17629
rect 16209 17595 16267 17601
rect 16209 17561 16221 17595
rect 16255 17561 16267 17595
rect 17586 17592 17592 17604
rect 17434 17564 17592 17592
rect 16209 17555 16267 17561
rect 14568 17496 15884 17524
rect 16224 17524 16252 17555
rect 17586 17552 17592 17564
rect 17644 17552 17650 17604
rect 17034 17524 17040 17536
rect 16224 17496 17040 17524
rect 14277 17487 14335 17493
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 17494 17484 17500 17536
rect 17552 17524 17558 17536
rect 17681 17527 17739 17533
rect 17681 17524 17693 17527
rect 17552 17496 17693 17524
rect 17552 17484 17558 17496
rect 17681 17493 17693 17496
rect 17727 17493 17739 17527
rect 18138 17524 18144 17536
rect 18099 17496 18144 17524
rect 17681 17487 17739 17493
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 18708 17524 18736 17623
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 21177 17663 21235 17669
rect 21177 17660 21189 17663
rect 20824 17632 21189 17660
rect 19797 17595 19855 17601
rect 19797 17561 19809 17595
rect 19843 17592 19855 17595
rect 20640 17592 20668 17620
rect 20824 17604 20852 17632
rect 21177 17629 21189 17632
rect 21223 17629 21235 17663
rect 22094 17660 22100 17672
rect 22055 17632 22100 17660
rect 21177 17623 21235 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 22278 17620 22284 17672
rect 22336 17660 22342 17672
rect 23109 17663 23167 17669
rect 23109 17660 23121 17663
rect 22336 17632 23121 17660
rect 22336 17620 22342 17632
rect 23109 17629 23121 17632
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 23566 17620 23572 17672
rect 23624 17660 23630 17672
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23624 17632 23673 17660
rect 23624 17620 23630 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23750 17620 23756 17672
rect 23808 17660 23814 17672
rect 24578 17660 24584 17672
rect 23808 17632 24584 17660
rect 23808 17620 23814 17632
rect 24578 17620 24584 17632
rect 24636 17660 24642 17672
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24636 17632 24685 17660
rect 24636 17620 24642 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 19843 17564 20668 17592
rect 19843 17561 19855 17564
rect 19797 17555 19855 17561
rect 20806 17552 20812 17604
rect 20864 17552 20870 17604
rect 19702 17524 19708 17536
rect 18708 17496 19708 17524
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19978 17524 19984 17536
rect 19939 17496 19984 17524
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20530 17524 20536 17536
rect 20491 17496 20536 17524
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 22002 17524 22008 17536
rect 21315 17496 22008 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 22922 17524 22928 17536
rect 22883 17496 22928 17524
rect 22922 17484 22928 17496
rect 22980 17484 22986 17536
rect 23845 17527 23903 17533
rect 23845 17493 23857 17527
rect 23891 17524 23903 17527
rect 23934 17524 23940 17536
rect 23891 17496 23940 17524
rect 23891 17493 23903 17496
rect 23845 17487 23903 17493
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24268 17496 24685 17524
rect 24268 17484 24274 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 25608 17524 25636 17827
rect 27062 17728 27068 17740
rect 27023 17700 27068 17728
rect 27062 17688 27068 17700
rect 27120 17688 27126 17740
rect 27338 17728 27344 17740
rect 27299 17700 27344 17728
rect 27338 17688 27344 17700
rect 27396 17688 27402 17740
rect 26510 17552 26516 17604
rect 26568 17552 26574 17604
rect 26326 17524 26332 17536
rect 25608 17496 26332 17524
rect 24673 17487 24731 17493
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 1104 17434 28032 17456
rect 1104 17382 7642 17434
rect 7694 17382 7706 17434
rect 7758 17382 7770 17434
rect 7822 17382 7834 17434
rect 7886 17382 7898 17434
rect 7950 17382 14334 17434
rect 14386 17382 14398 17434
rect 14450 17382 14462 17434
rect 14514 17382 14526 17434
rect 14578 17382 14590 17434
rect 14642 17382 21026 17434
rect 21078 17382 21090 17434
rect 21142 17382 21154 17434
rect 21206 17382 21218 17434
rect 21270 17382 21282 17434
rect 21334 17382 27718 17434
rect 27770 17382 27782 17434
rect 27834 17382 27846 17434
rect 27898 17382 27910 17434
rect 27962 17382 27974 17434
rect 28026 17382 28032 17434
rect 1104 17360 28032 17382
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2501 17323 2559 17329
rect 2501 17320 2513 17323
rect 2280 17292 2513 17320
rect 2280 17280 2286 17292
rect 2501 17289 2513 17292
rect 2547 17289 2559 17323
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 2501 17283 2559 17289
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 4062 17320 4068 17332
rect 4023 17292 4068 17320
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4614 17320 4620 17332
rect 4575 17292 4620 17320
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 6549 17323 6607 17329
rect 6549 17289 6561 17323
rect 6595 17320 6607 17323
rect 6638 17320 6644 17332
rect 6595 17292 6644 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 10042 17320 10048 17332
rect 9692 17292 10048 17320
rect 5074 17212 5080 17264
rect 5132 17252 5138 17264
rect 9692 17252 9720 17292
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 10836 17292 10977 17320
rect 10836 17280 10842 17292
rect 10965 17289 10977 17292
rect 11011 17289 11023 17323
rect 13722 17320 13728 17332
rect 10965 17283 11023 17289
rect 11808 17292 13728 17320
rect 5132 17224 9720 17252
rect 9861 17255 9919 17261
rect 5132 17212 5138 17224
rect 9861 17221 9873 17255
rect 9907 17252 9919 17255
rect 10686 17252 10692 17264
rect 9907 17224 10692 17252
rect 9907 17221 9919 17224
rect 9861 17215 9919 17221
rect 10686 17212 10692 17224
rect 10744 17252 10750 17264
rect 10873 17255 10931 17261
rect 10873 17252 10885 17255
rect 10744 17224 10885 17252
rect 10744 17212 10750 17224
rect 10873 17221 10885 17224
rect 10919 17221 10931 17255
rect 10873 17215 10931 17221
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11701 17255 11759 17261
rect 11701 17252 11713 17255
rect 11480 17224 11713 17252
rect 11480 17212 11486 17224
rect 11701 17221 11713 17224
rect 11747 17221 11759 17255
rect 11701 17215 11759 17221
rect 1578 17184 1584 17196
rect 1539 17156 1584 17184
rect 1578 17144 1584 17156
rect 1636 17144 1642 17196
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17153 3111 17187
rect 3053 17147 3111 17153
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17184 3295 17187
rect 3510 17184 3516 17196
rect 3283 17156 3516 17184
rect 3283 17153 3295 17156
rect 3237 17147 3295 17153
rect 3068 17116 3096 17147
rect 3510 17144 3516 17156
rect 3568 17184 3574 17196
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3568 17156 3893 17184
rect 3568 17144 3574 17156
rect 3881 17153 3893 17156
rect 3927 17153 3939 17187
rect 3881 17147 3939 17153
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 4080 17116 4108 17147
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4212 17156 4537 17184
rect 4212 17144 4218 17156
rect 4525 17153 4537 17156
rect 4571 17153 4583 17187
rect 4706 17184 4712 17196
rect 4667 17156 4712 17184
rect 4525 17147 4583 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 5644 17116 5672 17147
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7662 17187 7720 17193
rect 7662 17184 7674 17187
rect 6788 17156 7674 17184
rect 6788 17144 6794 17156
rect 7662 17153 7674 17156
rect 7708 17153 7720 17187
rect 7662 17147 7720 17153
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9398 17184 9404 17196
rect 8996 17156 9404 17184
rect 8996 17144 9002 17156
rect 9398 17144 9404 17156
rect 9456 17184 9462 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9456 17156 9781 17184
rect 9456 17144 9462 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10652 17156 10793 17184
rect 10652 17144 10658 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 7926 17116 7932 17128
rect 3068 17088 5672 17116
rect 7887 17088 7932 17116
rect 4172 17060 4200 17088
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 11149 17119 11207 17125
rect 10008 17088 10053 17116
rect 10008 17076 10014 17088
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 11808 17116 11836 17292
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 14277 17323 14335 17329
rect 14277 17289 14289 17323
rect 14323 17320 14335 17323
rect 15194 17320 15200 17332
rect 14323 17292 15200 17320
rect 14323 17289 14335 17292
rect 14277 17283 14335 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 18616 17292 19472 17320
rect 12894 17252 12900 17264
rect 11900 17224 12900 17252
rect 11900 17193 11928 17224
rect 12894 17212 12900 17224
rect 12952 17252 12958 17264
rect 13078 17252 13084 17264
rect 12952 17224 13084 17252
rect 12952 17212 12958 17224
rect 13078 17212 13084 17224
rect 13136 17212 13142 17264
rect 13446 17212 13452 17264
rect 13504 17212 13510 17264
rect 18138 17252 18144 17264
rect 14844 17224 18144 17252
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 11992 17116 12020 17147
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 14844 17193 14872 17224
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 14608 17156 14841 17184
rect 14608 17144 14614 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 16850 17184 16856 17196
rect 16811 17156 16856 17184
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17678 17184 17684 17196
rect 17639 17156 17684 17184
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 11195 17088 12020 17116
rect 12529 17119 12587 17125
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 12529 17085 12541 17119
rect 12575 17085 12587 17119
rect 12529 17079 12587 17085
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17116 12863 17119
rect 13814 17116 13820 17128
rect 12851 17088 13820 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 1762 17048 1768 17060
rect 1675 17020 1768 17048
rect 1762 17008 1768 17020
rect 1820 17048 1826 17060
rect 1820 17020 2774 17048
rect 1820 17008 1826 17020
rect 2746 16980 2774 17020
rect 4154 17008 4160 17060
rect 4212 17008 4218 17060
rect 4264 17020 7052 17048
rect 4264 16980 4292 17020
rect 5718 16980 5724 16992
rect 2746 16952 4292 16980
rect 5679 16952 5724 16980
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 7024 16980 7052 17020
rect 8294 17008 8300 17060
rect 8352 17048 8358 17060
rect 9401 17051 9459 17057
rect 9401 17048 9413 17051
rect 8352 17020 9413 17048
rect 8352 17008 8358 17020
rect 9401 17017 9413 17020
rect 9447 17017 9459 17051
rect 9401 17011 9459 17017
rect 10502 17008 10508 17060
rect 10560 17048 10566 17060
rect 10597 17051 10655 17057
rect 10597 17048 10609 17051
rect 10560 17020 10609 17048
rect 10560 17008 10566 17020
rect 10597 17017 10609 17020
rect 10643 17017 10655 17051
rect 12544 17048 12572 17079
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 15746 17116 15752 17128
rect 15707 17088 15752 17116
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 17310 17076 17316 17128
rect 17368 17116 17374 17128
rect 17589 17119 17647 17125
rect 17589 17116 17601 17119
rect 17368 17088 17601 17116
rect 17368 17076 17374 17088
rect 17589 17085 17601 17088
rect 17635 17085 17647 17119
rect 17589 17079 17647 17085
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18616 17116 18644 17292
rect 19334 17252 19340 17264
rect 19295 17224 19340 17252
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 19444 17184 19472 17292
rect 24578 17280 24584 17332
rect 24636 17320 24642 17332
rect 25685 17323 25743 17329
rect 25685 17320 25697 17323
rect 24636 17292 25697 17320
rect 24636 17280 24642 17292
rect 25685 17289 25697 17292
rect 25731 17289 25743 17323
rect 25685 17283 25743 17289
rect 19978 17212 19984 17264
rect 20036 17252 20042 17264
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 20036 17224 20453 17252
rect 20036 17212 20042 17224
rect 20441 17221 20453 17224
rect 20487 17221 20499 17255
rect 22186 17252 22192 17264
rect 20441 17215 20499 17221
rect 21192 17224 22192 17252
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 18782 17116 18788 17128
rect 18095 17088 18644 17116
rect 18743 17088 18788 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 19260 17116 19288 17170
rect 19444 17156 20085 17184
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20162 17144 20168 17196
rect 20220 17184 20226 17196
rect 20220 17156 20265 17184
rect 20220 17144 20226 17156
rect 20346 17144 20352 17196
rect 20404 17184 20410 17196
rect 20404 17156 20449 17184
rect 20404 17144 20410 17156
rect 20530 17144 20536 17196
rect 20588 17193 20594 17196
rect 21192 17193 21220 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 24210 17252 24216 17264
rect 24171 17224 24216 17252
rect 24210 17212 24216 17224
rect 24268 17212 24274 17264
rect 22376 17196 22428 17202
rect 20588 17184 20596 17193
rect 21177 17187 21235 17193
rect 20588 17156 20633 17184
rect 20588 17147 20596 17156
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 21284 17156 22376 17184
rect 20588 17144 20594 17147
rect 21284 17116 21312 17156
rect 23934 17184 23940 17196
rect 23895 17156 23940 17184
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 26418 17184 26424 17196
rect 25346 17156 25452 17184
rect 26379 17156 26424 17184
rect 22376 17138 22428 17144
rect 25424 17128 25452 17156
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 19208 17088 21312 17116
rect 21453 17119 21511 17125
rect 19208 17076 19214 17088
rect 21453 17085 21465 17119
rect 21499 17116 21511 17119
rect 22094 17116 22100 17128
rect 21499 17088 22100 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 22094 17076 22100 17088
rect 22152 17076 22158 17128
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17085 22523 17119
rect 23290 17116 23296 17128
rect 23251 17088 23296 17116
rect 22465 17079 22523 17085
rect 10597 17011 10655 17017
rect 11532 17020 12572 17048
rect 7190 16980 7196 16992
rect 7024 16952 7196 16980
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 8846 16980 8852 16992
rect 8807 16952 8852 16980
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 11532 16980 11560 17020
rect 13906 17008 13912 17060
rect 13964 17048 13970 17060
rect 17037 17051 17095 17057
rect 13964 17020 16988 17048
rect 13964 17008 13970 17020
rect 9548 16952 11560 16980
rect 9548 16940 9554 16952
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 14642 16980 14648 16992
rect 11756 16952 14648 16980
rect 11756 16940 11762 16952
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 16960 16980 16988 17020
rect 17037 17017 17049 17051
rect 17083 17048 17095 17051
rect 21082 17048 21088 17060
rect 17083 17020 21088 17048
rect 17083 17017 17095 17020
rect 17037 17011 17095 17017
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 21269 17051 21327 17057
rect 21269 17048 21281 17051
rect 21192 17020 21281 17048
rect 17402 16980 17408 16992
rect 16960 16952 17408 16980
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 20717 16983 20775 16989
rect 20717 16949 20729 16983
rect 20763 16980 20775 16983
rect 21192 16980 21220 17020
rect 21269 17017 21281 17020
rect 21315 17017 21327 17051
rect 21269 17011 21327 17017
rect 21910 17008 21916 17060
rect 21968 17048 21974 17060
rect 22480 17048 22508 17079
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 25406 17076 25412 17128
rect 25464 17076 25470 17128
rect 21968 17020 22508 17048
rect 21968 17008 21974 17020
rect 21358 16980 21364 16992
rect 20763 16952 21220 16980
rect 21319 16952 21364 16980
rect 20763 16949 20775 16952
rect 20717 16943 20775 16949
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 26326 16980 26332 16992
rect 26287 16952 26332 16980
rect 26326 16940 26332 16952
rect 26384 16940 26390 16992
rect 1104 16890 27876 16912
rect 1104 16838 4296 16890
rect 4348 16838 4360 16890
rect 4412 16838 4424 16890
rect 4476 16838 4488 16890
rect 4540 16838 4552 16890
rect 4604 16838 10988 16890
rect 11040 16838 11052 16890
rect 11104 16838 11116 16890
rect 11168 16838 11180 16890
rect 11232 16838 11244 16890
rect 11296 16838 17680 16890
rect 17732 16838 17744 16890
rect 17796 16838 17808 16890
rect 17860 16838 17872 16890
rect 17924 16838 17936 16890
rect 17988 16838 24372 16890
rect 24424 16838 24436 16890
rect 24488 16838 24500 16890
rect 24552 16838 24564 16890
rect 24616 16838 24628 16890
rect 24680 16838 27876 16890
rect 1104 16816 27876 16838
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 4157 16779 4215 16785
rect 4157 16776 4169 16779
rect 4120 16748 4169 16776
rect 4120 16736 4126 16748
rect 4157 16745 4169 16748
rect 4203 16776 4215 16779
rect 5994 16776 6000 16788
rect 4203 16748 6000 16776
rect 4203 16745 4215 16748
rect 4157 16739 4215 16745
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 6730 16776 6736 16788
rect 6691 16748 6736 16776
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 8754 16776 8760 16788
rect 7248 16748 8760 16776
rect 7248 16736 7254 16748
rect 8754 16736 8760 16748
rect 8812 16736 8818 16788
rect 8846 16736 8852 16788
rect 8904 16776 8910 16788
rect 10594 16776 10600 16788
rect 8904 16748 10600 16776
rect 8904 16736 8910 16748
rect 10594 16736 10600 16748
rect 10652 16776 10658 16788
rect 10689 16779 10747 16785
rect 10689 16776 10701 16779
rect 10652 16748 10701 16776
rect 10652 16736 10658 16748
rect 10689 16745 10701 16748
rect 10735 16745 10747 16779
rect 10689 16739 10747 16745
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 14550 16776 14556 16788
rect 13320 16748 14556 16776
rect 13320 16736 13326 16748
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 14700 16748 18460 16776
rect 14700 16736 14706 16748
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 14826 16708 14832 16720
rect 7984 16680 14832 16708
rect 7984 16668 7990 16680
rect 14826 16668 14832 16680
rect 14884 16668 14890 16720
rect 18432 16708 18460 16748
rect 18782 16736 18788 16788
rect 18840 16776 18846 16788
rect 19610 16776 19616 16788
rect 18840 16748 19616 16776
rect 18840 16736 18846 16748
rect 19610 16736 19616 16748
rect 19668 16776 19674 16788
rect 21910 16776 21916 16788
rect 19668 16748 21916 16776
rect 19668 16736 19674 16748
rect 21910 16736 21916 16748
rect 21968 16776 21974 16788
rect 21968 16748 22094 16776
rect 21968 16736 21974 16748
rect 20898 16708 20904 16720
rect 18432 16680 20904 16708
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16640 5043 16643
rect 5074 16640 5080 16652
rect 5031 16612 5080 16640
rect 5031 16609 5043 16612
rect 4985 16603 5043 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 8021 16643 8079 16649
rect 8021 16640 8033 16643
rect 6972 16612 8033 16640
rect 6972 16600 6978 16612
rect 8021 16609 8033 16612
rect 8067 16640 8079 16643
rect 8938 16640 8944 16652
rect 8067 16612 8944 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 8938 16600 8944 16612
rect 8996 16600 9002 16652
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 9950 16640 9956 16652
rect 9732 16612 9956 16640
rect 9732 16600 9738 16612
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 14277 16643 14335 16649
rect 14277 16640 14289 16643
rect 10744 16612 14289 16640
rect 10744 16600 10750 16612
rect 14277 16609 14289 16612
rect 14323 16609 14335 16643
rect 17586 16640 17592 16652
rect 17547 16612 17592 16640
rect 14277 16603 14335 16609
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 18432 16649 18460 16680
rect 20898 16668 20904 16680
rect 20956 16668 20962 16720
rect 22066 16708 22094 16748
rect 22462 16736 22468 16788
rect 22520 16776 22526 16788
rect 23385 16779 23443 16785
rect 23385 16776 23397 16779
rect 22520 16748 23397 16776
rect 22520 16736 22526 16748
rect 23385 16745 23397 16748
rect 23431 16745 23443 16779
rect 23385 16739 23443 16745
rect 22066 16680 23612 16708
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16609 18475 16643
rect 23474 16640 23480 16652
rect 23435 16612 23480 16640
rect 18417 16603 18475 16609
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 23584 16640 23612 16680
rect 24670 16640 24676 16652
rect 23584 16612 24676 16640
rect 24670 16600 24676 16612
rect 24728 16640 24734 16652
rect 24857 16643 24915 16649
rect 24857 16640 24869 16643
rect 24728 16612 24869 16640
rect 24728 16600 24734 16612
rect 24857 16609 24869 16612
rect 24903 16609 24915 16643
rect 24857 16603 24915 16609
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 26421 16643 26479 16649
rect 26421 16640 26433 16643
rect 26292 16612 26433 16640
rect 26292 16600 26298 16612
rect 26421 16609 26433 16612
rect 26467 16640 26479 16643
rect 27154 16640 27160 16652
rect 26467 16612 27160 16640
rect 26467 16609 26479 16612
rect 26421 16603 26479 16609
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 25320 16584 25372 16590
rect 2222 16572 2228 16584
rect 2183 16544 2228 16572
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3786 16572 3792 16584
rect 3007 16544 3792 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 3878 16532 3884 16584
rect 3936 16572 3942 16584
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3936 16544 3985 16572
rect 3936 16532 3942 16544
rect 3973 16541 3985 16544
rect 4019 16572 4031 16575
rect 4798 16572 4804 16584
rect 4019 16544 4804 16572
rect 4019 16541 4031 16544
rect 3973 16535 4031 16541
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 5721 16575 5779 16581
rect 5721 16541 5733 16575
rect 5767 16541 5779 16575
rect 6638 16572 6644 16584
rect 6599 16544 6644 16572
rect 5721 16535 5779 16541
rect 5736 16504 5764 16535
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 9490 16572 9496 16584
rect 6748 16544 9496 16572
rect 6748 16504 6776 16544
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 9769 16575 9827 16581
rect 9769 16541 9781 16575
rect 9815 16572 9827 16575
rect 10042 16572 10048 16584
rect 9815 16544 10048 16572
rect 9815 16541 9827 16544
rect 9769 16535 9827 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 13722 16572 13728 16584
rect 13683 16544 13728 16572
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 15010 16572 15016 16584
rect 14691 16544 15016 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 18690 16572 18696 16584
rect 18538 16544 18696 16572
rect 18690 16532 18696 16544
rect 18748 16572 18754 16584
rect 19150 16572 19156 16584
rect 18748 16544 19156 16572
rect 18748 16532 18754 16544
rect 19150 16532 19156 16544
rect 19208 16532 19214 16584
rect 19610 16572 19616 16584
rect 19571 16544 19616 16572
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16572 20499 16575
rect 20530 16572 20536 16584
rect 20487 16544 20536 16572
rect 20487 16541 20499 16544
rect 20441 16535 20499 16541
rect 20530 16532 20536 16544
rect 20588 16572 20594 16584
rect 20714 16572 20720 16584
rect 20588 16544 20720 16572
rect 20588 16532 20594 16544
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 21082 16532 21088 16584
rect 21140 16572 21146 16584
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 21140 16544 21189 16572
rect 21140 16532 21146 16544
rect 21177 16541 21189 16544
rect 21223 16541 21235 16575
rect 23661 16575 23719 16581
rect 23661 16572 23673 16575
rect 21177 16535 21235 16541
rect 22066 16544 23673 16572
rect 5736 16476 6776 16504
rect 7745 16507 7803 16513
rect 7745 16473 7757 16507
rect 7791 16504 7803 16507
rect 8110 16504 8116 16516
rect 7791 16476 8116 16504
rect 7791 16473 7803 16476
rect 7745 16467 7803 16473
rect 8110 16464 8116 16476
rect 8168 16464 8174 16516
rect 9861 16507 9919 16513
rect 9861 16473 9873 16507
rect 9907 16504 9919 16507
rect 11241 16507 11299 16513
rect 9907 16476 10824 16504
rect 9907 16473 9919 16476
rect 9861 16467 9919 16473
rect 10796 16448 10824 16476
rect 11241 16473 11253 16507
rect 11287 16504 11299 16507
rect 11330 16504 11336 16516
rect 11287 16476 11336 16504
rect 11287 16473 11299 16476
rect 11241 16467 11299 16473
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 11440 16476 14565 16504
rect 2038 16436 2044 16448
rect 1999 16408 2044 16436
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 5537 16439 5595 16445
rect 2832 16408 2877 16436
rect 2832 16396 2838 16408
rect 5537 16405 5549 16439
rect 5583 16436 5595 16439
rect 5994 16436 6000 16448
rect 5583 16408 6000 16436
rect 5583 16405 5595 16408
rect 5537 16399 5595 16405
rect 5994 16396 6000 16408
rect 6052 16396 6058 16448
rect 8018 16396 8024 16448
rect 8076 16436 8082 16448
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 8076 16408 9413 16436
rect 8076 16396 8082 16408
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 9401 16399 9459 16405
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 10962 16436 10968 16448
rect 10836 16408 10968 16436
rect 10836 16396 10842 16408
rect 10962 16396 10968 16408
rect 11020 16436 11026 16448
rect 11440 16436 11468 16476
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 14762 16507 14820 16513
rect 14762 16473 14774 16507
rect 14808 16473 14820 16507
rect 15378 16504 15384 16516
rect 15339 16476 15384 16504
rect 14762 16467 14820 16473
rect 11020 16408 11468 16436
rect 11020 16396 11026 16408
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 12529 16439 12587 16445
rect 12529 16436 12541 16439
rect 11848 16408 12541 16436
rect 11848 16396 11854 16408
rect 12529 16405 12541 16408
rect 12575 16405 12587 16439
rect 12529 16399 12587 16405
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 13504 16408 13553 16436
rect 13504 16396 13510 16408
rect 13541 16405 13553 16408
rect 13587 16405 13599 16439
rect 13541 16399 13599 16405
rect 13630 16396 13636 16448
rect 13688 16436 13694 16448
rect 14777 16436 14805 16467
rect 15378 16464 15384 16476
rect 15436 16464 15442 16516
rect 19702 16464 19708 16516
rect 19760 16504 19766 16516
rect 22066 16504 22094 16544
rect 23661 16541 23673 16544
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 25590 16572 25596 16584
rect 25372 16544 25596 16572
rect 25590 16532 25596 16544
rect 25648 16572 25654 16584
rect 25648 16544 26358 16572
rect 25648 16532 25654 16544
rect 25320 16526 25372 16532
rect 19760 16476 22094 16504
rect 19760 16464 19766 16476
rect 22186 16464 22192 16516
rect 22244 16504 22250 16516
rect 23382 16504 23388 16516
rect 22244 16476 23060 16504
rect 23343 16476 23388 16504
rect 22244 16464 22250 16476
rect 14918 16436 14924 16448
rect 13688 16408 14805 16436
rect 14879 16408 14924 16436
rect 13688 16396 13694 16408
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 15712 16408 16681 16436
rect 15712 16396 15718 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 16669 16399 16727 16405
rect 22370 16396 22376 16448
rect 22428 16436 22434 16448
rect 22465 16439 22523 16445
rect 22465 16436 22477 16439
rect 22428 16408 22477 16436
rect 22428 16396 22434 16408
rect 22465 16405 22477 16408
rect 22511 16405 22523 16439
rect 23032 16436 23060 16476
rect 23382 16464 23388 16476
rect 23440 16464 23446 16516
rect 23566 16464 23572 16516
rect 23624 16504 23630 16516
rect 23934 16504 23940 16516
rect 23624 16476 23940 16504
rect 23624 16464 23630 16476
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 25498 16464 25504 16516
rect 25556 16504 25562 16516
rect 25685 16507 25743 16513
rect 25685 16504 25697 16507
rect 25556 16476 25697 16504
rect 25556 16464 25562 16476
rect 25685 16473 25697 16476
rect 25731 16473 25743 16507
rect 26970 16504 26976 16516
rect 26931 16476 26976 16504
rect 25685 16467 25743 16473
rect 26970 16464 26976 16476
rect 27028 16464 27034 16516
rect 23845 16439 23903 16445
rect 23845 16436 23857 16439
rect 23032 16408 23857 16436
rect 22465 16399 22523 16405
rect 23845 16405 23857 16408
rect 23891 16405 23903 16439
rect 23845 16399 23903 16405
rect 1104 16346 28032 16368
rect 1104 16294 7642 16346
rect 7694 16294 7706 16346
rect 7758 16294 7770 16346
rect 7822 16294 7834 16346
rect 7886 16294 7898 16346
rect 7950 16294 14334 16346
rect 14386 16294 14398 16346
rect 14450 16294 14462 16346
rect 14514 16294 14526 16346
rect 14578 16294 14590 16346
rect 14642 16294 21026 16346
rect 21078 16294 21090 16346
rect 21142 16294 21154 16346
rect 21206 16294 21218 16346
rect 21270 16294 21282 16346
rect 21334 16294 27718 16346
rect 27770 16294 27782 16346
rect 27834 16294 27846 16346
rect 27898 16294 27910 16346
rect 27962 16294 27974 16346
rect 28026 16294 28032 16346
rect 1104 16272 28032 16294
rect 2222 16192 2228 16244
rect 2280 16232 2286 16244
rect 3605 16235 3663 16241
rect 3605 16232 3617 16235
rect 2280 16204 3617 16232
rect 2280 16192 2286 16204
rect 3605 16201 3617 16204
rect 3651 16201 3663 16235
rect 3605 16195 3663 16201
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 4249 16235 4307 16241
rect 4249 16232 4261 16235
rect 3844 16204 4261 16232
rect 3844 16192 3850 16204
rect 4249 16201 4261 16204
rect 4295 16232 4307 16235
rect 8205 16235 8263 16241
rect 4295 16204 6592 16232
rect 4295 16201 4307 16204
rect 4249 16195 4307 16201
rect 2038 16124 2044 16176
rect 2096 16164 2102 16176
rect 2133 16167 2191 16173
rect 2133 16164 2145 16167
rect 2096 16136 2145 16164
rect 2096 16124 2102 16136
rect 2133 16133 2145 16136
rect 2179 16133 2191 16167
rect 3694 16164 3700 16176
rect 3358 16136 3700 16164
rect 2133 16127 2191 16133
rect 3694 16124 3700 16136
rect 3752 16124 3758 16176
rect 5718 16164 5724 16176
rect 5290 16136 5724 16164
rect 5718 16124 5724 16136
rect 5776 16124 5782 16176
rect 5994 16056 6000 16108
rect 6052 16096 6058 16108
rect 6564 16105 6592 16204
rect 8205 16201 8217 16235
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 10594 16232 10600 16244
rect 10091 16204 10600 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 8220 16164 8248 16195
rect 10594 16192 10600 16204
rect 10652 16232 10658 16244
rect 10962 16232 10968 16244
rect 10652 16204 10968 16232
rect 10652 16192 10658 16204
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12802 16232 12808 16244
rect 12483 16204 12808 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 15930 16232 15936 16244
rect 15891 16204 15936 16232
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17310 16232 17316 16244
rect 17271 16204 17316 16232
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17402 16192 17408 16244
rect 17460 16232 17466 16244
rect 18690 16232 18696 16244
rect 17460 16204 17505 16232
rect 18651 16204 18696 16232
rect 17460 16192 17466 16204
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 20806 16232 20812 16244
rect 19536 16204 20812 16232
rect 8910 16167 8968 16173
rect 8910 16164 8922 16167
rect 8220 16136 8922 16164
rect 8910 16133 8922 16136
rect 8956 16133 8968 16167
rect 8910 16127 8968 16133
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 10873 16167 10931 16173
rect 10873 16164 10885 16167
rect 10744 16136 10885 16164
rect 10744 16124 10750 16136
rect 10873 16133 10885 16136
rect 10919 16133 10931 16167
rect 10873 16127 10931 16133
rect 13725 16167 13783 16173
rect 13725 16133 13737 16167
rect 13771 16164 13783 16167
rect 14182 16164 14188 16176
rect 13771 16136 14188 16164
rect 13771 16133 13783 16136
rect 13725 16127 13783 16133
rect 14182 16124 14188 16136
rect 14240 16124 14246 16176
rect 14461 16167 14519 16173
rect 14461 16133 14473 16167
rect 14507 16164 14519 16167
rect 14734 16164 14740 16176
rect 14507 16136 14740 16164
rect 14507 16133 14519 16136
rect 14461 16127 14519 16133
rect 14734 16124 14740 16136
rect 14792 16124 14798 16176
rect 15746 16164 15752 16176
rect 15686 16136 15752 16164
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 15948 16164 15976 16192
rect 19536 16176 19564 16204
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 21269 16235 21327 16241
rect 21269 16201 21281 16235
rect 21315 16232 21327 16235
rect 22278 16232 22284 16244
rect 21315 16204 22284 16232
rect 21315 16201 21327 16204
rect 21269 16195 21327 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 27154 16232 27160 16244
rect 22388 16204 24256 16232
rect 27115 16204 27160 16232
rect 22388 16176 22416 16204
rect 19518 16164 19524 16176
rect 15948 16136 19524 16164
rect 19518 16124 19524 16136
rect 19576 16124 19582 16176
rect 19981 16167 20039 16173
rect 19981 16133 19993 16167
rect 20027 16164 20039 16167
rect 22370 16164 22376 16176
rect 20027 16136 22376 16164
rect 20027 16133 20039 16136
rect 19981 16127 20039 16133
rect 22370 16124 22376 16136
rect 22428 16124 22434 16176
rect 23290 16124 23296 16176
rect 23348 16124 23354 16176
rect 24228 16173 24256 16204
rect 27154 16192 27160 16204
rect 27212 16192 27218 16244
rect 24213 16167 24271 16173
rect 24213 16133 24225 16167
rect 24259 16133 24271 16167
rect 26513 16167 26571 16173
rect 26513 16164 26525 16167
rect 24213 16127 24271 16133
rect 26206 16136 26525 16164
rect 6549 16099 6607 16105
rect 6052 16068 6097 16096
rect 6052 16056 6058 16068
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16065 7435 16099
rect 8018 16096 8024 16108
rect 7979 16068 8024 16096
rect 7377 16059 7435 16065
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 2774 16028 2780 16040
rect 1903 16000 2780 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 7392 16028 7420 16059
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 8812 16068 10793 16096
rect 8812 16056 8818 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 11020 16068 11161 16096
rect 11020 16056 11026 16068
rect 11149 16065 11161 16068
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 21634 16096 21640 16108
rect 20947 16068 21640 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 8294 16028 8300 16040
rect 5767 16000 5948 16028
rect 7392 16000 8300 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 5920 15960 5948 16000
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8662 16028 8668 16040
rect 8623 16000 8668 16028
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 10664 16031 10722 16037
rect 10664 16028 10676 16031
rect 10560 16000 10676 16028
rect 10560 15988 10566 16000
rect 10664 15997 10676 16000
rect 10710 16028 10722 16031
rect 14182 16028 14188 16040
rect 10710 16000 10824 16028
rect 14143 16000 14188 16028
rect 10710 15997 10722 16000
rect 10664 15991 10722 15997
rect 10796 15972 10824 16000
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 17218 16028 17224 16040
rect 17179 16000 17224 16028
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 15997 20683 16031
rect 20806 16028 20812 16040
rect 20767 16000 20812 16028
rect 20625 15991 20683 15997
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 5920 15932 6561 15960
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 6549 15923 6607 15929
rect 10042 15920 10048 15972
rect 10100 15960 10106 15972
rect 10100 15932 10640 15960
rect 10100 15920 10106 15932
rect 7561 15895 7619 15901
rect 7561 15861 7573 15895
rect 7607 15892 7619 15895
rect 9030 15892 9036 15904
rect 7607 15864 9036 15892
rect 7607 15861 7619 15864
rect 7561 15855 7619 15861
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 10502 15892 10508 15904
rect 10463 15864 10508 15892
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 10612 15892 10640 15932
rect 10778 15920 10784 15972
rect 10836 15920 10842 15972
rect 13538 15960 13544 15972
rect 12406 15932 13544 15960
rect 12406 15892 12434 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 17402 15920 17408 15972
rect 17460 15960 17466 15972
rect 20640 15960 20668 15991
rect 20806 15988 20812 16000
rect 20864 15988 20870 16040
rect 20898 15960 20904 15972
rect 17460 15932 19748 15960
rect 20640 15932 20904 15960
rect 17460 15920 17466 15932
rect 10612 15864 12434 15892
rect 17773 15895 17831 15901
rect 17773 15861 17785 15895
rect 17819 15892 17831 15895
rect 19610 15892 19616 15904
rect 17819 15864 19616 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 19720 15892 19748 15932
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 21652 15960 21680 16056
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 26206 16028 26234 16136
rect 26513 16133 26525 16136
rect 26559 16133 26571 16167
rect 26513 16127 26571 16133
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 22327 16000 26234 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 22002 15960 22008 15972
rect 21652 15932 22008 15960
rect 22002 15920 22008 15932
rect 22060 15920 22066 15972
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 23753 15963 23811 15969
rect 23753 15960 23765 15963
rect 23532 15932 23765 15960
rect 23532 15920 23538 15932
rect 23753 15929 23765 15932
rect 23799 15960 23811 15963
rect 23934 15960 23940 15972
rect 23799 15932 23940 15960
rect 23799 15929 23811 15932
rect 23753 15923 23811 15929
rect 23934 15920 23940 15932
rect 23992 15960 23998 15972
rect 26436 15960 26464 16059
rect 23992 15932 26464 15960
rect 23992 15920 23998 15932
rect 23290 15892 23296 15904
rect 19720 15864 23296 15892
rect 23290 15852 23296 15864
rect 23348 15852 23354 15904
rect 25501 15895 25559 15901
rect 25501 15861 25513 15895
rect 25547 15892 25559 15895
rect 25590 15892 25596 15904
rect 25547 15864 25596 15892
rect 25547 15861 25559 15864
rect 25501 15855 25559 15861
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 1104 15802 27876 15824
rect 1104 15750 4296 15802
rect 4348 15750 4360 15802
rect 4412 15750 4424 15802
rect 4476 15750 4488 15802
rect 4540 15750 4552 15802
rect 4604 15750 10988 15802
rect 11040 15750 11052 15802
rect 11104 15750 11116 15802
rect 11168 15750 11180 15802
rect 11232 15750 11244 15802
rect 11296 15750 17680 15802
rect 17732 15750 17744 15802
rect 17796 15750 17808 15802
rect 17860 15750 17872 15802
rect 17924 15750 17936 15802
rect 17988 15750 24372 15802
rect 24424 15750 24436 15802
rect 24488 15750 24500 15802
rect 24552 15750 24564 15802
rect 24616 15750 24628 15802
rect 24680 15750 27876 15802
rect 1104 15728 27876 15750
rect 4154 15688 4160 15700
rect 4115 15660 4160 15688
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 8846 15688 8852 15700
rect 8352 15660 8852 15688
rect 8352 15648 8358 15660
rect 8846 15648 8852 15660
rect 8904 15688 8910 15700
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 8904 15660 9229 15688
rect 8904 15648 8910 15660
rect 9217 15657 9229 15660
rect 9263 15657 9275 15691
rect 9217 15651 9275 15657
rect 6822 15580 6828 15632
rect 6880 15620 6886 15632
rect 7745 15623 7803 15629
rect 7745 15620 7757 15623
rect 6880 15592 7757 15620
rect 6880 15580 6886 15592
rect 7745 15589 7757 15592
rect 7791 15589 7803 15623
rect 9232 15620 9260 15651
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 12584 15660 13277 15688
rect 12584 15648 12590 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 14829 15691 14887 15697
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 15378 15688 15384 15700
rect 14875 15660 15384 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 11517 15623 11575 15629
rect 9232 15592 11284 15620
rect 7745 15583 7803 15589
rect 10686 15552 10692 15564
rect 10647 15524 10692 15552
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4890 15484 4896 15496
rect 4212 15456 4896 15484
rect 4212 15444 4218 15456
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 5534 15484 5540 15496
rect 5495 15456 5540 15484
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7156 15456 7757 15484
rect 7156 15444 7162 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9214 15484 9220 15496
rect 9171 15456 9220 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 10778 15444 10784 15496
rect 10836 15484 10842 15496
rect 11256 15493 11284 15592
rect 11517 15589 11529 15623
rect 11563 15620 11575 15623
rect 12618 15620 12624 15632
rect 11563 15592 12624 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 13280 15552 13308 15651
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 16850 15648 16856 15700
rect 16908 15688 16914 15700
rect 16945 15691 17003 15697
rect 16945 15688 16957 15691
rect 16908 15660 16957 15688
rect 16908 15648 16914 15660
rect 16945 15657 16957 15660
rect 16991 15657 17003 15691
rect 16945 15651 17003 15657
rect 18877 15691 18935 15697
rect 18877 15657 18889 15691
rect 18923 15688 18935 15691
rect 19702 15688 19708 15700
rect 18923 15660 19708 15688
rect 18923 15657 18935 15660
rect 18877 15651 18935 15657
rect 19702 15648 19708 15660
rect 19760 15648 19766 15700
rect 20073 15691 20131 15697
rect 20073 15657 20085 15691
rect 20119 15688 20131 15691
rect 20806 15688 20812 15700
rect 20119 15660 20812 15688
rect 20119 15657 20131 15660
rect 20073 15651 20131 15657
rect 20806 15648 20812 15660
rect 20864 15688 20870 15700
rect 22465 15691 22523 15697
rect 20864 15660 21496 15688
rect 20864 15648 20870 15660
rect 13280 15524 14596 15552
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10836 15456 10977 15484
rect 10836 15444 10842 15456
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11882 15484 11888 15496
rect 11287 15456 11888 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 1949 15419 2007 15425
rect 1949 15385 1961 15419
rect 1995 15385 2007 15419
rect 3326 15416 3332 15428
rect 3174 15388 3332 15416
rect 1949 15379 2007 15385
rect 1964 15348 1992 15379
rect 3326 15376 3332 15388
rect 3384 15376 3390 15428
rect 4062 15416 4068 15428
rect 4023 15388 4068 15416
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 5810 15416 5816 15428
rect 5771 15388 5816 15416
rect 5810 15376 5816 15388
rect 5868 15376 5874 15428
rect 9232 15416 9260 15444
rect 10980 15416 11008 15447
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 14568 15493 14596 15524
rect 17586 15512 17592 15564
rect 17644 15552 17650 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 17644 15524 18429 15552
rect 17644 15512 17650 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 21468 15552 21496 15660
rect 22465 15657 22477 15691
rect 22511 15688 22523 15691
rect 23382 15688 23388 15700
rect 22511 15660 23388 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 23382 15648 23388 15660
rect 23440 15648 23446 15700
rect 24854 15688 24860 15700
rect 24815 15660 24860 15688
rect 24854 15648 24860 15660
rect 24912 15648 24918 15700
rect 26326 15688 26332 15700
rect 25516 15660 26332 15688
rect 22094 15580 22100 15632
rect 22152 15620 22158 15632
rect 24581 15623 24639 15629
rect 24581 15620 24593 15623
rect 22152 15592 24593 15620
rect 22152 15580 22158 15592
rect 24581 15589 24593 15592
rect 24627 15589 24639 15623
rect 24581 15583 24639 15589
rect 22005 15555 22063 15561
rect 22005 15552 22017 15555
rect 21468 15524 22017 15552
rect 18417 15515 18475 15521
rect 22005 15521 22017 15524
rect 22051 15521 22063 15555
rect 23382 15552 23388 15564
rect 23343 15524 23388 15552
rect 22005 15515 22063 15521
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 25516 15561 25544 15660
rect 26326 15648 26332 15660
rect 26384 15648 26390 15700
rect 23661 15555 23719 15561
rect 23661 15521 23673 15555
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 25501 15555 25559 15561
rect 25501 15521 25513 15555
rect 25547 15521 25559 15555
rect 25774 15552 25780 15564
rect 25735 15524 25780 15552
rect 25501 15515 25559 15521
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 14016 15456 14289 15484
rect 11422 15416 11428 15428
rect 5920 15388 6302 15416
rect 9232 15388 11428 15416
rect 2866 15348 2872 15360
rect 1964 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3418 15348 3424 15360
rect 3379 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 4985 15351 5043 15357
rect 4985 15317 4997 15351
rect 5031 15348 5043 15351
rect 5920 15348 5948 15388
rect 11422 15376 11428 15388
rect 11480 15376 11486 15428
rect 11790 15376 11796 15428
rect 11848 15416 11854 15428
rect 11977 15419 12035 15425
rect 11977 15416 11989 15419
rect 11848 15388 11989 15416
rect 11848 15376 11854 15388
rect 11977 15385 11989 15388
rect 12023 15385 12035 15419
rect 11977 15379 12035 15385
rect 13446 15376 13452 15428
rect 13504 15416 13510 15428
rect 14016 15416 14044 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 14697 15487 14755 15493
rect 14697 15453 14709 15487
rect 14743 15484 14755 15487
rect 14826 15484 14832 15496
rect 14743 15456 14832 15484
rect 14743 15453 14755 15456
rect 14697 15447 14755 15453
rect 14826 15444 14832 15456
rect 14884 15484 14890 15496
rect 15654 15484 15660 15496
rect 14884 15456 15516 15484
rect 15615 15456 15660 15484
rect 14884 15444 14890 15456
rect 13504 15388 14044 15416
rect 13504 15376 13510 15388
rect 7282 15348 7288 15360
rect 5031 15320 5948 15348
rect 7243 15320 7288 15348
rect 5031 15317 5043 15320
rect 4985 15311 5043 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 8352 15320 8493 15348
rect 8352 15308 8358 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 8481 15311 8539 15317
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15348 9643 15351
rect 9674 15348 9680 15360
rect 9631 15320 9680 15348
rect 9631 15317 9643 15320
rect 9585 15311 9643 15317
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 14016 15348 14044 15388
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 14461 15419 14519 15425
rect 14461 15416 14473 15419
rect 14148 15388 14473 15416
rect 14148 15376 14154 15388
rect 14461 15385 14473 15388
rect 14507 15385 14519 15419
rect 15488 15416 15516 15456
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 17494 15444 17500 15496
rect 17552 15484 17558 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 17552 15456 18521 15484
rect 17552 15444 17558 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 18509 15447 18567 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 21358 15484 21364 15496
rect 19720 15456 21364 15484
rect 19720 15416 19748 15456
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 22097 15487 22155 15493
rect 21508 15456 21553 15484
rect 21508 15444 21514 15456
rect 22097 15453 22109 15487
rect 22143 15453 22155 15487
rect 22097 15447 22155 15453
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15484 23351 15487
rect 23474 15484 23480 15496
rect 23339 15456 23480 15484
rect 23339 15453 23351 15456
rect 23293 15447 23351 15453
rect 15488 15388 19748 15416
rect 21208 15419 21266 15425
rect 14461 15379 14519 15385
rect 21208 15385 21220 15419
rect 21254 15416 21266 15419
rect 22112 15416 22140 15447
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 23676 15484 23704 15515
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 26970 15512 26976 15564
rect 27028 15512 27034 15564
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 23676 15456 24777 15484
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 26988 15484 27016 15512
rect 24912 15456 24957 15484
rect 26910 15456 27016 15484
rect 24912 15444 24918 15456
rect 25038 15416 25044 15428
rect 21254 15388 21680 15416
rect 22112 15388 24716 15416
rect 24999 15388 25044 15416
rect 21254 15385 21266 15388
rect 21208 15379 21266 15385
rect 16390 15348 16396 15360
rect 14016 15320 16396 15348
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 19426 15348 19432 15360
rect 19387 15320 19432 15348
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 21652 15348 21680 15388
rect 22922 15348 22928 15360
rect 21652 15320 22928 15348
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 24688 15348 24716 15388
rect 25038 15376 25044 15388
rect 25096 15376 25102 15428
rect 26602 15348 26608 15360
rect 24688 15320 26608 15348
rect 26602 15308 26608 15320
rect 26660 15348 26666 15360
rect 27249 15351 27307 15357
rect 27249 15348 27261 15351
rect 26660 15320 27261 15348
rect 26660 15308 26666 15320
rect 27249 15317 27261 15320
rect 27295 15317 27307 15351
rect 27249 15311 27307 15317
rect 1104 15258 28032 15280
rect 1104 15206 7642 15258
rect 7694 15206 7706 15258
rect 7758 15206 7770 15258
rect 7822 15206 7834 15258
rect 7886 15206 7898 15258
rect 7950 15206 14334 15258
rect 14386 15206 14398 15258
rect 14450 15206 14462 15258
rect 14514 15206 14526 15258
rect 14578 15206 14590 15258
rect 14642 15206 21026 15258
rect 21078 15206 21090 15258
rect 21142 15206 21154 15258
rect 21206 15206 21218 15258
rect 21270 15206 21282 15258
rect 21334 15206 27718 15258
rect 27770 15206 27782 15258
rect 27834 15206 27846 15258
rect 27898 15206 27910 15258
rect 27962 15206 27974 15258
rect 28026 15206 28032 15258
rect 1104 15184 28032 15206
rect 3694 15144 3700 15156
rect 3655 15116 3700 15144
rect 3694 15104 3700 15116
rect 3752 15104 3758 15156
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 5868 15116 6653 15144
rect 5868 15104 5874 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 8021 15147 8079 15153
rect 8021 15113 8033 15147
rect 8067 15144 8079 15147
rect 8202 15144 8208 15156
rect 8067 15116 8208 15144
rect 8067 15113 8079 15116
rect 8021 15107 8079 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 10505 15147 10563 15153
rect 10505 15113 10517 15147
rect 10551 15144 10563 15147
rect 10686 15144 10692 15156
rect 10551 15116 10692 15144
rect 10551 15113 10563 15116
rect 10505 15107 10563 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 10836 15116 12081 15144
rect 10836 15104 10842 15116
rect 12069 15113 12081 15116
rect 12115 15144 12127 15147
rect 13449 15147 13507 15153
rect 12115 15116 12388 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 1670 15036 1676 15088
rect 1728 15076 1734 15088
rect 2133 15079 2191 15085
rect 2133 15076 2145 15079
rect 1728 15048 2145 15076
rect 1728 15036 1734 15048
rect 2133 15045 2145 15048
rect 2179 15045 2191 15079
rect 2866 15076 2872 15088
rect 2827 15048 2872 15076
rect 2133 15039 2191 15045
rect 2866 15036 2872 15048
rect 2924 15036 2930 15088
rect 4154 15036 4160 15088
rect 4212 15036 4218 15088
rect 4982 15036 4988 15088
rect 5040 15036 5046 15088
rect 8220 15076 8248 15104
rect 8220 15048 9536 15076
rect 2222 15008 2228 15020
rect 2183 14980 2228 15008
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 3145 15011 3203 15017
rect 3145 15008 3157 15011
rect 2832 14980 3157 15008
rect 2832 14968 2838 14980
rect 3145 14977 3157 14980
rect 3191 15008 3203 15011
rect 3418 15008 3424 15020
rect 3191 14980 3424 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 4172 15008 4200 15036
rect 3835 14980 4200 15008
rect 6733 15011 6791 15017
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 7282 15008 7288 15020
rect 6779 14980 7288 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 8478 15008 8484 15020
rect 8439 14980 8484 15008
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9381 15011 9439 15017
rect 9381 15008 9393 15011
rect 9088 14980 9393 15008
rect 9088 14968 9094 14980
rect 9381 14977 9393 14980
rect 9427 14977 9439 15011
rect 9508 15008 9536 15048
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 9732 15048 12296 15076
rect 9732 15036 9738 15048
rect 10778 15008 10784 15020
rect 9508 14980 10784 15008
rect 9381 14971 9439 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10928 14980 10977 15008
rect 10928 14968 10934 14980
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 4212 14912 4261 14940
rect 4212 14900 4218 14912
rect 4249 14909 4261 14912
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 6822 14940 6828 14952
rect 4571 14912 6828 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8720 14912 9137 14940
rect 8720 14900 8726 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 12158 14940 12164 14952
rect 12119 14912 12164 14940
rect 9125 14903 9183 14909
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 5997 14875 6055 14881
rect 5997 14872 6009 14875
rect 5868 14844 6009 14872
rect 5868 14832 5874 14844
rect 5997 14841 6009 14844
rect 6043 14872 6055 14875
rect 7098 14872 7104 14884
rect 6043 14844 7104 14872
rect 6043 14841 6055 14844
rect 5997 14835 6055 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 7377 14807 7435 14813
rect 7377 14773 7389 14807
rect 7423 14804 7435 14807
rect 7466 14804 7472 14816
rect 7423 14776 7472 14804
rect 7423 14773 7435 14776
rect 7377 14767 7435 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 9030 14804 9036 14816
rect 8619 14776 9036 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 9140 14804 9168 14903
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12268 14949 12296 15048
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14909 12311 14943
rect 12360 14940 12388 15116
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 15194 15144 15200 15156
rect 13495 15116 15200 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 17126 15144 17132 15156
rect 15764 15116 17132 15144
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15654 15076 15660 15088
rect 14783 15048 15660 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 15654 15036 15660 15048
rect 15712 15036 15718 15088
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 15764 15008 15792 15116
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 17310 15104 17316 15156
rect 17368 15144 17374 15156
rect 17497 15147 17555 15153
rect 17497 15144 17509 15147
rect 17368 15116 17509 15144
rect 17368 15104 17374 15116
rect 17497 15113 17509 15116
rect 17543 15113 17555 15147
rect 17497 15107 17555 15113
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20162 15144 20168 15156
rect 19751 15116 20168 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 26418 15144 26424 15156
rect 24412 15116 26424 15144
rect 15841 15079 15899 15085
rect 15841 15045 15853 15079
rect 15887 15076 15899 15079
rect 17586 15076 17592 15088
rect 15887 15048 17592 15076
rect 15887 15045 15899 15048
rect 15841 15039 15899 15045
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 18632 15079 18690 15085
rect 18632 15045 18644 15079
rect 18678 15076 18690 15079
rect 19426 15076 19432 15088
rect 18678 15048 19432 15076
rect 18678 15045 18690 15048
rect 18632 15039 18690 15045
rect 19426 15036 19432 15048
rect 19484 15036 19490 15088
rect 19518 15036 19524 15088
rect 19576 15076 19582 15088
rect 22462 15076 22468 15088
rect 19576 15048 19621 15076
rect 22375 15048 22468 15076
rect 19576 15036 19582 15048
rect 22462 15036 22468 15048
rect 22520 15076 22526 15088
rect 22520 15048 24348 15076
rect 22520 15036 22526 15048
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 13596 14980 15945 15008
rect 13596 14968 13602 14980
rect 15933 14977 15945 14980
rect 15979 14977 15991 15011
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 15933 14971 15991 14977
rect 16316 14980 17049 15008
rect 15654 14940 15660 14952
rect 12360 14912 15660 14940
rect 12253 14903 12311 14909
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14940 15807 14943
rect 15795 14912 16252 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 10410 14804 10416 14816
rect 9140 14776 10416 14804
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 11149 14807 11207 14813
rect 11149 14773 11161 14807
rect 11195 14804 11207 14807
rect 11606 14804 11612 14816
rect 11195 14776 11612 14804
rect 11195 14773 11207 14776
rect 11149 14767 11207 14773
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 16224 14804 16252 14912
rect 16316 14881 16344 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 17037 14971 17095 14977
rect 17144 14980 18889 15008
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 17144 14940 17172 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 19334 15008 19340 15020
rect 19295 14980 19340 15008
rect 18877 14971 18935 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 15008 20499 15011
rect 21450 15008 21456 15020
rect 20487 14980 21456 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 22373 15011 22431 15017
rect 22373 14977 22385 15011
rect 22419 15008 22431 15011
rect 22646 15008 22652 15020
rect 22419 14980 22652 15008
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 15008 23443 15011
rect 23474 15008 23480 15020
rect 23431 14980 23480 15008
rect 23431 14977 23443 14980
rect 23385 14971 23443 14977
rect 23474 14968 23480 14980
rect 23532 15008 23538 15020
rect 23750 15008 23756 15020
rect 23532 14980 23756 15008
rect 23532 14968 23538 14980
rect 23750 14968 23756 14980
rect 23808 14968 23814 15020
rect 20162 14940 20168 14952
rect 16448 14912 17172 14940
rect 20123 14912 20168 14940
rect 16448 14900 16454 14912
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20898 14900 20904 14952
rect 20956 14940 20962 14952
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 20956 14912 22569 14940
rect 20956 14900 20962 14912
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 23198 14900 23204 14952
rect 23256 14940 23262 14952
rect 24320 14949 24348 15048
rect 24412 15017 24440 15116
rect 26418 15104 26424 15116
rect 26476 15104 26482 15156
rect 27154 15144 27160 15156
rect 27115 15116 27160 15144
rect 27154 15104 27160 15116
rect 27212 15104 27218 15156
rect 25596 15020 25648 15026
rect 24397 15011 24455 15017
rect 24397 14977 24409 15011
rect 24443 14977 24455 15011
rect 24397 14971 24455 14977
rect 25314 14968 25320 15020
rect 25372 15008 25378 15020
rect 25501 15011 25559 15017
rect 25501 15008 25513 15011
rect 25372 14980 25513 15008
rect 25372 14968 25378 14980
rect 25501 14977 25513 14980
rect 25547 14977 25559 15011
rect 25501 14971 25559 14977
rect 25596 14962 25648 14968
rect 23293 14943 23351 14949
rect 23293 14940 23305 14943
rect 23256 14912 23305 14940
rect 23256 14900 23262 14912
rect 23293 14909 23305 14912
rect 23339 14909 23351 14943
rect 23293 14903 23351 14909
rect 24305 14943 24363 14949
rect 24305 14909 24317 14943
rect 24351 14909 24363 14943
rect 24305 14903 24363 14909
rect 24765 14943 24823 14949
rect 24765 14909 24777 14943
rect 24811 14940 24823 14943
rect 24854 14940 24860 14952
rect 24811 14912 24860 14940
rect 24811 14909 24823 14912
rect 24765 14903 24823 14909
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 26513 14943 26571 14949
rect 26513 14909 26525 14943
rect 26559 14940 26571 14943
rect 26602 14940 26608 14952
rect 26559 14912 26608 14940
rect 26559 14909 26571 14912
rect 26513 14903 26571 14909
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 16301 14875 16359 14881
rect 16301 14841 16313 14875
rect 16347 14841 16359 14875
rect 16301 14835 16359 14841
rect 16500 14844 17264 14872
rect 16500 14804 16528 14844
rect 17236 14816 17264 14844
rect 16850 14804 16856 14816
rect 11756 14776 11801 14804
rect 16224 14776 16528 14804
rect 16811 14776 16856 14804
rect 11756 14764 11762 14776
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17218 14764 17224 14816
rect 17276 14804 17282 14816
rect 20916 14804 20944 14900
rect 23753 14875 23811 14881
rect 23753 14841 23765 14875
rect 23799 14872 23811 14875
rect 25038 14872 25044 14884
rect 23799 14844 25044 14872
rect 23799 14841 23811 14844
rect 23753 14835 23811 14841
rect 25038 14832 25044 14844
rect 25096 14832 25102 14884
rect 17276 14776 20944 14804
rect 17276 14764 17282 14776
rect 21450 14764 21456 14816
rect 21508 14804 21514 14816
rect 22005 14807 22063 14813
rect 22005 14804 22017 14807
rect 21508 14776 22017 14804
rect 21508 14764 21514 14776
rect 22005 14773 22017 14776
rect 22051 14773 22063 14807
rect 22005 14767 22063 14773
rect 1104 14714 27876 14736
rect 1104 14662 4296 14714
rect 4348 14662 4360 14714
rect 4412 14662 4424 14714
rect 4476 14662 4488 14714
rect 4540 14662 4552 14714
rect 4604 14662 10988 14714
rect 11040 14662 11052 14714
rect 11104 14662 11116 14714
rect 11168 14662 11180 14714
rect 11232 14662 11244 14714
rect 11296 14662 17680 14714
rect 17732 14662 17744 14714
rect 17796 14662 17808 14714
rect 17860 14662 17872 14714
rect 17924 14662 17936 14714
rect 17988 14662 24372 14714
rect 24424 14662 24436 14714
rect 24488 14662 24500 14714
rect 24552 14662 24564 14714
rect 24616 14662 24628 14714
rect 24680 14662 27876 14714
rect 1104 14640 27876 14662
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4212 14572 4261 14600
rect 4212 14560 4218 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4982 14600 4988 14612
rect 4943 14572 4988 14600
rect 4249 14563 4307 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5592 14572 5641 14600
rect 5592 14560 5598 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 11698 14600 11704 14612
rect 5629 14563 5687 14569
rect 8496 14572 11704 14600
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 1728 14436 7021 14464
rect 1728 14424 1734 14436
rect 7009 14433 7021 14436
rect 7055 14464 7067 14467
rect 8294 14464 8300 14476
rect 7055 14436 8300 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 1854 14288 1860 14340
rect 1912 14328 1918 14340
rect 1912 14300 1978 14328
rect 1912 14288 1918 14300
rect 3050 14288 3056 14340
rect 3108 14328 3114 14340
rect 3145 14331 3203 14337
rect 3145 14328 3157 14331
rect 3108 14300 3157 14328
rect 3108 14288 3114 14300
rect 3145 14297 3157 14300
rect 3191 14297 3203 14331
rect 3145 14291 3203 14297
rect 1673 14263 1731 14269
rect 1673 14229 1685 14263
rect 1719 14260 1731 14263
rect 2130 14260 2136 14272
rect 1719 14232 2136 14260
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 3436 14260 3464 14359
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 4028 14368 4445 14396
rect 4028 14356 4034 14368
rect 4433 14365 4445 14368
rect 4479 14365 4491 14399
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 4433 14359 4491 14365
rect 4448 14328 4476 14359
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5810 14396 5816 14408
rect 5771 14368 5816 14396
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 6549 14399 6607 14405
rect 6549 14365 6561 14399
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 8389 14399 8447 14405
rect 7791 14368 8340 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 6564 14328 6592 14359
rect 8018 14328 8024 14340
rect 4448 14300 6408 14328
rect 6564 14300 8024 14328
rect 6380 14272 6408 14300
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 8312 14328 8340 14368
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 8496 14396 8524 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12400 14572 13124 14600
rect 12400 14560 12406 14572
rect 8573 14535 8631 14541
rect 8573 14501 8585 14535
rect 8619 14501 8631 14535
rect 8573 14495 8631 14501
rect 8588 14464 8616 14495
rect 8588 14436 9996 14464
rect 9490 14396 9496 14408
rect 8435 14368 8524 14396
rect 8588 14368 9496 14396
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 8588 14328 8616 14368
rect 9490 14356 9496 14368
rect 9548 14356 9554 14408
rect 9858 14396 9864 14408
rect 9819 14368 9864 14396
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 9968 14396 9996 14436
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 11664 14436 11836 14464
rect 11664 14424 11670 14436
rect 10117 14399 10175 14405
rect 10117 14396 10129 14399
rect 9968 14368 10129 14396
rect 10117 14365 10129 14368
rect 10163 14365 10175 14399
rect 10117 14359 10175 14365
rect 10410 14356 10416 14408
rect 10468 14396 10474 14408
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 10468 14368 11713 14396
rect 10468 14356 10474 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11808 14396 11836 14436
rect 11957 14399 12015 14405
rect 11957 14396 11969 14399
rect 11808 14368 11969 14396
rect 11701 14359 11759 14365
rect 11957 14365 11969 14368
rect 12003 14365 12015 14399
rect 11957 14359 12015 14365
rect 8312 14300 8616 14328
rect 9217 14331 9275 14337
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 10502 14328 10508 14340
rect 9263 14300 10508 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 10594 14288 10600 14340
rect 10652 14328 10658 14340
rect 12066 14328 12072 14340
rect 10652 14300 12072 14328
rect 10652 14288 10658 14300
rect 12066 14288 12072 14300
rect 12124 14328 12130 14340
rect 12986 14328 12992 14340
rect 12124 14300 12992 14328
rect 12124 14288 12130 14300
rect 12986 14288 12992 14300
rect 13044 14288 13050 14340
rect 13096 14328 13124 14572
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13725 14603 13783 14609
rect 13725 14600 13737 14603
rect 13596 14572 13737 14600
rect 13596 14560 13602 14572
rect 13725 14569 13737 14572
rect 13771 14569 13783 14603
rect 13725 14563 13783 14569
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 17586 14600 17592 14612
rect 14056 14572 15056 14600
rect 17547 14572 17592 14600
rect 14056 14560 14062 14572
rect 15028 14541 15056 14572
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 19521 14603 19579 14609
rect 19521 14569 19533 14603
rect 19567 14600 19579 14603
rect 20346 14600 20352 14612
rect 19567 14572 20352 14600
rect 19567 14569 19579 14572
rect 19521 14563 19579 14569
rect 20346 14560 20352 14572
rect 20404 14560 20410 14612
rect 22462 14600 22468 14612
rect 21100 14572 22094 14600
rect 22423 14572 22468 14600
rect 15013 14535 15071 14541
rect 15013 14501 15025 14535
rect 15059 14532 15071 14535
rect 18877 14535 18935 14541
rect 15059 14504 15884 14532
rect 15059 14501 15071 14504
rect 15013 14495 15071 14501
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 13504 14436 15117 14464
rect 13504 14424 13510 14436
rect 15105 14433 15117 14436
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 14553 14399 14611 14405
rect 14553 14396 14565 14399
rect 13688 14368 14565 14396
rect 13688 14356 13694 14368
rect 14553 14365 14565 14368
rect 14599 14365 14611 14399
rect 15010 14396 15016 14408
rect 14971 14368 15016 14396
rect 14553 14359 14611 14365
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 15396 14328 15424 14359
rect 15746 14328 15752 14340
rect 13096 14300 15752 14328
rect 13096 14272 13124 14300
rect 15746 14288 15752 14300
rect 15804 14288 15810 14340
rect 15856 14328 15884 14504
rect 18877 14501 18889 14535
rect 18923 14501 18935 14535
rect 18877 14495 18935 14501
rect 18322 14464 18328 14476
rect 18283 14436 18328 14464
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 18892 14464 18920 14495
rect 18966 14492 18972 14544
rect 19024 14532 19030 14544
rect 20073 14535 20131 14541
rect 20073 14532 20085 14535
rect 19024 14504 20085 14532
rect 19024 14492 19030 14504
rect 20073 14501 20085 14504
rect 20119 14501 20131 14535
rect 21100 14532 21128 14572
rect 20073 14495 20131 14501
rect 20364 14504 21128 14532
rect 22066 14532 22094 14572
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 22646 14560 22652 14612
rect 22704 14600 22710 14612
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 22704 14572 24593 14600
rect 22704 14560 22710 14572
rect 24581 14569 24593 14572
rect 24627 14569 24639 14603
rect 24581 14563 24639 14569
rect 22664 14532 22692 14560
rect 22066 14504 22692 14532
rect 18892 14436 20300 14464
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16298 14396 16304 14408
rect 16255 14368 16304 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16476 14399 16534 14405
rect 16476 14365 16488 14399
rect 16522 14396 16534 14399
rect 16850 14396 16856 14408
rect 16522 14368 16856 14396
rect 16522 14365 16534 14368
rect 16476 14359 16534 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14396 18475 14399
rect 19334 14396 19340 14408
rect 18463 14368 19340 14396
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 19334 14356 19340 14368
rect 19392 14396 19398 14408
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19392 14368 19441 14396
rect 19392 14356 19398 14368
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 20272 14405 20300 14436
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19576 14368 19625 14396
rect 19576 14356 19582 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 20257 14399 20315 14405
rect 20257 14365 20269 14399
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 19794 14328 19800 14340
rect 15856 14300 19800 14328
rect 19794 14288 19800 14300
rect 19852 14288 19858 14340
rect 20364 14328 20392 14504
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 23017 14467 23075 14473
rect 23017 14464 23029 14467
rect 22704 14436 23029 14464
rect 22704 14424 22710 14436
rect 23017 14433 23029 14436
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20956 14368 21097 14396
rect 20956 14356 20962 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 23290 14396 23296 14408
rect 23251 14368 23296 14396
rect 21085 14359 21143 14365
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 25038 14356 25044 14408
rect 25096 14396 25102 14408
rect 25314 14396 25320 14408
rect 25096 14368 25320 14396
rect 25096 14356 25102 14368
rect 25314 14356 25320 14368
rect 25372 14356 25378 14408
rect 25590 14356 25596 14408
rect 25648 14356 25654 14408
rect 26418 14356 26424 14408
rect 26476 14396 26482 14408
rect 26881 14399 26939 14405
rect 26881 14396 26893 14399
rect 26476 14368 26893 14396
rect 26476 14356 26482 14368
rect 26881 14365 26893 14368
rect 26927 14396 26939 14399
rect 27062 14396 27068 14408
rect 26927 14368 27068 14396
rect 26927 14365 26939 14368
rect 26881 14359 26939 14365
rect 27062 14356 27068 14368
rect 27120 14356 27126 14408
rect 21358 14337 21364 14340
rect 19904 14300 20392 14328
rect 6362 14260 6368 14272
rect 2280 14232 3464 14260
rect 6323 14232 6368 14260
rect 2280 14220 2286 14232
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 7558 14220 7564 14272
rect 7616 14260 7622 14272
rect 7745 14263 7803 14269
rect 7745 14260 7757 14263
rect 7616 14232 7757 14260
rect 7616 14220 7622 14232
rect 7745 14229 7757 14232
rect 7791 14229 7803 14263
rect 7745 14223 7803 14229
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 10042 14260 10048 14272
rect 9355 14232 10048 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 11241 14263 11299 14269
rect 11241 14229 11253 14263
rect 11287 14260 11299 14263
rect 12158 14260 12164 14272
rect 11287 14232 12164 14260
rect 11287 14229 11299 14232
rect 11241 14223 11299 14229
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 13078 14260 13084 14272
rect 12991 14232 13084 14260
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 15712 14232 18521 14260
rect 15712 14220 15718 14232
rect 18509 14229 18521 14232
rect 18555 14260 18567 14263
rect 19058 14260 19064 14272
rect 18555 14232 19064 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 19058 14220 19064 14232
rect 19116 14260 19122 14272
rect 19904 14260 19932 14300
rect 21352 14291 21364 14337
rect 21416 14328 21422 14340
rect 26326 14328 26332 14340
rect 21416 14300 21452 14328
rect 26287 14300 26332 14328
rect 21358 14288 21364 14291
rect 21416 14288 21422 14300
rect 26326 14288 26332 14300
rect 26384 14288 26390 14340
rect 26786 14328 26792 14340
rect 26747 14300 26792 14328
rect 26786 14288 26792 14300
rect 26844 14288 26850 14340
rect 23198 14260 23204 14272
rect 19116 14232 19932 14260
rect 23159 14232 23204 14260
rect 19116 14220 19122 14232
rect 23198 14220 23204 14232
rect 23256 14220 23262 14272
rect 23661 14263 23719 14269
rect 23661 14229 23673 14263
rect 23707 14260 23719 14263
rect 24026 14260 24032 14272
rect 23707 14232 24032 14260
rect 23707 14229 23719 14232
rect 23661 14223 23719 14229
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 1104 14170 28032 14192
rect 1104 14118 7642 14170
rect 7694 14118 7706 14170
rect 7758 14118 7770 14170
rect 7822 14118 7834 14170
rect 7886 14118 7898 14170
rect 7950 14118 14334 14170
rect 14386 14118 14398 14170
rect 14450 14118 14462 14170
rect 14514 14118 14526 14170
rect 14578 14118 14590 14170
rect 14642 14118 21026 14170
rect 21078 14118 21090 14170
rect 21142 14118 21154 14170
rect 21206 14118 21218 14170
rect 21270 14118 21282 14170
rect 21334 14118 27718 14170
rect 27770 14118 27782 14170
rect 27834 14118 27846 14170
rect 27898 14118 27910 14170
rect 27962 14118 27974 14170
rect 28026 14118 28032 14170
rect 1104 14096 28032 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 1762 14056 1768 14068
rect 1719 14028 1768 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 2222 14056 2228 14068
rect 2183 14028 2228 14056
rect 2222 14016 2228 14028
rect 2280 14016 2286 14068
rect 3050 14056 3056 14068
rect 3011 14028 3056 14056
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3326 14016 3332 14068
rect 3384 14056 3390 14068
rect 3697 14059 3755 14065
rect 3697 14056 3709 14059
rect 3384 14028 3709 14056
rect 3384 14016 3390 14028
rect 3697 14025 3709 14028
rect 3743 14025 3755 14059
rect 3697 14019 3755 14025
rect 5997 14059 6055 14065
rect 5997 14025 6009 14059
rect 6043 14056 6055 14059
rect 7282 14056 7288 14068
rect 6043 14028 7288 14056
rect 6043 14025 6055 14028
rect 5997 14019 6055 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7558 14016 7564 14068
rect 7616 14016 7622 14068
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 9180 14028 9229 14056
rect 9180 14016 9186 14028
rect 9217 14025 9229 14028
rect 9263 14056 9275 14059
rect 9490 14056 9496 14068
rect 9263 14028 9496 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 12158 14056 12164 14068
rect 12071 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14056 12222 14068
rect 13446 14056 13452 14068
rect 12216 14028 13452 14056
rect 12216 14016 12222 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 18877 14059 18935 14065
rect 14332 14028 15700 14056
rect 14332 14016 14338 14028
rect 2130 13948 2136 14000
rect 2188 13988 2194 14000
rect 2498 13988 2504 14000
rect 2188 13960 2504 13988
rect 2188 13948 2194 13960
rect 2498 13948 2504 13960
rect 2556 13988 2562 14000
rect 7374 13988 7380 14000
rect 2556 13960 2912 13988
rect 2556 13948 2562 13960
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 2774 13920 2780 13932
rect 2455 13892 2780 13920
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 2884 13929 2912 13960
rect 5828 13960 7380 13988
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 3835 13892 4445 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4433 13889 4445 13892
rect 4479 13920 4491 13923
rect 4890 13920 4896 13932
rect 4479 13892 4896 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 1762 13744 1768 13796
rect 1820 13784 1826 13796
rect 3804 13784 3832 13883
rect 4890 13880 4896 13892
rect 4948 13920 4954 13932
rect 5828 13929 5856 13960
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 7576 13988 7604 14016
rect 7745 13991 7803 13997
rect 7745 13988 7757 13991
rect 7576 13960 7757 13988
rect 7745 13957 7757 13960
rect 7791 13957 7803 13991
rect 9030 13988 9036 14000
rect 8943 13960 9036 13988
rect 7745 13951 7803 13957
rect 9030 13948 9036 13960
rect 9088 13988 9094 14000
rect 9088 13960 15424 13988
rect 9088 13948 9094 13960
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 4948 13892 5181 13920
rect 4948 13880 4954 13892
rect 5169 13889 5181 13892
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6420 13892 6561 13920
rect 6420 13880 6426 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 7466 13920 7472 13932
rect 7427 13892 7472 13920
rect 6549 13883 6607 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 10042 13920 10048 13932
rect 10003 13892 10048 13920
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 10594 13920 10600 13932
rect 10367 13892 10600 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10594 13880 10600 13892
rect 10652 13880 10658 13932
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13920 11207 13923
rect 11422 13920 11428 13932
rect 11195 13892 11428 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4341 13855 4399 13861
rect 4341 13852 4353 13855
rect 4212 13824 4353 13852
rect 4212 13812 4218 13824
rect 4341 13821 4353 13824
rect 4387 13821 4399 13855
rect 4341 13815 4399 13821
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 6730 13852 6736 13864
rect 5307 13824 6736 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 9950 13852 9956 13864
rect 9911 13824 9956 13852
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10060 13852 10088 13880
rect 10796 13852 10824 13883
rect 10870 13852 10876 13864
rect 10060 13824 10876 13852
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11072 13852 11100 13883
rect 11422 13880 11428 13892
rect 11480 13880 11486 13932
rect 12066 13920 12072 13932
rect 12027 13892 12072 13920
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12342 13920 12348 13932
rect 12299 13892 12348 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12802 13920 12808 13932
rect 12483 13892 12808 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12952 13892 13001 13920
rect 12952 13880 12958 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 15194 13920 15200 13932
rect 15155 13892 15200 13920
rect 12989 13883 13047 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 12820 13852 12848 13880
rect 13814 13852 13820 13864
rect 11072 13824 12756 13852
rect 12820 13824 13820 13852
rect 1820 13756 3832 13784
rect 1820 13744 1826 13756
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 5408 13756 7604 13784
rect 5408 13744 5414 13756
rect 6270 13676 6276 13728
rect 6328 13716 6334 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6328 13688 6561 13716
rect 6328 13676 6334 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 7576 13716 7604 13756
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 11885 13787 11943 13793
rect 11885 13784 11897 13787
rect 11572 13756 11897 13784
rect 11572 13744 11578 13756
rect 11885 13753 11897 13756
rect 11931 13784 11943 13787
rect 11974 13784 11980 13796
rect 11931 13756 11980 13784
rect 11931 13753 11943 13756
rect 11885 13747 11943 13753
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 12728 13784 12756 13824
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13998 13852 14004 13864
rect 13924 13824 14004 13852
rect 13924 13784 13952 13824
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14734 13852 14740 13864
rect 14695 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15396 13861 15424 13960
rect 15672 13929 15700 14028
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 19334 14056 19340 14068
rect 18923 14028 19340 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 20898 14056 20904 14068
rect 19536 14028 20904 14056
rect 17764 13991 17822 13997
rect 17764 13957 17776 13991
rect 17810 13988 17822 13991
rect 18966 13988 18972 14000
rect 17810 13960 18972 13988
rect 17810 13957 17822 13960
rect 17764 13951 17822 13957
rect 18966 13948 18972 13960
rect 19024 13948 19030 14000
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 15804 13892 16865 13920
rect 15804 13880 15810 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 17497 13923 17555 13929
rect 17497 13889 17509 13923
rect 17543 13920 17555 13923
rect 17586 13920 17592 13932
rect 17543 13892 17592 13920
rect 17543 13889 17555 13892
rect 17497 13883 17555 13889
rect 17586 13880 17592 13892
rect 17644 13880 17650 13932
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13920 19395 13923
rect 19536 13920 19564 14028
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 21499 14028 22094 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 22066 13988 22094 14028
rect 25038 14016 25044 14068
rect 25096 14056 25102 14068
rect 27154 14056 27160 14068
rect 25096 14028 27160 14056
rect 25096 14016 25102 14028
rect 27154 14016 27160 14028
rect 27212 14016 27218 14068
rect 22250 13991 22308 13997
rect 22250 13988 22262 13991
rect 22066 13960 22262 13988
rect 22250 13957 22262 13960
rect 22296 13957 22308 13991
rect 26326 13988 26332 14000
rect 26266 13960 26332 13988
rect 22250 13951 22308 13957
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 19610 13929 19616 13932
rect 19383 13892 19564 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 19604 13883 19616 13929
rect 19668 13920 19674 13932
rect 21269 13923 21327 13929
rect 19668 13892 19704 13920
rect 19610 13880 19616 13883
rect 19668 13880 19674 13892
rect 21269 13889 21281 13923
rect 21315 13920 21327 13923
rect 21910 13920 21916 13932
rect 21315 13892 21916 13920
rect 21315 13889 21327 13892
rect 21269 13883 21327 13889
rect 21910 13880 21916 13892
rect 21968 13880 21974 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 23532 13892 24041 13920
rect 23532 13880 23538 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 15381 13855 15439 13861
rect 15381 13821 15393 13855
rect 15427 13821 15439 13855
rect 15381 13815 15439 13821
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 17310 13852 17316 13864
rect 15611 13824 17316 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 12728 13756 13952 13784
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 14642 13784 14648 13796
rect 14148 13756 14648 13784
rect 14148 13744 14154 13756
rect 14642 13744 14648 13756
rect 14700 13784 14706 13796
rect 15102 13784 15108 13796
rect 14700 13756 15108 13784
rect 14700 13744 14706 13756
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 15488 13784 15516 13815
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 20898 13812 20904 13864
rect 20956 13852 20962 13864
rect 22002 13852 22008 13864
rect 20956 13824 22008 13852
rect 20956 13812 20962 13824
rect 22002 13812 22008 13824
rect 22060 13812 22066 13864
rect 24305 13855 24363 13861
rect 24305 13821 24317 13855
rect 24351 13852 24363 13855
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 24351 13824 24777 13852
rect 24351 13821 24363 13824
rect 24305 13815 24363 13821
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 24765 13815 24823 13821
rect 25130 13812 25136 13864
rect 25188 13852 25194 13864
rect 26513 13855 26571 13861
rect 26513 13852 26525 13855
rect 25188 13824 26525 13852
rect 25188 13812 25194 13824
rect 26513 13821 26525 13824
rect 26559 13821 26571 13855
rect 26513 13815 26571 13821
rect 17402 13784 17408 13796
rect 15488 13756 17408 13784
rect 17402 13744 17408 13756
rect 17460 13744 17466 13796
rect 9122 13716 9128 13728
rect 7576 13688 9128 13716
rect 6549 13679 6607 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 12434 13716 12440 13728
rect 12216 13688 12440 13716
rect 12216 13676 12222 13688
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 12986 13716 12992 13728
rect 12676 13688 12992 13716
rect 12676 13676 12682 13688
rect 12986 13676 12992 13688
rect 13044 13716 13050 13728
rect 15286 13716 15292 13728
rect 13044 13688 15292 13716
rect 13044 13676 13050 13688
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 15838 13716 15844 13728
rect 15799 13688 15844 13716
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 16942 13716 16948 13728
rect 16903 13688 16948 13716
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 20714 13716 20720 13728
rect 20675 13688 20720 13716
rect 20714 13676 20720 13688
rect 20772 13676 20778 13728
rect 23382 13716 23388 13728
rect 23343 13688 23388 13716
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 24762 13676 24768 13728
rect 24820 13716 24826 13728
rect 25022 13719 25080 13725
rect 25022 13716 25034 13719
rect 24820 13688 25034 13716
rect 24820 13676 24826 13688
rect 25022 13685 25034 13688
rect 25068 13685 25080 13719
rect 25022 13679 25080 13685
rect 1104 13626 27876 13648
rect 1104 13574 4296 13626
rect 4348 13574 4360 13626
rect 4412 13574 4424 13626
rect 4476 13574 4488 13626
rect 4540 13574 4552 13626
rect 4604 13574 10988 13626
rect 11040 13574 11052 13626
rect 11104 13574 11116 13626
rect 11168 13574 11180 13626
rect 11232 13574 11244 13626
rect 11296 13574 17680 13626
rect 17732 13574 17744 13626
rect 17796 13574 17808 13626
rect 17860 13574 17872 13626
rect 17924 13574 17936 13626
rect 17988 13574 24372 13626
rect 24424 13574 24436 13626
rect 24488 13574 24500 13626
rect 24552 13574 24564 13626
rect 24616 13574 24628 13626
rect 24680 13574 27876 13626
rect 1104 13552 27876 13574
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 8294 13512 8300 13524
rect 5592 13484 8300 13512
rect 5592 13472 5598 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 9122 13512 9128 13524
rect 8628 13484 9128 13512
rect 8628 13472 8634 13484
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 11701 13515 11759 13521
rect 9916 13484 10548 13512
rect 9916 13472 9922 13484
rect 4816 13416 6040 13444
rect 4816 13385 4844 13416
rect 6012 13385 6040 13416
rect 10520 13388 10548 13484
rect 11701 13481 11713 13515
rect 11747 13512 11759 13515
rect 12434 13512 12440 13524
rect 11747 13484 12440 13512
rect 11747 13481 11759 13484
rect 11701 13475 11759 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 12618 13512 12624 13524
rect 12575 13484 12624 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 15194 13512 15200 13524
rect 12768 13484 15200 13512
rect 12768 13472 12774 13484
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 16853 13515 16911 13521
rect 15344 13484 16804 13512
rect 15344 13472 15350 13484
rect 13722 13444 13728 13456
rect 11532 13416 13216 13444
rect 13683 13416 13728 13444
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13345 6055 13379
rect 6270 13376 6276 13388
rect 6231 13348 6276 13376
rect 5997 13339 6055 13345
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 7340 13348 8432 13376
rect 7340 13336 7346 13348
rect 1946 13308 1952 13320
rect 1907 13280 1952 13308
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4706 13308 4712 13320
rect 4111 13280 4712 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 1857 13243 1915 13249
rect 1857 13209 1869 13243
rect 1903 13240 1915 13243
rect 2774 13240 2780 13252
rect 1903 13212 2780 13240
rect 1903 13209 1915 13212
rect 1857 13203 1915 13209
rect 2774 13200 2780 13212
rect 2832 13200 2838 13252
rect 3252 13240 3280 13271
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5258 13308 5264 13320
rect 4939 13280 5264 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 5408 13280 5453 13308
rect 5408 13268 5414 13280
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 8294 13308 8300 13320
rect 5592 13280 5637 13308
rect 8255 13280 8300 13308
rect 5592 13268 5598 13280
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 8404 13308 8432 13348
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 11532 13385 11560 13416
rect 11517 13379 11575 13385
rect 10560 13348 10653 13376
rect 10560 13336 10566 13348
rect 11517 13345 11529 13379
rect 11563 13345 11575 13379
rect 12066 13376 12072 13388
rect 11517 13339 11575 13345
rect 11624 13348 12072 13376
rect 10238 13311 10296 13317
rect 10238 13308 10250 13311
rect 8404 13280 10250 13308
rect 10238 13277 10250 13280
rect 10284 13277 10296 13311
rect 10238 13271 10296 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13308 11115 13311
rect 11624 13308 11652 13348
rect 12066 13336 12072 13348
rect 12124 13376 12130 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12124 13348 12725 13376
rect 12124 13336 12130 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 13188 13376 13216 13416
rect 13722 13404 13728 13416
rect 13780 13444 13786 13456
rect 14090 13444 14096 13456
rect 13780 13416 14096 13444
rect 13780 13404 13786 13416
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 16776 13444 16804 13484
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 17218 13512 17224 13524
rect 16899 13484 17224 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 18322 13512 18328 13524
rect 18187 13484 18328 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18322 13472 18328 13484
rect 18380 13512 18386 13524
rect 21177 13515 21235 13521
rect 18380 13484 20116 13512
rect 18380 13472 18386 13484
rect 16776 13416 18092 13444
rect 13906 13376 13912 13388
rect 13188 13348 13912 13376
rect 12713 13339 12771 13345
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14277 13379 14335 13385
rect 14277 13345 14289 13379
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15194 13376 15200 13388
rect 14599 13348 15200 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 11103 13280 11652 13308
rect 11977 13311 12035 13317
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 12158 13308 12164 13320
rect 12023 13280 12164 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 14182 13308 14188 13320
rect 12820 13280 14188 13308
rect 6546 13240 6552 13252
rect 3252 13212 6552 13240
rect 6546 13200 6552 13212
rect 6604 13200 6610 13252
rect 6730 13200 6736 13252
rect 6788 13200 6794 13252
rect 8573 13243 8631 13249
rect 8573 13209 8585 13243
rect 8619 13240 8631 13243
rect 9398 13240 9404 13252
rect 8619 13212 9404 13240
rect 8619 13209 8631 13212
rect 8573 13203 8631 13209
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 12820 13240 12848 13280
rect 14182 13268 14188 13280
rect 14240 13308 14246 13320
rect 14292 13308 14320 13339
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 17310 13336 17316 13388
rect 17368 13376 17374 13388
rect 17368 13348 17632 13376
rect 17368 13336 17374 13348
rect 16758 13308 16764 13320
rect 14240 13280 14320 13308
rect 16719 13280 16764 13308
rect 14240 13268 14246 13280
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 17402 13308 17408 13320
rect 17363 13280 17408 13308
rect 16853 13271 16911 13277
rect 9508 13212 12848 13240
rect 12897 13243 12955 13249
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 2501 13175 2559 13181
rect 2501 13172 2513 13175
rect 2280 13144 2513 13172
rect 2280 13132 2286 13144
rect 2501 13141 2513 13144
rect 2547 13141 2559 13175
rect 2501 13135 2559 13141
rect 3421 13175 3479 13181
rect 3421 13141 3433 13175
rect 3467 13172 3479 13175
rect 4154 13172 4160 13184
rect 3467 13144 4160 13172
rect 3467 13141 3479 13144
rect 3421 13135 3479 13141
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 5350 13172 5356 13184
rect 4295 13144 5356 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 7558 13172 7564 13184
rect 5583 13144 7564 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 7745 13175 7803 13181
rect 7745 13141 7757 13175
rect 7791 13172 7803 13175
rect 8018 13172 8024 13184
rect 7791 13144 8024 13172
rect 7791 13141 7803 13144
rect 7745 13135 7803 13141
rect 8018 13132 8024 13144
rect 8076 13172 8082 13184
rect 9508 13172 9536 13212
rect 12897 13209 12909 13243
rect 12943 13240 12955 13243
rect 13078 13240 13084 13252
rect 12943 13212 13084 13240
rect 12943 13209 12955 13212
rect 12897 13203 12955 13209
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13173 13243 13231 13249
rect 13173 13209 13185 13243
rect 13219 13240 13231 13243
rect 13446 13240 13452 13252
rect 13219 13212 13452 13240
rect 13219 13209 13231 13212
rect 13173 13203 13231 13209
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 14274 13240 14280 13252
rect 13596 13212 14280 13240
rect 13596 13200 13602 13212
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 15286 13200 15292 13252
rect 15344 13200 15350 13252
rect 16868 13240 16896 13271
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 17604 13317 17632 13348
rect 18064 13317 18092 13416
rect 20088 13388 20116 13484
rect 21177 13481 21189 13515
rect 21223 13512 21235 13515
rect 21223 13484 22968 13512
rect 21223 13481 21235 13484
rect 21177 13475 21235 13481
rect 22940 13444 22968 13484
rect 23198 13472 23204 13524
rect 23256 13512 23262 13524
rect 23385 13515 23443 13521
rect 23385 13512 23397 13515
rect 23256 13484 23397 13512
rect 23256 13472 23262 13484
rect 23385 13481 23397 13484
rect 23431 13481 23443 13515
rect 24762 13512 24768 13524
rect 24723 13484 24768 13512
rect 23385 13475 23443 13481
rect 24762 13472 24768 13484
rect 24820 13472 24826 13524
rect 27062 13512 27068 13524
rect 27023 13484 27068 13512
rect 27062 13472 27068 13484
rect 27120 13472 27126 13524
rect 23658 13444 23664 13456
rect 22940 13416 23664 13444
rect 23658 13404 23664 13416
rect 23716 13404 23722 13456
rect 19978 13376 19984 13388
rect 18524 13348 19984 13376
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18524 13308 18552 13348
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 20070 13336 20076 13388
rect 20128 13376 20134 13388
rect 20714 13376 20720 13388
rect 20128 13348 20173 13376
rect 20627 13348 20720 13376
rect 20128 13336 20134 13348
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 22002 13376 22008 13388
rect 21963 13348 22008 13376
rect 22002 13336 22008 13348
rect 22060 13336 22066 13388
rect 25593 13379 25651 13385
rect 23860 13348 24624 13376
rect 18279 13280 18552 13308
rect 18693 13311 18751 13317
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 18693 13277 18705 13311
rect 18739 13277 18751 13311
rect 18874 13308 18880 13320
rect 18835 13280 18880 13308
rect 18693 13271 18751 13277
rect 17494 13240 17500 13252
rect 15856 13212 16896 13240
rect 17455 13212 17500 13240
rect 8076 13144 9536 13172
rect 8076 13132 8082 13144
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 11698 13172 11704 13184
rect 10284 13144 11704 13172
rect 10284 13132 10290 13144
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 11882 13172 11888 13184
rect 11843 13144 11888 13172
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12805 13175 12863 13181
rect 12805 13172 12817 13175
rect 12032 13144 12817 13172
rect 12032 13132 12038 13144
rect 12805 13141 12817 13144
rect 12851 13172 12863 13175
rect 14182 13172 14188 13184
rect 12851 13144 14188 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 15856 13172 15884 13212
rect 16022 13172 16028 13184
rect 14700 13144 15884 13172
rect 15983 13144 16028 13172
rect 14700 13132 14706 13144
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16868 13172 16896 13212
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18248 13172 18276 13271
rect 18708 13240 18736 13271
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 19484 13280 19809 13308
rect 19484 13268 19490 13280
rect 19797 13277 19809 13280
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 20732 13308 20760 13336
rect 19935 13280 20760 13308
rect 20809 13311 20867 13317
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20809 13277 20821 13311
rect 20855 13277 20867 13311
rect 23860 13308 23888 13348
rect 24026 13308 24032 13320
rect 20809 13271 20867 13277
rect 22204 13280 23888 13308
rect 23987 13280 24032 13308
rect 19518 13240 19524 13252
rect 18708 13212 19524 13240
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 20824 13240 20852 13271
rect 22204 13240 22232 13280
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 24596 13317 24624 13348
rect 25593 13345 25605 13379
rect 25639 13376 25651 13379
rect 26786 13376 26792 13388
rect 25639 13348 26792 13376
rect 25639 13345 25651 13348
rect 25593 13339 25651 13345
rect 26786 13336 26792 13348
rect 26844 13336 26850 13388
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13308 24639 13311
rect 25130 13308 25136 13320
rect 24627 13280 25136 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 25314 13308 25320 13320
rect 25275 13280 25320 13308
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 20824 13212 22232 13240
rect 22272 13243 22330 13249
rect 22272 13209 22284 13243
rect 22318 13240 22330 13243
rect 22318 13212 23888 13240
rect 22318 13209 22330 13212
rect 22272 13203 22330 13209
rect 16868 13144 18276 13172
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 18564 13144 18705 13172
rect 18564 13132 18570 13144
rect 18693 13141 18705 13144
rect 18739 13141 18751 13175
rect 18693 13135 18751 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 19392 13144 19441 13172
rect 19392 13132 19398 13144
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 20070 13132 20076 13184
rect 20128 13172 20134 13184
rect 22646 13172 22652 13184
rect 20128 13144 22652 13172
rect 20128 13132 20134 13144
rect 22646 13132 22652 13144
rect 22704 13132 22710 13184
rect 23860 13181 23888 13212
rect 26602 13200 26608 13252
rect 26660 13200 26666 13252
rect 23845 13175 23903 13181
rect 23845 13141 23857 13175
rect 23891 13141 23903 13175
rect 23845 13135 23903 13141
rect 1104 13082 28032 13104
rect 1104 13030 7642 13082
rect 7694 13030 7706 13082
rect 7758 13030 7770 13082
rect 7822 13030 7834 13082
rect 7886 13030 7898 13082
rect 7950 13030 14334 13082
rect 14386 13030 14398 13082
rect 14450 13030 14462 13082
rect 14514 13030 14526 13082
rect 14578 13030 14590 13082
rect 14642 13030 21026 13082
rect 21078 13030 21090 13082
rect 21142 13030 21154 13082
rect 21206 13030 21218 13082
rect 21270 13030 21282 13082
rect 21334 13030 27718 13082
rect 27770 13030 27782 13082
rect 27834 13030 27846 13082
rect 27898 13030 27910 13082
rect 27962 13030 27974 13082
rect 28026 13030 28032 13082
rect 1104 13008 28032 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 1854 12968 1860 12980
rect 1719 12940 1860 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 1946 12928 1952 12980
rect 2004 12968 2010 12980
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 2004 12940 3985 12968
rect 2004 12928 2010 12940
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 4246 12968 4252 12980
rect 3973 12931 4031 12937
rect 4080 12940 4252 12968
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 2774 12900 2780 12912
rect 2547 12872 2780 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 4080 12900 4108 12940
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 4764 12940 6561 12968
rect 4764 12928 4770 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 7098 12968 7104 12980
rect 6696 12940 7104 12968
rect 6696 12928 6702 12940
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 10318 12968 10324 12980
rect 10279 12940 10324 12968
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 11514 12968 11520 12980
rect 10560 12940 11520 12968
rect 10560 12928 10566 12940
rect 11514 12928 11520 12940
rect 11572 12968 11578 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11572 12940 11897 12968
rect 11572 12928 11578 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 11885 12931 11943 12937
rect 12897 12971 12955 12977
rect 12897 12937 12909 12971
rect 12943 12968 12955 12971
rect 13538 12968 13544 12980
rect 12943 12940 13544 12968
rect 12943 12937 12955 12940
rect 12897 12931 12955 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 13998 12968 14004 12980
rect 13771 12940 14004 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 13998 12928 14004 12940
rect 14056 12968 14062 12980
rect 16942 12968 16948 12980
rect 14056 12940 16948 12968
rect 14056 12928 14062 12940
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 17184 12940 17233 12968
rect 17184 12928 17190 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17221 12931 17279 12937
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 17368 12940 18245 12968
rect 17368 12928 17374 12940
rect 18233 12937 18245 12940
rect 18279 12937 18291 12971
rect 18233 12931 18291 12937
rect 19521 12971 19579 12977
rect 19521 12937 19533 12971
rect 19567 12968 19579 12971
rect 19610 12968 19616 12980
rect 19567 12940 19616 12968
rect 19567 12937 19579 12940
rect 19521 12931 19579 12937
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 19978 12928 19984 12980
rect 20036 12928 20042 12980
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 21358 12968 21364 12980
rect 21315 12940 21364 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 21910 12928 21916 12980
rect 21968 12968 21974 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 21968 12940 22017 12968
rect 21968 12928 21974 12940
rect 22005 12937 22017 12940
rect 22051 12937 22063 12971
rect 22005 12931 22063 12937
rect 22465 12971 22523 12977
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 23382 12968 23388 12980
rect 22511 12940 23388 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 25314 12928 25320 12980
rect 25372 12968 25378 12980
rect 25409 12971 25467 12977
rect 25409 12968 25421 12971
rect 25372 12940 25421 12968
rect 25372 12928 25378 12940
rect 25409 12937 25421 12940
rect 25455 12937 25467 12971
rect 25409 12931 25467 12937
rect 3726 12872 4108 12900
rect 4154 12860 4160 12912
rect 4212 12900 4218 12912
rect 4862 12903 4920 12909
rect 4862 12900 4874 12903
rect 4212 12872 4874 12900
rect 4212 12860 4218 12872
rect 4862 12869 4874 12872
rect 4908 12869 4920 12903
rect 4862 12863 4920 12869
rect 5258 12860 5264 12912
rect 5316 12900 5322 12912
rect 7837 12903 7895 12909
rect 7837 12900 7849 12903
rect 5316 12872 7849 12900
rect 5316 12860 5322 12872
rect 7837 12869 7849 12872
rect 7883 12900 7895 12903
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 7883 12872 10364 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 2222 12832 2228 12844
rect 2183 12804 2228 12832
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4706 12832 4712 12844
rect 4663 12804 4712 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12832 6975 12835
rect 7282 12832 7288 12844
rect 6963 12804 7288 12832
rect 6963 12801 6975 12804
rect 6917 12795 6975 12801
rect 7282 12792 7288 12804
rect 7340 12832 7346 12844
rect 9585 12835 9643 12841
rect 7340 12804 8800 12832
rect 7340 12792 7346 12804
rect 7009 12767 7067 12773
rect 7009 12764 7021 12767
rect 6932 12736 7021 12764
rect 6932 12708 6960 12736
rect 7009 12733 7021 12736
rect 7055 12733 7067 12767
rect 7009 12727 7067 12733
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12764 7251 12767
rect 7650 12764 7656 12776
rect 7239 12736 7656 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 6914 12656 6920 12708
rect 6972 12656 6978 12708
rect 8772 12696 8800 12804
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10226 12832 10232 12844
rect 9631 12804 10232 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10336 12841 10364 12872
rect 10428 12872 12112 12900
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 9674 12764 9680 12776
rect 9364 12736 9680 12764
rect 9364 12724 9370 12736
rect 9674 12724 9680 12736
rect 9732 12764 9738 12776
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 9732 12736 10149 12764
rect 9732 12724 9738 12736
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10137 12727 10195 12733
rect 10428 12696 10456 12872
rect 12084 12832 12112 12872
rect 13648 12872 13829 12900
rect 12434 12832 12440 12844
rect 12084 12804 12440 12832
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 12526 12792 12532 12844
rect 12584 12832 12590 12844
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12584 12804 12817 12832
rect 12584 12792 12590 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 13538 12832 13544 12844
rect 13228 12804 13544 12832
rect 13228 12792 13234 12804
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 12253 12767 12311 12773
rect 10735 12736 11744 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 11716 12705 11744 12736
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12710 12764 12716 12776
rect 12299 12736 12716 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 13648 12764 13676 12872
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 14093 12903 14151 12909
rect 14093 12869 14105 12903
rect 14139 12900 14151 12903
rect 14182 12900 14188 12912
rect 14139 12872 14188 12900
rect 14139 12869 14151 12872
rect 14093 12863 14151 12869
rect 14182 12860 14188 12872
rect 14240 12900 14246 12912
rect 15010 12900 15016 12912
rect 14240 12872 15016 12900
rect 14240 12860 14246 12872
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 15838 12860 15844 12912
rect 15896 12900 15902 12912
rect 16301 12903 16359 12909
rect 16301 12900 16313 12903
rect 15896 12872 16313 12900
rect 15896 12860 15902 12872
rect 16301 12869 16313 12872
rect 16347 12869 16359 12903
rect 16301 12863 16359 12869
rect 17402 12860 17408 12912
rect 17460 12900 17466 12912
rect 18138 12900 18144 12912
rect 17460 12872 18144 12900
rect 17460 12860 17466 12872
rect 18138 12860 18144 12872
rect 18196 12860 18202 12912
rect 18506 12900 18512 12912
rect 18467 12872 18512 12900
rect 18506 12860 18512 12872
rect 18564 12860 18570 12912
rect 18601 12903 18659 12909
rect 18601 12869 18613 12903
rect 18647 12900 18659 12903
rect 19702 12900 19708 12912
rect 18647 12872 19708 12900
rect 18647 12869 18659 12872
rect 18601 12863 18659 12869
rect 19702 12860 19708 12872
rect 19760 12860 19766 12912
rect 19996 12900 20024 12928
rect 23290 12900 23296 12912
rect 19996 12872 20852 12900
rect 23251 12872 23296 12900
rect 13722 12792 13728 12844
rect 13780 12832 13786 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13780 12804 13921 12832
rect 13780 12792 13786 12804
rect 13909 12801 13921 12804
rect 13955 12801 13967 12835
rect 13909 12795 13967 12801
rect 18412 12835 18470 12841
rect 18412 12801 18424 12835
rect 18458 12832 18470 12835
rect 18458 12804 18552 12832
rect 18458 12801 18470 12804
rect 18412 12795 18470 12801
rect 14550 12764 14556 12776
rect 13504 12736 13676 12764
rect 14511 12736 14556 12764
rect 13504 12724 13510 12736
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 8772 12668 10456 12696
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12665 11759 12699
rect 11701 12659 11759 12665
rect 17328 12640 17356 12727
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 17460 12736 17505 12764
rect 17460 12724 17466 12736
rect 18524 12696 18552 12804
rect 18690 12792 18696 12844
rect 18748 12841 18754 12844
rect 18748 12835 18787 12841
rect 18775 12801 18787 12835
rect 18748 12795 18787 12801
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12801 18935 12835
rect 19334 12832 19340 12844
rect 19295 12804 19340 12832
rect 18877 12795 18935 12801
rect 18748 12792 18754 12795
rect 18892 12764 18920 12795
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 20180 12841 20208 12872
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19852 12804 19993 12832
rect 19852 12792 19858 12804
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 20438 12792 20444 12844
rect 20496 12832 20502 12844
rect 20824 12841 20852 12872
rect 23290 12860 23296 12872
rect 23348 12860 23354 12912
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20496 12804 20637 12832
rect 20496 12792 20502 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12801 20867 12835
rect 21450 12832 21456 12844
rect 21411 12804 21456 12832
rect 20809 12795 20867 12801
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 22152 12804 22385 12832
rect 22152 12792 22158 12804
rect 22373 12801 22385 12804
rect 22419 12832 22431 12835
rect 23382 12832 23388 12844
rect 22419 12804 23388 12832
rect 22419 12801 22431 12804
rect 22373 12795 22431 12801
rect 23382 12792 23388 12804
rect 23440 12792 23446 12844
rect 25130 12792 25136 12844
rect 25188 12832 25194 12844
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 25188 12804 25421 12832
rect 25188 12792 25194 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 22462 12764 22468 12776
rect 18892 12736 22468 12764
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 22646 12764 22652 12776
rect 22607 12736 22652 12764
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 19058 12696 19064 12708
rect 18524 12668 19064 12696
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 5994 12628 6000 12640
rect 5955 12600 6000 12628
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10226 12628 10232 12640
rect 9824 12600 10232 12628
rect 9824 12588 9830 12600
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10870 12588 10876 12640
rect 10928 12628 10934 12640
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 10928 12600 11897 12628
rect 10928 12588 10934 12600
rect 11885 12597 11897 12600
rect 11931 12628 11943 12631
rect 12342 12628 12348 12640
rect 11931 12600 12348 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12986 12628 12992 12640
rect 12492 12600 12992 12628
rect 12492 12588 12498 12600
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 16724 12600 16865 12628
rect 16724 12588 16730 12600
rect 16853 12597 16865 12600
rect 16899 12597 16911 12631
rect 16853 12591 16911 12597
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 18874 12628 18880 12640
rect 17368 12600 18880 12628
rect 17368 12588 17374 12600
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 19024 12600 20085 12628
rect 19024 12588 19030 12600
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 20714 12628 20720 12640
rect 20675 12600 20720 12628
rect 20073 12591 20131 12597
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 23382 12588 23388 12640
rect 23440 12628 23446 12640
rect 23753 12631 23811 12637
rect 23753 12628 23765 12631
rect 23440 12600 23765 12628
rect 23440 12588 23446 12600
rect 23753 12597 23765 12600
rect 23799 12597 23811 12631
rect 23753 12591 23811 12597
rect 1104 12538 27876 12560
rect 1104 12486 4296 12538
rect 4348 12486 4360 12538
rect 4412 12486 4424 12538
rect 4476 12486 4488 12538
rect 4540 12486 4552 12538
rect 4604 12486 10988 12538
rect 11040 12486 11052 12538
rect 11104 12486 11116 12538
rect 11168 12486 11180 12538
rect 11232 12486 11244 12538
rect 11296 12486 17680 12538
rect 17732 12486 17744 12538
rect 17796 12486 17808 12538
rect 17860 12486 17872 12538
rect 17924 12486 17936 12538
rect 17988 12486 24372 12538
rect 24424 12486 24436 12538
rect 24488 12486 24500 12538
rect 24552 12486 24564 12538
rect 24616 12486 24628 12538
rect 24680 12486 27876 12538
rect 1104 12464 27876 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 6549 12427 6607 12433
rect 1995 12396 6132 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 5166 12356 5172 12368
rect 4448 12328 5172 12356
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12288 2651 12291
rect 4448 12288 4476 12328
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 6104 12356 6132 12396
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 6914 12424 6920 12436
rect 6595 12396 6920 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7009 12427 7067 12433
rect 7009 12393 7021 12427
rect 7055 12424 7067 12427
rect 7098 12424 7104 12436
rect 7055 12396 7104 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8386 12424 8392 12436
rect 8260 12396 8392 12424
rect 8260 12384 8266 12396
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 16758 12424 16764 12436
rect 10008 12396 12434 12424
rect 10008 12384 10014 12396
rect 9122 12356 9128 12368
rect 6104 12328 9128 12356
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 10594 12316 10600 12368
rect 10652 12356 10658 12368
rect 10652 12328 12296 12356
rect 10652 12316 10658 12328
rect 4614 12288 4620 12300
rect 2639 12260 4476 12288
rect 4575 12260 4620 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2832 12192 3065 12220
rect 2832 12180 2838 12192
rect 3053 12189 3065 12192
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 4448 12220 4476 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6972 12260 7481 12288
rect 6972 12248 6978 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7650 12288 7656 12300
rect 7611 12260 7656 12288
rect 7469 12251 7527 12257
rect 7650 12248 7656 12260
rect 7708 12288 7714 12300
rect 8110 12288 8116 12300
rect 7708 12260 8116 12288
rect 7708 12248 7714 12260
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 11330 12288 11336 12300
rect 9048 12260 11336 12288
rect 4387 12192 4476 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 1578 12112 1584 12164
rect 1636 12152 1642 12164
rect 1673 12155 1731 12161
rect 1673 12152 1685 12155
rect 1636 12124 1685 12152
rect 1636 12112 1642 12124
rect 1673 12121 1685 12124
rect 1719 12121 1731 12155
rect 1673 12115 1731 12121
rect 2038 12112 2044 12164
rect 2096 12152 2102 12164
rect 3252 12152 3280 12183
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 5166 12220 5172 12232
rect 4764 12192 5172 12220
rect 4764 12180 4770 12192
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 9048 12220 9076 12260
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11664 12260 12173 12288
rect 11664 12248 11670 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 5276 12192 9076 12220
rect 9125 12223 9183 12229
rect 2096 12124 3280 12152
rect 3421 12155 3479 12161
rect 2096 12112 2102 12124
rect 3421 12121 3433 12155
rect 3467 12152 3479 12155
rect 5276 12152 5304 12192
rect 9125 12189 9137 12223
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 5442 12161 5448 12164
rect 5436 12152 5448 12161
rect 3467 12124 5304 12152
rect 5403 12124 5448 12152
rect 3467 12121 3479 12124
rect 3421 12115 3479 12121
rect 5436 12115 5448 12124
rect 5442 12112 5448 12115
rect 5500 12112 5506 12164
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6638 12152 6644 12164
rect 6052 12124 6644 12152
rect 6052 12112 6058 12124
rect 6638 12112 6644 12124
rect 6696 12152 6702 12164
rect 6914 12152 6920 12164
rect 6696 12124 6920 12152
rect 6696 12112 6702 12124
rect 6914 12112 6920 12124
rect 6972 12112 6978 12164
rect 7377 12155 7435 12161
rect 7377 12152 7389 12155
rect 7024 12124 7389 12152
rect 3970 12084 3976 12096
rect 3931 12056 3976 12084
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4430 12084 4436 12096
rect 4391 12056 4436 12084
rect 4430 12044 4436 12056
rect 4488 12044 4494 12096
rect 4890 12044 4896 12096
rect 4948 12084 4954 12096
rect 7024 12084 7052 12124
rect 7377 12121 7389 12124
rect 7423 12121 7435 12155
rect 7377 12115 7435 12121
rect 8294 12112 8300 12164
rect 8352 12152 8358 12164
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 8352 12124 8401 12152
rect 8352 12112 8358 12124
rect 8389 12121 8401 12124
rect 8435 12121 8447 12155
rect 8570 12152 8576 12164
rect 8531 12124 8576 12152
rect 8389 12115 8447 12121
rect 4948 12056 7052 12084
rect 4948 12044 4954 12056
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7524 12056 8217 12084
rect 7524 12044 7530 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8404 12084 8432 12115
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 9140 12152 9168 12183
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 10744 12192 11989 12220
rect 10744 12180 10750 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 12268 12220 12296 12328
rect 12406 12288 12434 12396
rect 15028 12396 16764 12424
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 15028 12356 15056 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17310 12424 17316 12436
rect 17267 12396 17316 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 19058 12384 19064 12436
rect 19116 12424 19122 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19116 12396 19809 12424
rect 19116 12384 19122 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19797 12387 19855 12393
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 22520 12396 22845 12424
rect 22520 12384 22526 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 22833 12387 22891 12393
rect 13872 12328 15056 12356
rect 18432 12328 20668 12356
rect 13872 12316 13878 12328
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 12406 12260 13369 12288
rect 13357 12257 13369 12260
rect 13403 12257 13415 12291
rect 14734 12288 14740 12300
rect 14695 12260 14740 12288
rect 13357 12251 13415 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15286 12288 15292 12300
rect 15247 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 13906 12220 13912 12232
rect 12268 12192 13912 12220
rect 11977 12183 12035 12189
rect 13906 12180 13912 12192
rect 13964 12220 13970 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13964 12192 14565 12220
rect 13964 12180 13970 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12220 15899 12223
rect 15930 12220 15936 12232
rect 15887 12192 15936 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 18432 12220 18460 12328
rect 18506 12248 18512 12300
rect 18564 12288 18570 12300
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 18564 12260 18613 12288
rect 18564 12248 18570 12260
rect 18601 12257 18613 12260
rect 18647 12288 18659 12291
rect 18966 12288 18972 12300
rect 18647 12260 18972 12288
rect 18647 12257 18659 12260
rect 18601 12251 18659 12257
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 16040 12192 18460 12220
rect 9398 12152 9404 12164
rect 9088 12124 9168 12152
rect 9359 12124 9404 12152
rect 9088 12112 9094 12124
rect 9398 12112 9404 12124
rect 9456 12112 9462 12164
rect 10410 12112 10416 12164
rect 10468 12112 10474 12164
rect 11790 12112 11796 12164
rect 11848 12152 11854 12164
rect 12069 12155 12127 12161
rect 12069 12152 12081 12155
rect 11848 12124 12081 12152
rect 11848 12112 11854 12124
rect 12069 12121 12081 12124
rect 12115 12121 12127 12155
rect 12069 12115 12127 12121
rect 12618 12112 12624 12164
rect 12676 12152 12682 12164
rect 16040 12152 16068 12192
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 18932 12192 19441 12220
rect 18932 12180 18938 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 20640 12229 20668 12328
rect 23106 12288 23112 12300
rect 23067 12260 23112 12288
rect 23106 12248 23112 12260
rect 23164 12248 23170 12300
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19576 12192 19625 12220
rect 19576 12180 19582 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 21726 12220 21732 12232
rect 21687 12192 21732 12220
rect 20625 12183 20683 12189
rect 16114 12161 16120 12164
rect 12676 12124 16068 12152
rect 12676 12112 12682 12124
rect 13188 12096 13216 12124
rect 16108 12115 16120 12161
rect 16172 12152 16178 12164
rect 16172 12124 16208 12152
rect 16114 12112 16120 12115
rect 16172 12112 16178 12124
rect 17126 12112 17132 12164
rect 17184 12152 17190 12164
rect 18417 12155 18475 12161
rect 18417 12152 18429 12155
rect 17184 12124 18429 12152
rect 17184 12112 17190 12124
rect 18417 12121 18429 12124
rect 18463 12152 18475 12155
rect 19334 12152 19340 12164
rect 18463 12124 19340 12152
rect 18463 12121 18475 12124
rect 18417 12115 18475 12121
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 20640 12152 20668 12183
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 23198 12220 23204 12232
rect 23159 12192 23204 12220
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 23845 12155 23903 12161
rect 23845 12152 23857 12155
rect 20640 12124 23857 12152
rect 23845 12121 23857 12124
rect 23891 12121 23903 12155
rect 23845 12115 23903 12121
rect 10778 12084 10784 12096
rect 8404 12056 10784 12084
rect 8205 12047 8263 12053
rect 10778 12044 10784 12056
rect 10836 12084 10842 12096
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 10836 12056 10885 12084
rect 10836 12044 10842 12056
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 10873 12047 10931 12053
rect 11609 12087 11667 12093
rect 11609 12053 11621 12087
rect 11655 12084 11667 12087
rect 11698 12084 11704 12096
rect 11655 12056 11704 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12584 12056 12817 12084
rect 12584 12044 12590 12056
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 12805 12047 12863 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13630 12084 13636 12096
rect 13311 12056 13636 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 18046 12084 18052 12096
rect 18007 12056 18052 12084
rect 18046 12044 18052 12056
rect 18104 12044 18110 12096
rect 18509 12087 18567 12093
rect 18509 12053 18521 12087
rect 18555 12084 18567 12087
rect 18966 12084 18972 12096
rect 18555 12056 18972 12084
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 20809 12087 20867 12093
rect 20809 12084 20821 12087
rect 20496 12056 20821 12084
rect 20496 12044 20502 12056
rect 20809 12053 20821 12056
rect 20855 12053 20867 12087
rect 21910 12084 21916 12096
rect 21871 12056 21916 12084
rect 20809 12047 20867 12053
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 1104 11994 28032 12016
rect 1104 11942 7642 11994
rect 7694 11942 7706 11994
rect 7758 11942 7770 11994
rect 7822 11942 7834 11994
rect 7886 11942 7898 11994
rect 7950 11942 14334 11994
rect 14386 11942 14398 11994
rect 14450 11942 14462 11994
rect 14514 11942 14526 11994
rect 14578 11942 14590 11994
rect 14642 11942 21026 11994
rect 21078 11942 21090 11994
rect 21142 11942 21154 11994
rect 21206 11942 21218 11994
rect 21270 11942 21282 11994
rect 21334 11942 27718 11994
rect 27770 11942 27782 11994
rect 27834 11942 27846 11994
rect 27898 11942 27910 11994
rect 27962 11942 27974 11994
rect 28026 11942 28032 11994
rect 1104 11920 28032 11942
rect 2225 11883 2283 11889
rect 2225 11849 2237 11883
rect 2271 11880 2283 11883
rect 4065 11883 4123 11889
rect 2271 11852 2774 11880
rect 2271 11849 2283 11852
rect 2225 11843 2283 11849
rect 2746 11812 2774 11852
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4430 11880 4436 11892
rect 4111 11852 4436 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4430 11840 4436 11852
rect 4488 11880 4494 11892
rect 7926 11880 7932 11892
rect 4488 11852 5304 11880
rect 4488 11840 4494 11852
rect 2930 11815 2988 11821
rect 2930 11812 2942 11815
rect 2746 11784 2942 11812
rect 2930 11781 2942 11784
rect 2976 11781 2988 11815
rect 2930 11775 2988 11781
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 4672 11784 5212 11812
rect 4672 11772 4678 11784
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 3970 11744 3976 11756
rect 2087 11716 3976 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 4890 11744 4896 11756
rect 4851 11716 4896 11744
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11645 2743 11679
rect 4982 11676 4988 11688
rect 4943 11648 4988 11676
rect 2685 11639 2743 11645
rect 2700 11540 2728 11639
rect 4982 11636 4988 11648
rect 5040 11636 5046 11688
rect 5184 11685 5212 11784
rect 5276 11744 5304 11852
rect 5920 11852 7932 11880
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 5920 11812 5948 11852
rect 7926 11840 7932 11852
rect 7984 11880 7990 11892
rect 10410 11880 10416 11892
rect 7984 11852 10088 11880
rect 10371 11852 10416 11880
rect 7984 11840 7990 11852
rect 7006 11812 7012 11824
rect 5500 11784 5948 11812
rect 6840 11784 7012 11812
rect 5500 11772 5506 11784
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5276 11716 5825 11744
rect 5813 11713 5825 11716
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6362 11744 6368 11756
rect 6043 11716 6368 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 5169 11679 5227 11685
rect 5169 11645 5181 11679
rect 5215 11676 5227 11679
rect 5828 11676 5856 11707
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6512 11716 6745 11744
rect 6512 11704 6518 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6546 11676 6552 11688
rect 5215 11648 5304 11676
rect 5828 11648 6552 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 4706 11608 4712 11620
rect 3620 11580 4712 11608
rect 2866 11540 2872 11552
rect 2700 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11540 2930 11552
rect 3620 11540 3648 11580
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 2924 11512 3648 11540
rect 2924 11500 2930 11512
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4212 11512 4537 11540
rect 4212 11500 4218 11512
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 5276 11540 5304 11648
rect 6546 11636 6552 11648
rect 6604 11636 6610 11688
rect 6840 11685 6868 11784
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 7466 11772 7472 11824
rect 7524 11812 7530 11824
rect 7524 11784 7788 11812
rect 7524 11772 7530 11784
rect 7760 11753 7788 11784
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 8021 11815 8079 11821
rect 8021 11812 8033 11815
rect 7892 11784 8033 11812
rect 7892 11772 7898 11784
rect 8021 11781 8033 11784
rect 8067 11781 8079 11815
rect 8846 11812 8852 11824
rect 8807 11784 8852 11812
rect 8021 11775 8079 11781
rect 8846 11772 8852 11784
rect 8904 11772 8910 11824
rect 9950 11812 9956 11824
rect 9508 11784 9956 11812
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7116 11716 7665 11744
rect 7116 11685 7144 11716
rect 7653 11713 7665 11716
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 7746 11747 7804 11753
rect 7746 11713 7758 11747
rect 7792 11713 7804 11747
rect 7746 11707 7804 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8118 11747 8176 11753
rect 8118 11713 8130 11747
rect 8164 11713 8176 11747
rect 9508 11744 9536 11784
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10060 11812 10088 11852
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 11790 11840 11796 11892
rect 11848 11880 11854 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 11848 11852 13093 11880
rect 11848 11840 11854 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13081 11843 13139 11849
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 15010 11880 15016 11892
rect 14507 11852 15016 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 15194 11880 15200 11892
rect 15155 11852 15200 11880
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 16114 11880 16120 11892
rect 16071 11852 16120 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 18966 11880 18972 11892
rect 18927 11852 18972 11880
rect 18966 11840 18972 11852
rect 19024 11880 19030 11892
rect 19024 11852 19472 11880
rect 19024 11840 19030 11852
rect 10686 11812 10692 11824
rect 10060 11784 10692 11812
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 12434 11812 12440 11824
rect 11164 11784 12440 11812
rect 8118 11707 8176 11713
rect 8220 11716 9536 11744
rect 9769 11747 9827 11753
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 7944 11676 7972 11707
rect 7616 11648 7972 11676
rect 7616 11636 7622 11648
rect 5905 11611 5963 11617
rect 5905 11577 5917 11611
rect 5951 11608 5963 11611
rect 8128 11608 8156 11707
rect 5951 11580 8156 11608
rect 5951 11577 5963 11580
rect 5905 11571 5963 11577
rect 8220 11540 8248 11716
rect 9769 11713 9781 11747
rect 9815 11744 9827 11747
rect 10226 11744 10232 11756
rect 9815 11716 10232 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10226 11704 10232 11716
rect 10284 11744 10290 11756
rect 10594 11744 10600 11756
rect 10284 11716 10600 11744
rect 10284 11704 10290 11716
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11164 11753 11192 11784
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 14553 11815 14611 11821
rect 14553 11781 14565 11815
rect 14599 11812 14611 11815
rect 14918 11812 14924 11824
rect 14599 11784 14924 11812
rect 14599 11781 14611 11784
rect 14553 11775 14611 11781
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 17586 11772 17592 11824
rect 17644 11812 17650 11824
rect 19444 11821 19472 11852
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 19797 11883 19855 11889
rect 19797 11880 19809 11883
rect 19760 11852 19809 11880
rect 19760 11840 19766 11852
rect 19797 11849 19809 11852
rect 19843 11849 19855 11883
rect 19797 11843 19855 11849
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 20257 11883 20315 11889
rect 20257 11880 20269 11883
rect 20220 11852 20269 11880
rect 20220 11840 20226 11852
rect 20257 11849 20269 11852
rect 20303 11849 20315 11883
rect 20257 11843 20315 11849
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 22738 11880 22744 11892
rect 20496 11852 22744 11880
rect 20496 11840 20502 11852
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 17834 11815 17892 11821
rect 17834 11812 17846 11815
rect 17644 11784 17846 11812
rect 17644 11772 17650 11784
rect 17834 11781 17846 11784
rect 17880 11781 17892 11815
rect 17834 11775 17892 11781
rect 19429 11815 19487 11821
rect 19429 11781 19441 11815
rect 19475 11781 19487 11815
rect 19429 11775 19487 11781
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 22250 11815 22308 11821
rect 22250 11812 22262 11815
rect 21968 11784 22262 11812
rect 21968 11772 21974 11784
rect 22250 11781 22262 11784
rect 22296 11781 22308 11815
rect 22250 11775 22308 11781
rect 11974 11753 11980 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10928 11716 10977 11744
rect 10928 11704 10934 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11968 11707 11980 11753
rect 12032 11744 12038 11756
rect 12032 11716 12068 11744
rect 11974 11704 11980 11707
rect 12032 11704 12038 11716
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 12400 11716 13553 11744
rect 12400 11704 12406 11716
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13814 11744 13820 11756
rect 13775 11716 13820 11744
rect 13541 11707 13599 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 15378 11744 15384 11756
rect 15291 11716 15384 11744
rect 15378 11704 15384 11716
rect 15436 11744 15442 11756
rect 16022 11744 16028 11756
rect 15436 11716 16028 11744
rect 15436 11704 15442 11716
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11744 16267 11747
rect 16666 11744 16672 11756
rect 16255 11716 16672 11744
rect 16255 11713 16267 11716
rect 16209 11707 16267 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 16850 11744 16856 11756
rect 16811 11716 16856 11744
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 17678 11744 17684 11756
rect 17368 11716 17684 11744
rect 17368 11704 17374 11716
rect 17678 11704 17684 11716
rect 17736 11744 17742 11756
rect 17736 11716 18644 11744
rect 17736 11704 17742 11716
rect 8294 11636 8300 11688
rect 8352 11636 8358 11688
rect 9674 11676 9680 11688
rect 9635 11648 9680 11676
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11572 11648 11713 11676
rect 11572 11636 11578 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 13998 11676 14004 11688
rect 13955 11648 14004 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 13998 11636 14004 11648
rect 14056 11676 14062 11688
rect 15286 11676 15292 11688
rect 14056 11648 15292 11676
rect 14056 11636 14062 11648
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 17494 11636 17500 11688
rect 17552 11676 17558 11688
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 17552 11648 17601 11676
rect 17552 11636 17558 11648
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 18616 11676 18644 11716
rect 18782 11704 18788 11756
rect 18840 11744 18846 11756
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 18840 11716 19625 11744
rect 18840 11704 18846 11716
rect 19613 11713 19625 11716
rect 19659 11744 19671 11747
rect 22554 11744 22560 11756
rect 19659 11716 22560 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 23198 11704 23204 11756
rect 23256 11744 23262 11756
rect 24397 11747 24455 11753
rect 24397 11744 24409 11747
rect 23256 11716 24409 11744
rect 23256 11704 23262 11716
rect 24397 11713 24409 11716
rect 24443 11744 24455 11747
rect 26326 11744 26332 11756
rect 24443 11716 26332 11744
rect 24443 11713 24455 11716
rect 24397 11707 24455 11713
rect 26326 11704 26332 11716
rect 26384 11704 26390 11756
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 18616 11648 22017 11676
rect 17589 11639 17647 11645
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 8312 11608 8340 11636
rect 11057 11611 11115 11617
rect 11057 11608 11069 11611
rect 8312 11580 11069 11608
rect 11057 11577 11069 11580
rect 11103 11608 11115 11611
rect 11606 11608 11612 11620
rect 11103 11580 11612 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 19702 11608 19708 11620
rect 18892 11580 19708 11608
rect 5276 11512 8248 11540
rect 8297 11543 8355 11549
rect 4525 11503 4583 11509
rect 8297 11509 8309 11543
rect 8343 11540 8355 11543
rect 9214 11540 9220 11552
rect 8343 11512 9220 11540
rect 8343 11509 8355 11512
rect 8297 11503 8355 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11540 17095 11543
rect 18892 11540 18920 11580
rect 19702 11568 19708 11580
rect 19760 11568 19766 11620
rect 20438 11568 20444 11620
rect 20496 11608 20502 11620
rect 21361 11611 21419 11617
rect 21361 11608 21373 11611
rect 20496 11580 21373 11608
rect 20496 11568 20502 11580
rect 21361 11577 21373 11580
rect 21407 11577 21419 11611
rect 21361 11571 21419 11577
rect 17083 11512 18920 11540
rect 17083 11509 17095 11512
rect 17037 11503 17095 11509
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 20809 11543 20867 11549
rect 20809 11540 20821 11543
rect 20680 11512 20821 11540
rect 20680 11500 20686 11512
rect 20809 11509 20821 11512
rect 20855 11509 20867 11543
rect 20809 11503 20867 11509
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 23106 11540 23112 11552
rect 22244 11512 23112 11540
rect 22244 11500 22250 11512
rect 23106 11500 23112 11512
rect 23164 11540 23170 11552
rect 23385 11543 23443 11549
rect 23385 11540 23397 11543
rect 23164 11512 23397 11540
rect 23164 11500 23170 11512
rect 23385 11509 23397 11512
rect 23431 11509 23443 11543
rect 23385 11503 23443 11509
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 24854 11540 24860 11552
rect 24443 11512 24860 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 24854 11500 24860 11512
rect 24912 11500 24918 11552
rect 1104 11450 27876 11472
rect 1104 11398 4296 11450
rect 4348 11398 4360 11450
rect 4412 11398 4424 11450
rect 4476 11398 4488 11450
rect 4540 11398 4552 11450
rect 4604 11398 10988 11450
rect 11040 11398 11052 11450
rect 11104 11398 11116 11450
rect 11168 11398 11180 11450
rect 11232 11398 11244 11450
rect 11296 11398 17680 11450
rect 17732 11398 17744 11450
rect 17796 11398 17808 11450
rect 17860 11398 17872 11450
rect 17924 11398 17936 11450
rect 17988 11398 24372 11450
rect 24424 11398 24436 11450
rect 24488 11398 24500 11450
rect 24552 11398 24564 11450
rect 24616 11398 24628 11450
rect 24680 11398 27876 11450
rect 1104 11376 27876 11398
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 4982 11336 4988 11348
rect 3467 11308 4988 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 7285 11339 7343 11345
rect 5224 11308 7236 11336
rect 5224 11296 5230 11308
rect 4709 11271 4767 11277
rect 4709 11237 4721 11271
rect 4755 11237 4767 11271
rect 4709 11231 4767 11237
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4614 11200 4620 11212
rect 4203 11172 4620 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 4724 11200 4752 11231
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 6273 11271 6331 11277
rect 6273 11268 6285 11271
rect 4856 11240 6285 11268
rect 4856 11228 4862 11240
rect 6273 11237 6285 11240
rect 6319 11237 6331 11271
rect 6273 11231 6331 11237
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 6420 11240 6592 11268
rect 6420 11228 6426 11240
rect 4724 11172 6500 11200
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2866 11132 2872 11144
rect 2087 11104 2872 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 5074 11132 5080 11144
rect 4387 11104 5080 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 5074 11092 5080 11104
rect 5132 11092 5138 11144
rect 6472 11141 6500 11172
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11132 5871 11135
rect 6457 11135 6515 11141
rect 5859 11104 6408 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2286 11067 2344 11073
rect 2286 11064 2298 11067
rect 2188 11036 2298 11064
rect 2188 11024 2194 11036
rect 2286 11033 2298 11036
rect 2332 11033 2344 11067
rect 4246 11064 4252 11076
rect 4207 11036 4252 11064
rect 2286 11027 2344 11033
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 5626 10996 5632 11008
rect 5587 10968 5632 10996
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 6380 10996 6408 11104
rect 6457 11101 6469 11135
rect 6503 11101 6515 11135
rect 6564 11132 6592 11240
rect 6822 11132 6828 11144
rect 6564 11104 6828 11132
rect 6457 11095 6515 11101
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6880 11104 7113 11132
rect 6880 11092 6886 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6604 11036 6929 11064
rect 6604 11024 6610 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 7208 11064 7236 11308
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7742 11336 7748 11348
rect 7331 11308 7748 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 17126 11336 17132 11348
rect 17087 11308 17132 11336
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 17586 11296 17592 11348
rect 17644 11336 17650 11348
rect 17865 11339 17923 11345
rect 17865 11336 17877 11339
rect 17644 11308 17877 11336
rect 17644 11296 17650 11308
rect 17865 11305 17877 11308
rect 17911 11305 17923 11339
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 17865 11299 17923 11305
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 19981 11339 20039 11345
rect 19981 11336 19993 11339
rect 19392 11308 19993 11336
rect 19392 11296 19398 11308
rect 19981 11305 19993 11308
rect 20027 11336 20039 11339
rect 20622 11336 20628 11348
rect 20027 11308 20628 11336
rect 20027 11305 20039 11308
rect 19981 11299 20039 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21726 11336 21732 11348
rect 21687 11308 21732 11336
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 22738 11296 22744 11348
rect 22796 11336 22802 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22796 11308 22937 11336
rect 22796 11296 22802 11308
rect 22925 11305 22937 11308
rect 22971 11305 22983 11339
rect 22925 11299 22983 11305
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 23477 11339 23535 11345
rect 23477 11336 23489 11339
rect 23348 11308 23489 11336
rect 23348 11296 23354 11308
rect 23477 11305 23489 11308
rect 23523 11305 23535 11339
rect 26326 11336 26332 11348
rect 26287 11308 26332 11336
rect 23477 11299 23535 11305
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 7432 11240 7849 11268
rect 7432 11228 7438 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 9214 11268 9220 11280
rect 9175 11240 9220 11268
rect 7837 11231 7895 11237
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9490 11228 9496 11280
rect 9548 11268 9554 11280
rect 16485 11271 16543 11277
rect 9548 11240 12296 11268
rect 9548 11228 9554 11240
rect 8386 11200 8392 11212
rect 8220 11172 8392 11200
rect 8220 11141 8248 11172
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 10134 11200 10140 11212
rect 8527 11172 10140 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 12268 11209 12296 11240
rect 16485 11237 16497 11271
rect 16531 11237 16543 11271
rect 16485 11231 16543 11237
rect 22066 11240 22416 11268
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11169 12311 11203
rect 16500 11200 16528 11231
rect 18966 11200 18972 11212
rect 12253 11163 12311 11169
rect 15948 11172 16528 11200
rect 18616 11172 18972 11200
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 8570 11132 8576 11144
rect 8343 11104 8576 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 9122 11132 9128 11144
rect 9083 11104 9128 11132
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9490 11132 9496 11144
rect 9232 11104 9496 11132
rect 8478 11064 8484 11076
rect 7208 11036 8484 11064
rect 6917 11027 6975 11033
rect 8478 11024 8484 11036
rect 8536 11064 8542 11076
rect 9232 11064 9260 11104
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 10318 11132 10324 11144
rect 10091 11104 10324 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 15769 11135 15827 11141
rect 12406 11104 12664 11132
rect 8536 11036 9260 11064
rect 9401 11067 9459 11073
rect 8536 11024 8542 11036
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 12406 11064 12434 11104
rect 9447 11036 12434 11064
rect 12520 11067 12578 11073
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 12520 11033 12532 11067
rect 12566 11033 12578 11067
rect 12636 11064 12664 11104
rect 15769 11101 15781 11135
rect 15815 11132 15827 11135
rect 15948 11132 15976 11172
rect 15815 11104 15976 11132
rect 16025 11135 16083 11141
rect 15815 11101 15827 11104
rect 15769 11095 15827 11101
rect 16025 11101 16037 11135
rect 16071 11101 16083 11135
rect 16666 11132 16672 11144
rect 16627 11104 16672 11132
rect 16025 11095 16083 11101
rect 12710 11064 12716 11076
rect 12636 11036 12716 11064
rect 12520 11027 12578 11033
rect 7006 10996 7012 11008
rect 6380 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 11330 10996 11336 11008
rect 11291 10968 11336 10996
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12544 10996 12572 11027
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 14568 11036 14964 11064
rect 13630 10996 13636 11008
rect 12492 10968 12572 10996
rect 13591 10968 13636 10996
rect 12492 10956 12498 10968
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14568 10996 14596 11036
rect 14148 10968 14596 10996
rect 14645 10999 14703 11005
rect 14148 10956 14154 10968
rect 14645 10965 14657 10999
rect 14691 10996 14703 10999
rect 14826 10996 14832 11008
rect 14691 10968 14832 10996
rect 14691 10965 14703 10968
rect 14645 10959 14703 10965
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 14936 10996 14964 11036
rect 15930 11024 15936 11076
rect 15988 11064 15994 11076
rect 16040 11064 16068 11095
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18616 11141 18644 11172
rect 18966 11160 18972 11172
rect 19024 11160 19030 11212
rect 20714 11200 20720 11212
rect 20675 11172 20720 11200
rect 20714 11160 20720 11172
rect 20772 11200 20778 11212
rect 22066 11200 22094 11240
rect 22186 11200 22192 11212
rect 20772 11172 22094 11200
rect 22147 11172 22192 11200
rect 20772 11160 20778 11172
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 22388 11209 22416 11240
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 23106 11200 23112 11212
rect 22419 11172 23112 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 24854 11200 24860 11212
rect 24815 11172 24860 11200
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11101 18659 11135
rect 18782 11132 18788 11144
rect 18743 11104 18788 11132
rect 18601 11095 18659 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 20162 11132 20168 11144
rect 19352 11104 20168 11132
rect 17310 11064 17316 11076
rect 15988 11036 17316 11064
rect 15988 11024 15994 11036
rect 17310 11024 17316 11036
rect 17368 11024 17374 11076
rect 19352 10996 19380 11104
rect 20162 11092 20168 11104
rect 20220 11092 20226 11144
rect 20809 11135 20867 11141
rect 20809 11101 20821 11135
rect 20855 11132 20867 11135
rect 22094 11132 22100 11144
rect 20855 11104 22100 11132
rect 20855 11101 20867 11104
rect 20809 11095 20867 11101
rect 22094 11092 22100 11104
rect 22152 11092 22158 11144
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 19521 11067 19579 11073
rect 19521 11033 19533 11067
rect 19567 11064 19579 11067
rect 19610 11064 19616 11076
rect 19567 11036 19616 11064
rect 19567 11033 19579 11036
rect 19521 11027 19579 11033
rect 19610 11024 19616 11036
rect 19668 11064 19674 11076
rect 20438 11064 20444 11076
rect 19668 11036 20444 11064
rect 19668 11024 19674 11036
rect 20438 11024 20444 11036
rect 20496 11064 20502 11076
rect 20901 11067 20959 11073
rect 20901 11064 20913 11067
rect 20496 11036 20913 11064
rect 20496 11024 20502 11036
rect 20901 11033 20913 11036
rect 20947 11033 20959 11067
rect 23290 11064 23296 11076
rect 20901 11027 20959 11033
rect 21008 11036 23296 11064
rect 14936 10968 19380 10996
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 21008 10996 21036 11036
rect 19852 10968 21036 10996
rect 21269 10999 21327 11005
rect 19852 10956 19858 10968
rect 21269 10965 21281 10999
rect 21315 10996 21327 10999
rect 21358 10996 21364 11008
rect 21315 10968 21364 10996
rect 21315 10965 21327 10968
rect 21269 10959 21327 10965
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 22112 11005 22140 11036
rect 23290 11024 23296 11036
rect 23348 11024 23354 11076
rect 24596 11064 24624 11095
rect 24762 11064 24768 11076
rect 24596 11036 24768 11064
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 24946 11024 24952 11076
rect 25004 11064 25010 11076
rect 25004 11036 25346 11064
rect 25004 11024 25010 11036
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10965 22155 10999
rect 22097 10959 22155 10965
rect 1104 10906 28032 10928
rect 1104 10854 7642 10906
rect 7694 10854 7706 10906
rect 7758 10854 7770 10906
rect 7822 10854 7834 10906
rect 7886 10854 7898 10906
rect 7950 10854 14334 10906
rect 14386 10854 14398 10906
rect 14450 10854 14462 10906
rect 14514 10854 14526 10906
rect 14578 10854 14590 10906
rect 14642 10854 21026 10906
rect 21078 10854 21090 10906
rect 21142 10854 21154 10906
rect 21206 10854 21218 10906
rect 21270 10854 21282 10906
rect 21334 10854 27718 10906
rect 27770 10854 27782 10906
rect 27834 10854 27846 10906
rect 27898 10854 27910 10906
rect 27962 10854 27974 10906
rect 28026 10854 28032 10906
rect 1104 10832 28032 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 9674 10792 9680 10804
rect 8343 10764 9680 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11974 10792 11980 10804
rect 11931 10764 11980 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12345 10795 12403 10801
rect 12345 10761 12357 10795
rect 12391 10792 12403 10795
rect 12434 10792 12440 10804
rect 12391 10764 12440 10792
rect 12391 10761 12403 10764
rect 12345 10755 12403 10761
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 13906 10792 13912 10804
rect 13867 10764 13912 10792
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 15841 10795 15899 10801
rect 15841 10761 15853 10795
rect 15887 10792 15899 10795
rect 16666 10792 16672 10804
rect 15887 10764 16672 10792
rect 15887 10761 15899 10764
rect 15841 10755 15899 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 20441 10795 20499 10801
rect 20441 10761 20453 10795
rect 20487 10761 20499 10795
rect 20441 10755 20499 10761
rect 2860 10727 2918 10733
rect 2860 10693 2872 10727
rect 2906 10724 2918 10727
rect 4798 10724 4804 10736
rect 2906 10696 4804 10724
rect 2906 10693 2918 10696
rect 2860 10687 2918 10693
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 6914 10724 6920 10736
rect 5184 10696 6920 10724
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 4154 10656 4160 10668
rect 1995 10628 4160 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 5184 10665 5212 10696
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 10318 10724 10324 10736
rect 9631 10696 10324 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 10318 10684 10324 10696
rect 10376 10724 10382 10736
rect 11330 10724 11336 10736
rect 10376 10696 11336 10724
rect 10376 10684 10382 10696
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14461 10727 14519 10733
rect 14461 10724 14473 10727
rect 14148 10696 14473 10724
rect 14148 10684 14154 10696
rect 14461 10693 14473 10696
rect 14507 10693 14519 10727
rect 18325 10727 18383 10733
rect 18325 10724 18337 10727
rect 14461 10687 14519 10693
rect 15488 10696 18337 10724
rect 15488 10668 15516 10696
rect 18325 10693 18337 10696
rect 18371 10724 18383 10727
rect 19610 10724 19616 10736
rect 18371 10696 19616 10724
rect 18371 10693 18383 10696
rect 18325 10687 18383 10693
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 20456 10724 20484 10755
rect 20530 10752 20536 10804
rect 20588 10792 20594 10804
rect 24946 10792 24952 10804
rect 20588 10764 24072 10792
rect 24907 10764 24952 10792
rect 20588 10752 20594 10764
rect 22250 10727 22308 10733
rect 22250 10724 22262 10727
rect 20456 10696 22262 10724
rect 22250 10693 22262 10696
rect 22296 10693 22308 10727
rect 22250 10687 22308 10693
rect 24044 10724 24072 10764
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 25314 10724 25320 10736
rect 24044 10696 25320 10724
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 8110 10656 8116 10668
rect 6779 10628 8116 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 9766 10656 9772 10668
rect 8220 10628 9772 10656
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10557 2651 10591
rect 2593 10551 2651 10557
rect 2608 10452 2636 10551
rect 4982 10548 4988 10600
rect 5040 10588 5046 10600
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 5040 10560 5089 10588
rect 5040 10548 5046 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 6638 10588 6644 10600
rect 6599 10560 6644 10588
rect 5077 10551 5135 10557
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 8220 10532 8248 10628
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 10042 10656 10048 10668
rect 9955 10628 10048 10656
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9968 10588 9996 10628
rect 10042 10616 10048 10628
rect 10100 10656 10106 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10100 10628 10425 10656
rect 10100 10616 10106 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 11698 10656 11704 10668
rect 11659 10628 11704 10656
rect 10413 10619 10471 10625
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 12526 10656 12532 10668
rect 12487 10628 12532 10656
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 10134 10588 10140 10600
rect 9732 10560 9996 10588
rect 10095 10560 10140 10588
rect 9732 10548 9738 10560
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 4525 10523 4583 10529
rect 4525 10489 4537 10523
rect 4571 10520 4583 10523
rect 8202 10520 8208 10532
rect 4571 10492 8208 10520
rect 4571 10489 4583 10492
rect 4525 10483 4583 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10336 10520 10364 10551
rect 12158 10548 12164 10600
rect 12216 10588 12222 10600
rect 13188 10588 13216 10619
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14884 10628 15393 10656
rect 14884 10616 14890 10628
rect 15381 10625 15393 10628
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 15470 10616 15476 10668
rect 15528 10656 15534 10668
rect 17310 10656 17316 10668
rect 15528 10628 15573 10656
rect 17271 10628 17316 10656
rect 15528 10616 15534 10628
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 19518 10656 19524 10668
rect 19479 10628 19524 10656
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 20254 10656 20260 10668
rect 20215 10628 20260 10656
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 21085 10659 21143 10665
rect 21085 10625 21097 10659
rect 21131 10656 21143 10659
rect 21358 10656 21364 10668
rect 21131 10628 21364 10656
rect 21131 10625 21143 10628
rect 21085 10619 21143 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 24044 10656 24072 10696
rect 25314 10684 25320 10696
rect 25372 10724 25378 10736
rect 25409 10727 25467 10733
rect 25409 10724 25421 10727
rect 25372 10696 25421 10724
rect 25372 10684 25378 10696
rect 25409 10693 25421 10696
rect 25455 10693 25467 10727
rect 25409 10687 25467 10693
rect 24121 10659 24179 10665
rect 24121 10656 24133 10659
rect 24044 10628 24133 10656
rect 24121 10625 24133 10628
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25130 10656 25136 10668
rect 24627 10628 25136 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25130 10616 25136 10628
rect 25188 10616 25194 10668
rect 15286 10588 15292 10600
rect 12216 10560 13216 10588
rect 15247 10560 15292 10588
rect 12216 10548 12222 10560
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 17494 10588 17500 10600
rect 17455 10560 17500 10588
rect 17494 10548 17500 10560
rect 17552 10548 17558 10600
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18506 10548 18512 10600
rect 18564 10588 18570 10600
rect 18564 10560 18609 10588
rect 18564 10548 18570 10560
rect 14090 10520 14096 10532
rect 9824 10492 10364 10520
rect 10704 10492 14096 10520
rect 9824 10480 9830 10492
rect 2866 10452 2872 10464
rect 2608 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 3973 10455 4031 10461
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 4246 10452 4252 10464
rect 4019 10424 4252 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4246 10412 4252 10424
rect 4304 10452 4310 10464
rect 4614 10452 4620 10464
rect 4304 10424 4620 10452
rect 4304 10412 4310 10424
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 7101 10455 7159 10461
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 7650 10452 7656 10464
rect 7147 10424 7656 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 10042 10412 10048 10464
rect 10100 10452 10106 10464
rect 10704 10452 10732 10492
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10520 14703 10523
rect 15194 10520 15200 10532
rect 14691 10492 15200 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 15194 10480 15200 10492
rect 15252 10520 15258 10532
rect 15930 10520 15936 10532
rect 15252 10492 15936 10520
rect 15252 10480 15258 10492
rect 15930 10480 15936 10492
rect 15988 10480 15994 10532
rect 16758 10480 16764 10532
rect 16816 10520 16822 10532
rect 17957 10523 18015 10529
rect 17957 10520 17969 10523
rect 16816 10492 17969 10520
rect 16816 10480 16822 10492
rect 17957 10489 17969 10492
rect 18003 10489 18015 10523
rect 17957 10483 18015 10489
rect 10100 10424 10732 10452
rect 10781 10455 10839 10461
rect 10100 10412 10106 10424
rect 10781 10421 10793 10455
rect 10827 10452 10839 10455
rect 11330 10452 11336 10464
rect 10827 10424 11336 10452
rect 10827 10421 10839 10424
rect 10781 10415 10839 10421
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 19337 10455 19395 10461
rect 19337 10421 19349 10455
rect 19383 10452 19395 10455
rect 19426 10452 19432 10464
rect 19383 10424 19432 10452
rect 19383 10421 19395 10424
rect 19337 10415 19395 10421
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 20901 10455 20959 10461
rect 20901 10421 20913 10455
rect 20947 10452 20959 10455
rect 20990 10452 20996 10464
rect 20947 10424 20996 10452
rect 20947 10421 20959 10424
rect 20901 10415 20959 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 23290 10412 23296 10464
rect 23348 10452 23354 10464
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 23348 10424 23397 10452
rect 23348 10412 23354 10424
rect 23385 10421 23397 10424
rect 23431 10421 23443 10455
rect 23385 10415 23443 10421
rect 1104 10362 27876 10384
rect 1104 10310 4296 10362
rect 4348 10310 4360 10362
rect 4412 10310 4424 10362
rect 4476 10310 4488 10362
rect 4540 10310 4552 10362
rect 4604 10310 10988 10362
rect 11040 10310 11052 10362
rect 11104 10310 11116 10362
rect 11168 10310 11180 10362
rect 11232 10310 11244 10362
rect 11296 10310 17680 10362
rect 17732 10310 17744 10362
rect 17796 10310 17808 10362
rect 17860 10310 17872 10362
rect 17924 10310 17936 10362
rect 17988 10310 24372 10362
rect 24424 10310 24436 10362
rect 24488 10310 24500 10362
rect 24552 10310 24564 10362
rect 24616 10310 24628 10362
rect 24680 10310 27876 10362
rect 1104 10288 27876 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 7377 10251 7435 10257
rect 7377 10248 7389 10251
rect 5592 10220 7389 10248
rect 5592 10208 5598 10220
rect 7377 10217 7389 10220
rect 7423 10217 7435 10251
rect 7377 10211 7435 10217
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 9122 10248 9128 10260
rect 7883 10220 9128 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12860 10220 12909 10248
rect 12860 10208 12866 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 13722 10248 13728 10260
rect 13683 10220 13728 10248
rect 12897 10211 12955 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 18322 10248 18328 10260
rect 15151 10220 18328 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 19429 10251 19487 10257
rect 19429 10217 19441 10251
rect 19475 10248 19487 10251
rect 19518 10248 19524 10260
rect 19475 10220 19524 10248
rect 19475 10217 19487 10220
rect 19429 10211 19487 10217
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 20254 10208 20260 10260
rect 20312 10248 20318 10260
rect 22557 10251 22615 10257
rect 22557 10248 22569 10251
rect 20312 10220 22569 10248
rect 20312 10208 20318 10220
rect 22557 10217 22569 10220
rect 22603 10217 22615 10251
rect 24762 10248 24768 10260
rect 24723 10220 24768 10248
rect 22557 10211 22615 10217
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 8573 10183 8631 10189
rect 8573 10149 8585 10183
rect 8619 10180 8631 10183
rect 11514 10180 11520 10192
rect 8619 10152 11520 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 13630 10180 13636 10192
rect 11992 10152 13636 10180
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 4706 10112 4712 10124
rect 2915 10084 4712 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5445 10115 5503 10121
rect 5445 10081 5457 10115
rect 5491 10112 5503 10115
rect 5534 10112 5540 10124
rect 5491 10084 5540 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 7466 10112 7472 10124
rect 7427 10084 7472 10112
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 11992 10121 12020 10152
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 22094 10180 22100 10192
rect 22055 10152 22100 10180
rect 22094 10140 22100 10152
rect 22152 10140 22158 10192
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10081 12035 10115
rect 11977 10075 12035 10081
rect 12253 10115 12311 10121
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12299 10084 13001 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 14826 10112 14832 10124
rect 14787 10084 14832 10112
rect 12989 10075 13047 10081
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15344 10084 15761 10112
rect 15344 10072 15350 10084
rect 15749 10081 15761 10084
rect 15795 10112 15807 10115
rect 17310 10112 17316 10124
rect 15795 10084 17316 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18506 10072 18512 10124
rect 18564 10112 18570 10124
rect 19981 10115 20039 10121
rect 19981 10112 19993 10115
rect 18564 10084 19993 10112
rect 18564 10072 18570 10084
rect 19981 10081 19993 10084
rect 20027 10081 20039 10115
rect 23106 10112 23112 10124
rect 23067 10084 23112 10112
rect 19981 10075 20039 10081
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2685 10047 2743 10053
rect 2685 10044 2697 10047
rect 2188 10016 2697 10044
rect 2188 10004 2194 10016
rect 2685 10013 2697 10016
rect 2731 10013 2743 10047
rect 2958 10044 2964 10056
rect 2919 10016 2964 10044
rect 2685 10007 2743 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 4522 10044 4528 10056
rect 4483 10016 4528 10044
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10013 9643 10047
rect 9858 10044 9864 10056
rect 9819 10016 9864 10044
rect 9585 10007 9643 10013
rect 1949 9979 2007 9985
rect 1949 9945 1961 9979
rect 1995 9976 2007 9979
rect 7374 9976 7380 9988
rect 1995 9948 3004 9976
rect 7335 9948 7380 9976
rect 1995 9945 2007 9948
rect 1949 9939 2007 9945
rect 2976 9920 3004 9948
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 8386 9976 8392 9988
rect 8347 9948 8392 9976
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 9600 9976 9628 10007
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10778 10044 10784 10056
rect 10739 10016 10784 10044
rect 10778 10004 10784 10016
rect 10836 10044 10842 10056
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 10836 10016 11897 10044
rect 10836 10004 10842 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10044 12955 10047
rect 13078 10044 13084 10056
rect 12943 10016 13084 10044
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 15378 10044 15384 10056
rect 14783 10016 15384 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 16758 10044 16764 10056
rect 16719 10016 16764 10044
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17494 10044 17500 10056
rect 17451 10016 17500 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 19794 10044 19800 10056
rect 19576 10016 19800 10044
rect 19576 10004 19582 10016
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 20990 10053 20996 10056
rect 20717 10047 20775 10053
rect 20717 10013 20729 10047
rect 20763 10013 20775 10047
rect 20984 10044 20996 10053
rect 20951 10016 20996 10044
rect 20717 10007 20775 10013
rect 20984 10007 20996 10016
rect 10686 9976 10692 9988
rect 8536 9948 10364 9976
rect 10647 9948 10692 9976
rect 8536 9936 8542 9948
rect 2498 9908 2504 9920
rect 2459 9880 2504 9908
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 2958 9868 2964 9920
rect 3016 9868 3022 9920
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 4154 9908 4160 9920
rect 4019 9880 4160 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 10226 9908 10232 9920
rect 6972 9880 7017 9908
rect 10187 9880 10232 9908
rect 6972 9868 6978 9880
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10336 9908 10364 9948
rect 10686 9936 10692 9948
rect 10744 9936 10750 9988
rect 13173 9979 13231 9985
rect 10796 9948 12434 9976
rect 10796 9908 10824 9948
rect 10336 9880 10824 9908
rect 12406 9908 12434 9948
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 14182 9976 14188 9988
rect 13219 9948 14188 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 14826 9936 14832 9988
rect 14884 9976 14890 9988
rect 15933 9979 15991 9985
rect 15933 9976 15945 9979
rect 14884 9948 15945 9976
rect 14884 9936 14890 9948
rect 15933 9945 15945 9948
rect 15979 9976 15991 9979
rect 16574 9976 16580 9988
rect 15979 9948 16580 9976
rect 15979 9945 15991 9948
rect 15933 9939 15991 9945
rect 16574 9936 16580 9948
rect 16632 9936 16638 9988
rect 17650 9979 17708 9985
rect 17650 9976 17662 9979
rect 16960 9948 17662 9976
rect 13262 9908 13268 9920
rect 12406 9880 13268 9908
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 15838 9908 15844 9920
rect 15799 9880 15844 9908
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 16960 9917 16988 9948
rect 17650 9945 17662 9948
rect 17696 9945 17708 9979
rect 17650 9939 17708 9945
rect 19242 9936 19248 9988
rect 19300 9976 19306 9988
rect 20732 9976 20760 10007
rect 20990 10004 20996 10007
rect 21048 10004 21054 10056
rect 23750 10044 23756 10056
rect 23711 10016 23756 10044
rect 23750 10004 23756 10016
rect 23808 10044 23814 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 23808 10016 24593 10044
rect 23808 10004 23814 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 20806 9976 20812 9988
rect 19300 9948 20812 9976
rect 19300 9936 19306 9948
rect 20806 9936 20812 9948
rect 20864 9976 20870 9988
rect 22002 9976 22008 9988
rect 20864 9948 22008 9976
rect 20864 9936 20870 9948
rect 22002 9936 22008 9948
rect 22060 9936 22066 9988
rect 23382 9976 23388 9988
rect 22940 9948 23388 9976
rect 22940 9920 22968 9948
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 24029 9979 24087 9985
rect 24029 9945 24041 9979
rect 24075 9976 24087 9979
rect 25222 9976 25228 9988
rect 24075 9948 25228 9976
rect 24075 9945 24087 9948
rect 24029 9939 24087 9945
rect 25222 9936 25228 9948
rect 25280 9936 25286 9988
rect 16301 9911 16359 9917
rect 16301 9908 16313 9911
rect 16172 9880 16313 9908
rect 16172 9868 16178 9880
rect 16301 9877 16313 9880
rect 16347 9877 16359 9911
rect 16301 9871 16359 9877
rect 16945 9911 17003 9917
rect 16945 9877 16957 9911
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18472 9880 18797 9908
rect 18472 9868 18478 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18785 9871 18843 9877
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20530 9908 20536 9920
rect 19935 9880 20536 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 22922 9908 22928 9920
rect 22883 9880 22928 9908
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 23017 9911 23075 9917
rect 23017 9877 23029 9911
rect 23063 9908 23075 9911
rect 23290 9908 23296 9920
rect 23063 9880 23296 9908
rect 23063 9877 23075 9880
rect 23017 9871 23075 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 23400 9908 23428 9936
rect 25317 9911 25375 9917
rect 25317 9908 25329 9911
rect 23400 9880 25329 9908
rect 25317 9877 25329 9880
rect 25363 9877 25375 9911
rect 25317 9871 25375 9877
rect 1104 9818 28032 9840
rect 1104 9766 7642 9818
rect 7694 9766 7706 9818
rect 7758 9766 7770 9818
rect 7822 9766 7834 9818
rect 7886 9766 7898 9818
rect 7950 9766 14334 9818
rect 14386 9766 14398 9818
rect 14450 9766 14462 9818
rect 14514 9766 14526 9818
rect 14578 9766 14590 9818
rect 14642 9766 21026 9818
rect 21078 9766 21090 9818
rect 21142 9766 21154 9818
rect 21206 9766 21218 9818
rect 21270 9766 21282 9818
rect 21334 9766 27718 9818
rect 27770 9766 27782 9818
rect 27834 9766 27846 9818
rect 27898 9766 27910 9818
rect 27962 9766 27974 9818
rect 28026 9766 28032 9818
rect 1104 9744 28032 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 10042 9704 10048 9716
rect 4580 9676 10048 9704
rect 4580 9664 4586 9676
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 10134 9664 10140 9716
rect 10192 9704 10198 9716
rect 11422 9704 11428 9716
rect 10192 9676 11428 9704
rect 10192 9664 10198 9676
rect 11422 9664 11428 9676
rect 11480 9704 11486 9716
rect 12710 9704 12716 9716
rect 11480 9676 12716 9704
rect 11480 9664 11486 9676
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 16298 9704 16304 9716
rect 15896 9676 16304 9704
rect 15896 9664 15902 9676
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 20530 9704 20536 9716
rect 20491 9676 20536 9704
rect 20530 9664 20536 9676
rect 20588 9664 20594 9716
rect 2308 9639 2366 9645
rect 2308 9605 2320 9639
rect 2354 9636 2366 9639
rect 2498 9636 2504 9648
rect 2354 9608 2504 9636
rect 2354 9605 2366 9608
rect 2308 9599 2366 9605
rect 2498 9596 2504 9608
rect 2556 9596 2562 9648
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3936 9608 3985 9636
rect 3936 9596 3942 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 4154 9636 4160 9648
rect 4115 9608 4160 9636
rect 3973 9599 4031 9605
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 3988 9568 4016 9599
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 6546 9636 6552 9648
rect 5092 9608 5396 9636
rect 6507 9608 6552 9636
rect 5092 9568 5120 9608
rect 5258 9568 5264 9580
rect 3988 9540 5120 9568
rect 5219 9540 5264 9568
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5368 9568 5396 9608
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 8386 9636 8392 9648
rect 6886 9608 8392 9636
rect 6886 9568 6914 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 12805 9639 12863 9645
rect 12805 9605 12817 9639
rect 12851 9636 12863 9639
rect 13814 9636 13820 9648
rect 12851 9608 13820 9636
rect 12851 9605 12863 9608
rect 12805 9599 12863 9605
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9636 14519 9639
rect 15470 9636 15476 9648
rect 14507 9608 15476 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 15470 9596 15476 9608
rect 15528 9596 15534 9648
rect 17494 9596 17500 9648
rect 17552 9636 17558 9648
rect 23014 9636 23020 9648
rect 17552 9608 18455 9636
rect 17552 9596 17558 9608
rect 7006 9568 7012 9580
rect 5368 9540 6914 9568
rect 6967 9540 7012 9568
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7248 9540 7389 9568
rect 7248 9528 7254 9540
rect 7377 9537 7389 9540
rect 7423 9568 7435 9571
rect 8297 9571 8355 9577
rect 7423 9540 8248 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 4672 9472 5181 9500
rect 4672 9460 4678 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 4522 9432 4528 9444
rect 3620 9404 4528 9432
rect 3620 9376 3648 9404
rect 4522 9392 4528 9404
rect 4580 9392 4586 9444
rect 5629 9435 5687 9441
rect 5629 9401 5641 9435
rect 5675 9432 5687 9435
rect 7466 9432 7472 9444
rect 5675 9404 7472 9432
rect 5675 9401 5687 9404
rect 5629 9395 5687 9401
rect 7466 9392 7472 9404
rect 7524 9392 7530 9444
rect 8220 9432 8248 9540
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8754 9568 8760 9580
rect 8343 9540 8760 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 12713 9571 12771 9577
rect 11747 9540 12388 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8435 9472 8861 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 10686 9500 10692 9512
rect 9171 9472 10692 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 8478 9432 8484 9444
rect 8220 9404 8484 9432
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 12360 9441 12388 9540
rect 12713 9537 12725 9571
rect 12759 9568 12771 9571
rect 13722 9568 13728 9580
rect 12759 9540 13584 9568
rect 13683 9540 13728 9568
rect 12759 9537 12771 9540
rect 12713 9531 12771 9537
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9469 12955 9503
rect 13556 9500 13584 9540
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15010 9568 15016 9580
rect 14967 9540 15016 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 15188 9571 15246 9577
rect 15188 9537 15200 9571
rect 15234 9568 15246 9571
rect 15930 9568 15936 9580
rect 15234 9540 15936 9568
rect 15234 9537 15246 9540
rect 15188 9531 15246 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 17144 9540 17233 9568
rect 14826 9500 14832 9512
rect 13556 9472 14832 9500
rect 12897 9463 12955 9469
rect 12345 9435 12403 9441
rect 12345 9401 12357 9435
rect 12391 9401 12403 9435
rect 12345 9395 12403 9401
rect 12710 9392 12716 9444
rect 12768 9432 12774 9444
rect 12912 9432 12940 9463
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 12768 9404 12940 9432
rect 15856 9404 16865 9432
rect 12768 9392 12774 9404
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 3602 9364 3608 9376
rect 3467 9336 3608 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10192 9336 10609 9364
rect 10192 9324 10198 9336
rect 10597 9333 10609 9336
rect 10643 9364 10655 9367
rect 10778 9364 10784 9376
rect 10643 9336 10784 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 13538 9364 13544 9376
rect 13499 9336 13544 9364
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 15856 9364 15884 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 17144 9432 17172 9540
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17586 9528 17592 9580
rect 17644 9568 17650 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17644 9540 18245 9568
rect 17644 9528 17650 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 17310 9500 17316 9512
rect 17271 9472 17316 9500
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 18322 9500 18328 9512
rect 17460 9472 17505 9500
rect 18283 9472 18328 9500
rect 17460 9460 17466 9472
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 18427 9500 18455 9608
rect 18524 9608 23020 9636
rect 18524 9577 18552 9608
rect 23014 9596 23020 9608
rect 23072 9596 23078 9648
rect 24762 9596 24768 9648
rect 24820 9596 24826 9648
rect 25222 9636 25228 9648
rect 25183 9608 25228 9636
rect 25222 9596 25228 9608
rect 25280 9596 25286 9648
rect 18509 9571 18567 9577
rect 18509 9537 18521 9571
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 19242 9528 19248 9580
rect 19300 9528 19306 9580
rect 19426 9577 19432 9580
rect 19420 9568 19432 9577
rect 19387 9540 19432 9568
rect 19420 9531 19432 9540
rect 19426 9528 19432 9531
rect 19484 9528 19490 9580
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 19852 9540 21189 9568
rect 19852 9528 19858 9540
rect 21177 9537 21189 9540
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 22373 9571 22431 9577
rect 22373 9537 22385 9571
rect 22419 9568 22431 9571
rect 22646 9568 22652 9580
rect 22419 9540 22652 9568
rect 22419 9537 22431 9540
rect 22373 9531 22431 9537
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 23198 9568 23204 9580
rect 23159 9540 23204 9568
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18427 9472 19165 9500
rect 19153 9469 19165 9472
rect 19199 9500 19211 9503
rect 19260 9500 19288 9528
rect 19199 9472 19288 9500
rect 19199 9469 19211 9472
rect 19153 9463 19211 9469
rect 20530 9460 20536 9512
rect 20588 9500 20594 9512
rect 22281 9503 22339 9509
rect 22281 9500 22293 9503
rect 20588 9472 22293 9500
rect 20588 9460 20594 9472
rect 22281 9469 22293 9472
rect 22327 9469 22339 9503
rect 25498 9500 25504 9512
rect 25459 9472 25504 9500
rect 22281 9463 22339 9469
rect 25498 9460 25504 9472
rect 25556 9460 25562 9512
rect 18046 9432 18052 9444
rect 17144 9404 18052 9432
rect 16853 9395 16911 9401
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 22830 9432 22836 9444
rect 18524 9404 19012 9432
rect 18524 9373 18552 9404
rect 14608 9336 15884 9364
rect 18509 9367 18567 9373
rect 14608 9324 14614 9336
rect 18509 9333 18521 9367
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 18693 9367 18751 9373
rect 18693 9333 18705 9367
rect 18739 9364 18751 9367
rect 18874 9364 18880 9376
rect 18739 9336 18880 9364
rect 18739 9333 18751 9336
rect 18693 9327 18751 9333
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 18984 9364 19012 9404
rect 20180 9404 22836 9432
rect 20180 9364 20208 9404
rect 22830 9392 22836 9404
rect 22888 9392 22894 9444
rect 18984 9336 20208 9364
rect 20714 9324 20720 9376
rect 20772 9364 20778 9376
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 20772 9336 21005 9364
rect 20772 9324 20778 9336
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 20993 9327 21051 9333
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21140 9336 22017 9364
rect 21140 9324 21146 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 23293 9367 23351 9373
rect 23293 9333 23305 9367
rect 23339 9364 23351 9367
rect 23566 9364 23572 9376
rect 23339 9336 23572 9364
rect 23339 9333 23351 9336
rect 23293 9327 23351 9333
rect 23566 9324 23572 9336
rect 23624 9324 23630 9376
rect 23750 9364 23756 9376
rect 23711 9336 23756 9364
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 1104 9274 27876 9296
rect 1104 9222 4296 9274
rect 4348 9222 4360 9274
rect 4412 9222 4424 9274
rect 4476 9222 4488 9274
rect 4540 9222 4552 9274
rect 4604 9222 10988 9274
rect 11040 9222 11052 9274
rect 11104 9222 11116 9274
rect 11168 9222 11180 9274
rect 11232 9222 11244 9274
rect 11296 9222 17680 9274
rect 17732 9222 17744 9274
rect 17796 9222 17808 9274
rect 17860 9222 17872 9274
rect 17924 9222 17936 9274
rect 17988 9222 24372 9274
rect 24424 9222 24436 9274
rect 24488 9222 24500 9274
rect 24552 9222 24564 9274
rect 24616 9222 24628 9274
rect 24680 9222 27876 9274
rect 1104 9200 27876 9222
rect 2038 9160 2044 9172
rect 1872 9132 2044 9160
rect 1872 9033 1900 9132
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 5077 9163 5135 9169
rect 5077 9129 5089 9163
rect 5123 9160 5135 9163
rect 5166 9160 5172 9172
rect 5123 9132 5172 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 7282 9160 7288 9172
rect 5276 9132 7288 9160
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9061 3295 9095
rect 4982 9092 4988 9104
rect 3237 9055 3295 9061
rect 4172 9064 4988 9092
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 8993 1915 9027
rect 1857 8987 1915 8993
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 3252 9024 3280 9055
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 3200 8996 3985 9024
rect 3200 8984 3206 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 4172 8968 4200 9064
rect 4982 9052 4988 9064
rect 5040 9092 5046 9104
rect 5276 9092 5304 9132
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7432 9132 8033 9160
rect 7432 9120 7438 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 8021 9123 8079 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9766 9160 9772 9172
rect 9171 9132 9772 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 5040 9064 5304 9092
rect 5040 9052 5046 9064
rect 8481 9027 8539 9033
rect 5092 8996 8340 9024
rect 4154 8956 4160 8968
rect 4067 8928 4160 8956
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 5092 8965 5120 8996
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5077 8919 5135 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 2124 8891 2182 8897
rect 2124 8857 2136 8891
rect 2170 8888 2182 8891
rect 2682 8888 2688 8900
rect 2170 8860 2688 8888
rect 2170 8857 2182 8860
rect 2124 8851 2182 8857
rect 2682 8848 2688 8860
rect 2740 8848 2746 8900
rect 5810 8888 5816 8900
rect 5771 8860 5816 8888
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 6546 8848 6552 8900
rect 6604 8848 6610 8900
rect 8312 8888 8340 8996
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 9140 9024 9168 9123
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11609 9163 11667 9169
rect 11609 9129 11621 9163
rect 11655 9160 11667 9163
rect 12802 9160 12808 9172
rect 11655 9132 12808 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 16577 9163 16635 9169
rect 13320 9132 16528 9160
rect 13320 9120 13326 9132
rect 16500 9092 16528 9132
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 16942 9160 16948 9172
rect 16623 9132 16948 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 16942 9120 16948 9132
rect 17000 9160 17006 9172
rect 17310 9160 17316 9172
rect 17000 9132 17316 9160
rect 17000 9120 17006 9132
rect 17310 9120 17316 9132
rect 17368 9120 17374 9172
rect 17586 9160 17592 9172
rect 17547 9132 17592 9160
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18417 9163 18475 9169
rect 18417 9160 18429 9163
rect 18196 9132 18429 9160
rect 18196 9120 18202 9132
rect 18417 9129 18429 9132
rect 18463 9129 18475 9163
rect 18417 9123 18475 9129
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 21082 9160 21088 9172
rect 18923 9132 21088 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 22830 9160 22836 9172
rect 22791 9132 22836 9160
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 23845 9095 23903 9101
rect 23845 9092 23857 9095
rect 16500 9064 19012 9092
rect 8527 8996 9168 9024
rect 11333 9027 11391 9033
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 11333 8993 11345 9027
rect 11379 9024 11391 9027
rect 11790 9024 11796 9036
rect 11379 8996 11796 9024
rect 11379 8993 11391 8996
rect 11333 8987 11391 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 15194 9024 15200 9036
rect 11940 8996 12204 9024
rect 15155 8996 15200 9024
rect 11940 8984 11946 8996
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8754 8956 8760 8968
rect 8435 8928 8760 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 11241 8959 11299 8965
rect 10551 8928 11100 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10134 8888 10140 8900
rect 8312 8860 10140 8888
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 10260 8891 10318 8897
rect 10260 8857 10272 8891
rect 10306 8888 10318 8891
rect 10962 8888 10968 8900
rect 10306 8860 10968 8888
rect 10306 8857 10318 8860
rect 10260 8851 10318 8857
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11072 8888 11100 8928
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11422 8956 11428 8968
rect 11287 8928 11428 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 12066 8956 12072 8968
rect 12027 8928 12072 8956
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12176 8956 12204 8996
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 16356 8996 17141 9024
rect 16356 8984 16362 8996
rect 17129 8993 17141 8996
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 12325 8959 12383 8965
rect 12325 8956 12337 8959
rect 12176 8928 12337 8956
rect 12325 8925 12337 8928
rect 12371 8925 12383 8959
rect 14550 8956 14556 8968
rect 14511 8928 14556 8956
rect 12325 8919 12383 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 17218 8956 17224 8968
rect 17179 8928 17224 8956
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 18598 8956 18604 8968
rect 18559 8928 18604 8956
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 18874 8956 18880 8968
rect 18748 8928 18793 8956
rect 18835 8928 18880 8956
rect 18748 8916 18754 8928
rect 18874 8916 18880 8928
rect 18932 8916 18938 8968
rect 18984 8956 19012 9064
rect 21560 9064 23857 9092
rect 20806 9024 20812 9036
rect 20767 8996 20812 9024
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 20553 8959 20611 8965
rect 18984 8928 20484 8956
rect 11514 8888 11520 8900
rect 11072 8860 11520 8888
rect 11514 8848 11520 8860
rect 11572 8888 11578 8900
rect 12084 8888 12112 8916
rect 15442 8891 15500 8897
rect 15442 8888 15454 8891
rect 11572 8860 12112 8888
rect 14752 8860 15454 8888
rect 11572 8848 11578 8860
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 4614 8820 4620 8832
rect 4387 8792 4620 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 4614 8780 4620 8792
rect 4672 8780 4678 8832
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 6880 8792 7297 8820
rect 6880 8780 6886 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 13449 8823 13507 8829
rect 13449 8789 13461 8823
rect 13495 8820 13507 8823
rect 13814 8820 13820 8832
rect 13495 8792 13820 8820
rect 13495 8789 13507 8792
rect 13449 8783 13507 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14752 8829 14780 8860
rect 15442 8857 15454 8860
rect 15488 8857 15500 8891
rect 15442 8851 15500 8857
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8789 14795 8823
rect 19426 8820 19432 8832
rect 19387 8792 19432 8820
rect 14737 8783 14795 8789
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 20456 8820 20484 8928
rect 20553 8925 20565 8959
rect 20599 8956 20611 8959
rect 20714 8956 20720 8968
rect 20599 8928 20720 8956
rect 20599 8925 20611 8928
rect 20553 8919 20611 8925
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 21560 8965 21588 9064
rect 23845 9061 23857 9064
rect 23891 9092 23903 9095
rect 24946 9092 24952 9104
rect 23891 9064 24952 9092
rect 23891 9061 23903 9064
rect 23845 9055 23903 9061
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 23109 9027 23167 9033
rect 23109 9024 23121 9027
rect 22152 8996 23121 9024
rect 22152 8984 22158 8996
rect 23109 8993 23121 8996
rect 23155 8993 23167 9027
rect 23109 8987 23167 8993
rect 24673 9027 24731 9033
rect 24673 8993 24685 9027
rect 24719 9024 24731 9027
rect 24762 9024 24768 9036
rect 24719 8996 24768 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 24762 8984 24768 8996
rect 24820 8984 24826 9036
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 20916 8928 21557 8956
rect 20916 8820 20944 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 22002 8956 22008 8968
rect 21915 8928 22008 8956
rect 21545 8919 21603 8925
rect 22002 8916 22008 8928
rect 22060 8956 22066 8968
rect 23198 8956 23204 8968
rect 22060 8928 22140 8956
rect 23159 8928 23204 8956
rect 22060 8916 22066 8928
rect 22112 8888 22140 8928
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 25130 8956 25136 8968
rect 25091 8928 25136 8956
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 25314 8956 25320 8968
rect 25275 8928 25320 8956
rect 25314 8916 25320 8928
rect 25372 8956 25378 8968
rect 26142 8956 26148 8968
rect 25372 8928 26148 8956
rect 25372 8916 25378 8928
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 25148 8888 25176 8916
rect 22112 8860 25176 8888
rect 20456 8792 20944 8820
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 22373 8823 22431 8829
rect 22373 8820 22385 8823
rect 22336 8792 22385 8820
rect 22336 8780 22342 8792
rect 22373 8789 22385 8792
rect 22419 8789 22431 8823
rect 22373 8783 22431 8789
rect 1104 8730 28032 8752
rect 1104 8678 7642 8730
rect 7694 8678 7706 8730
rect 7758 8678 7770 8730
rect 7822 8678 7834 8730
rect 7886 8678 7898 8730
rect 7950 8678 14334 8730
rect 14386 8678 14398 8730
rect 14450 8678 14462 8730
rect 14514 8678 14526 8730
rect 14578 8678 14590 8730
rect 14642 8678 21026 8730
rect 21078 8678 21090 8730
rect 21142 8678 21154 8730
rect 21206 8678 21218 8730
rect 21270 8678 21282 8730
rect 21334 8678 27718 8730
rect 27770 8678 27782 8730
rect 27834 8678 27846 8730
rect 27898 8678 27910 8730
rect 27962 8678 27974 8730
rect 28026 8678 28032 8730
rect 1104 8656 28032 8678
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 3697 8619 3755 8625
rect 3697 8616 3709 8619
rect 2832 8588 3709 8616
rect 2832 8576 2838 8588
rect 3697 8585 3709 8588
rect 3743 8616 3755 8619
rect 4062 8616 4068 8628
rect 3743 8588 4068 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 5592 8588 5641 8616
rect 5592 8576 5598 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 6546 8616 6552 8628
rect 6507 8588 6552 8616
rect 5629 8579 5687 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 10962 8616 10968 8628
rect 10923 8588 10968 8616
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 12529 8619 12587 8625
rect 12529 8585 12541 8619
rect 12575 8616 12587 8619
rect 13170 8616 13176 8628
rect 12575 8588 13176 8616
rect 12575 8585 12587 8588
rect 12529 8579 12587 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 15930 8616 15936 8628
rect 15891 8588 15936 8616
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 19245 8619 19303 8625
rect 16632 8588 16988 8616
rect 16632 8576 16638 8588
rect 1949 8551 2007 8557
rect 1949 8517 1961 8551
rect 1995 8548 2007 8551
rect 2314 8548 2320 8560
rect 1995 8520 2320 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 4614 8548 4620 8560
rect 2792 8520 4620 8548
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2792 8480 2820 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5718 8548 5724 8560
rect 5092 8520 5724 8548
rect 2271 8452 2820 8480
rect 2869 8483 2927 8489
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 3142 8480 3148 8492
rect 3103 8452 3148 8480
rect 2869 8443 2927 8449
rect 2148 8412 2176 8443
rect 2774 8412 2780 8424
rect 2148 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2884 8412 2912 8443
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3878 8480 3884 8492
rect 3839 8452 3884 8480
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 5092 8489 5120 8520
rect 5718 8508 5724 8520
rect 5776 8548 5782 8560
rect 6454 8548 6460 8560
rect 5776 8520 6460 8548
rect 5776 8508 5782 8520
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 6880 8520 8340 8548
rect 6880 8508 6886 8520
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6914 8480 6920 8492
rect 5859 8452 6920 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7190 8480 7196 8492
rect 7064 8452 7109 8480
rect 7151 8452 7196 8480
rect 7064 8440 7070 8452
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 8312 8489 8340 8520
rect 9214 8508 9220 8560
rect 9272 8508 9278 8560
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12952 8520 13001 8548
rect 12952 8508 12958 8520
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 12989 8511 13047 8517
rect 14737 8551 14795 8557
rect 14737 8517 14749 8551
rect 14783 8548 14795 8551
rect 16850 8548 16856 8560
rect 14783 8520 16856 8548
rect 14783 8517 14795 8520
rect 14737 8511 14795 8517
rect 16850 8508 16856 8520
rect 16908 8508 16914 8560
rect 16960 8557 16988 8588
rect 19245 8585 19257 8619
rect 19291 8616 19303 8619
rect 19794 8616 19800 8628
rect 19291 8588 19800 8616
rect 19291 8585 19303 8588
rect 19245 8579 19303 8585
rect 19794 8576 19800 8588
rect 19852 8576 19858 8628
rect 23198 8576 23204 8628
rect 23256 8616 23262 8628
rect 25041 8619 25099 8625
rect 25041 8616 25053 8619
rect 23256 8588 25053 8616
rect 23256 8576 23262 8588
rect 25041 8585 25053 8588
rect 25087 8585 25099 8619
rect 25041 8579 25099 8585
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8548 17003 8551
rect 19518 8548 19524 8560
rect 16991 8520 19524 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 19518 8508 19524 8520
rect 19576 8508 19582 8560
rect 19702 8548 19708 8560
rect 19663 8520 19708 8548
rect 19702 8508 19708 8520
rect 19760 8508 19766 8560
rect 22922 8548 22928 8560
rect 19812 8520 22928 8548
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7340 8452 8125 8480
rect 7340 8440 7346 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8480 11207 8483
rect 11330 8480 11336 8492
rect 11195 8452 11336 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 13446 8480 13452 8492
rect 12023 8452 13452 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 15378 8480 15384 8492
rect 15339 8452 15384 8480
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18506 8480 18512 8492
rect 18095 8452 18512 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 4706 8412 4712 8424
rect 2884 8384 4712 8412
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 5902 8412 5908 8424
rect 5092 8384 5908 8412
rect 1949 8347 2007 8353
rect 1949 8313 1961 8347
rect 1995 8344 2007 8347
rect 2130 8344 2136 8356
rect 1995 8316 2136 8344
rect 1995 8313 2007 8316
rect 1949 8307 2007 8313
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 4154 8344 4160 8356
rect 3099 8316 4160 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 5092 8353 5120 8384
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11664 8384 11713 8412
rect 11664 8372 11670 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 17880 8412 17908 8443
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18966 8480 18972 8492
rect 18923 8452 18972 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18966 8440 18972 8452
rect 19024 8480 19030 8492
rect 19812 8480 19840 8520
rect 22922 8508 22928 8520
rect 22980 8508 22986 8560
rect 23566 8548 23572 8560
rect 23527 8520 23572 8548
rect 23566 8508 23572 8520
rect 23624 8508 23630 8560
rect 19024 8452 19840 8480
rect 19024 8440 19030 8452
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 22373 8483 22431 8489
rect 22373 8480 22385 8483
rect 21416 8452 22385 8480
rect 21416 8440 21422 8452
rect 22373 8449 22385 8452
rect 22419 8449 22431 8483
rect 25056 8480 25084 8579
rect 25498 8576 25504 8628
rect 25556 8616 25562 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 25556 8588 25697 8616
rect 25556 8576 25562 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 25501 8483 25559 8489
rect 25501 8480 25513 8483
rect 22373 8443 22431 8449
rect 18322 8412 18328 8424
rect 17880 8384 18328 8412
rect 11701 8375 11759 8381
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 18414 8372 18420 8424
rect 18472 8412 18478 8424
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 18472 8384 18613 8412
rect 18472 8372 18478 8384
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8412 18843 8415
rect 19426 8412 19432 8424
rect 18831 8384 19432 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 19426 8372 19432 8384
rect 19484 8412 19490 8424
rect 22281 8415 22339 8421
rect 22281 8412 22293 8415
rect 19484 8384 22293 8412
rect 19484 8372 19490 8384
rect 22281 8381 22293 8384
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23934 8412 23940 8424
rect 23339 8384 23940 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23934 8372 23940 8384
rect 23992 8372 23998 8424
rect 24688 8412 24716 8466
rect 25056 8452 25513 8480
rect 25501 8449 25513 8452
rect 25547 8449 25559 8483
rect 25501 8443 25559 8449
rect 24762 8412 24768 8424
rect 24688 8384 24768 8412
rect 24762 8372 24768 8384
rect 24820 8372 24826 8424
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8313 5135 8347
rect 5077 8307 5135 8313
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 8113 8347 8171 8353
rect 8113 8344 8125 8347
rect 5684 8316 8125 8344
rect 5684 8304 5690 8316
rect 8113 8313 8125 8316
rect 8159 8313 8171 8347
rect 8754 8344 8760 8356
rect 8715 8316 8760 8344
rect 8113 8307 8171 8313
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 18690 8304 18696 8356
rect 18748 8344 18754 8356
rect 22005 8347 22063 8353
rect 22005 8344 22017 8347
rect 18748 8316 22017 8344
rect 18748 8304 18754 8316
rect 22005 8313 22017 8316
rect 22051 8313 22063 8347
rect 22005 8307 22063 8313
rect 15286 8276 15292 8288
rect 15247 8248 15292 8276
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 17957 8279 18015 8285
rect 17957 8245 17969 8279
rect 18003 8276 18015 8279
rect 18230 8276 18236 8288
rect 18003 8248 18236 8276
rect 18003 8245 18015 8248
rect 17957 8239 18015 8245
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 20806 8236 20812 8288
rect 20864 8276 20870 8288
rect 20993 8279 21051 8285
rect 20993 8276 21005 8279
rect 20864 8248 21005 8276
rect 20864 8236 20870 8248
rect 20993 8245 21005 8248
rect 21039 8245 21051 8279
rect 20993 8239 21051 8245
rect 1104 8186 27876 8208
rect 1104 8134 4296 8186
rect 4348 8134 4360 8186
rect 4412 8134 4424 8186
rect 4476 8134 4488 8186
rect 4540 8134 4552 8186
rect 4604 8134 10988 8186
rect 11040 8134 11052 8186
rect 11104 8134 11116 8186
rect 11168 8134 11180 8186
rect 11232 8134 11244 8186
rect 11296 8134 17680 8186
rect 17732 8134 17744 8186
rect 17796 8134 17808 8186
rect 17860 8134 17872 8186
rect 17924 8134 17936 8186
rect 17988 8134 24372 8186
rect 24424 8134 24436 8186
rect 24488 8134 24500 8186
rect 24552 8134 24564 8186
rect 24616 8134 24628 8186
rect 24680 8134 27876 8186
rect 1104 8112 27876 8134
rect 2038 8072 2044 8084
rect 1999 8044 2044 8072
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5868 8044 6009 8072
rect 5868 8032 5874 8044
rect 5997 8041 6009 8044
rect 6043 8041 6055 8075
rect 5997 8035 6055 8041
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7374 8072 7380 8084
rect 7248 8044 7380 8072
rect 7248 8032 7254 8044
rect 7374 8032 7380 8044
rect 7432 8072 7438 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7432 8044 8033 8072
rect 7432 8032 7438 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8996 8044 9137 8072
rect 8996 8032 9002 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 10226 8072 10232 8084
rect 9907 8044 10232 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13722 8072 13728 8084
rect 13403 8044 13728 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14240 8044 14289 8072
rect 14240 8032 14246 8044
rect 14277 8041 14289 8044
rect 14323 8041 14335 8075
rect 14277 8035 14335 8041
rect 18509 8075 18567 8081
rect 18509 8041 18521 8075
rect 18555 8072 18567 8075
rect 18598 8072 18604 8084
rect 18555 8044 18604 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 19518 8072 19524 8084
rect 19479 8044 19524 8072
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 22097 8075 22155 8081
rect 22097 8072 22109 8075
rect 22060 8044 22109 8072
rect 22060 8032 22066 8044
rect 22097 8041 22109 8044
rect 22143 8041 22155 8075
rect 23014 8072 23020 8084
rect 22975 8044 23020 8072
rect 22097 8035 22155 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 26142 8072 26148 8084
rect 26103 8044 26148 8072
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 6730 7936 6736 7948
rect 6196 7908 6736 7936
rect 6196 7880 6224 7908
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 12158 7936 12164 7948
rect 12119 7908 12164 7936
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12710 7936 12716 7948
rect 12671 7908 12716 7936
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 14553 7939 14611 7945
rect 14553 7936 14565 7939
rect 13872 7908 14565 7936
rect 13872 7896 13878 7908
rect 14553 7905 14565 7908
rect 14599 7905 14611 7939
rect 23290 7936 23296 7948
rect 23251 7908 23296 7936
rect 14553 7899 14611 7905
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 24673 7939 24731 7945
rect 24673 7905 24685 7939
rect 24719 7936 24731 7939
rect 24762 7936 24768 7948
rect 24719 7908 24768 7936
rect 24719 7905 24731 7908
rect 24673 7899 24731 7905
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 2188 7840 3985 7868
rect 2188 7828 2194 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 4120 7840 4169 7868
rect 4120 7828 4126 7840
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 4157 7831 4215 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 6178 7868 6184 7880
rect 6091 7840 6184 7868
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 8812 7840 9689 7868
rect 8812 7828 8818 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10376 7840 10425 7868
rect 10376 7828 10382 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 13964 7840 14657 7868
rect 13964 7828 13970 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 15068 7840 15761 7868
rect 15068 7828 15074 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 16942 7868 16948 7880
rect 16903 7840 16948 7868
rect 15749 7831 15807 7837
rect 3326 7800 3332 7812
rect 3287 7772 3332 7800
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 4341 7803 4399 7809
rect 4341 7769 4353 7803
rect 4387 7800 4399 7803
rect 6733 7803 6791 7809
rect 6733 7800 6745 7803
rect 4387 7772 6745 7800
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 6733 7769 6745 7772
rect 6779 7800 6791 7803
rect 7558 7800 7564 7812
rect 6779 7772 7564 7800
rect 6779 7769 6791 7772
rect 6733 7763 6791 7769
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 12989 7803 13047 7809
rect 12989 7769 13001 7803
rect 13035 7800 13047 7803
rect 15194 7800 15200 7812
rect 13035 7772 15200 7800
rect 13035 7769 13047 7772
rect 12989 7763 13047 7769
rect 15194 7760 15200 7772
rect 15252 7760 15258 7812
rect 15764 7800 15792 7831
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7868 17371 7871
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17359 7840 17969 7868
rect 17359 7837 17371 7840
rect 17313 7831 17371 7837
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 17957 7831 18015 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7868 18383 7871
rect 18414 7868 18420 7880
rect 18371 7840 18420 7868
rect 18371 7837 18383 7840
rect 18325 7831 18383 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 23385 7871 23443 7877
rect 20395 7840 22094 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 17129 7803 17187 7809
rect 17129 7800 17141 7803
rect 15764 7772 17141 7800
rect 17129 7769 17141 7772
rect 17175 7769 17187 7803
rect 18138 7800 18144 7812
rect 18099 7772 18144 7800
rect 17129 7763 17187 7769
rect 18138 7760 18144 7772
rect 18196 7760 18202 7812
rect 20806 7800 20812 7812
rect 20767 7772 20812 7800
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 22066 7800 22094 7840
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 23750 7868 23756 7880
rect 23431 7840 23756 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 23750 7828 23756 7840
rect 23808 7828 23814 7880
rect 25130 7868 25136 7880
rect 25091 7840 25136 7868
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 25222 7828 25228 7880
rect 25280 7868 25286 7880
rect 25409 7871 25467 7877
rect 25409 7868 25421 7871
rect 25280 7840 25421 7868
rect 25280 7828 25286 7840
rect 25409 7837 25421 7840
rect 25455 7868 25467 7871
rect 26142 7868 26148 7880
rect 25455 7840 26148 7868
rect 25455 7837 25467 7840
rect 25409 7831 25467 7837
rect 26142 7828 26148 7840
rect 26200 7828 26206 7880
rect 22646 7800 22652 7812
rect 22066 7772 22652 7800
rect 22646 7760 22652 7772
rect 22704 7760 22710 7812
rect 5350 7732 5356 7744
rect 5311 7704 5356 7732
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 12894 7732 12900 7744
rect 12855 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15749 7735 15807 7741
rect 15749 7732 15761 7735
rect 14884 7704 15761 7732
rect 14884 7692 14890 7704
rect 15749 7701 15761 7704
rect 15795 7701 15807 7735
rect 16482 7732 16488 7744
rect 16395 7704 16488 7732
rect 15749 7695 15807 7701
rect 16482 7692 16488 7704
rect 16540 7732 16546 7744
rect 17954 7732 17960 7744
rect 16540 7704 17960 7732
rect 16540 7692 16546 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 20162 7732 20168 7744
rect 20123 7704 20168 7732
rect 20162 7692 20168 7704
rect 20220 7692 20226 7744
rect 1104 7642 28032 7664
rect 1104 7590 7642 7642
rect 7694 7590 7706 7642
rect 7758 7590 7770 7642
rect 7822 7590 7834 7642
rect 7886 7590 7898 7642
rect 7950 7590 14334 7642
rect 14386 7590 14398 7642
rect 14450 7590 14462 7642
rect 14514 7590 14526 7642
rect 14578 7590 14590 7642
rect 14642 7590 21026 7642
rect 21078 7590 21090 7642
rect 21142 7590 21154 7642
rect 21206 7590 21218 7642
rect 21270 7590 21282 7642
rect 21334 7590 27718 7642
rect 27770 7590 27782 7642
rect 27834 7590 27846 7642
rect 27898 7590 27910 7642
rect 27962 7590 27974 7642
rect 28026 7590 28032 7642
rect 1104 7568 28032 7590
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3384 7500 3893 7528
rect 3384 7488 3390 7500
rect 3881 7497 3893 7500
rect 3927 7497 3939 7531
rect 3881 7491 3939 7497
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 13354 7528 13360 7540
rect 12952 7500 13360 7528
rect 12952 7488 12958 7500
rect 13354 7488 13360 7500
rect 13412 7528 13418 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13412 7500 13553 7528
rect 13412 7488 13418 7500
rect 13541 7497 13553 7500
rect 13587 7497 13599 7531
rect 14090 7528 14096 7540
rect 14051 7500 14096 7528
rect 13541 7491 13599 7497
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 18138 7528 18144 7540
rect 17175 7500 18144 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 18138 7488 18144 7500
rect 18196 7488 18202 7540
rect 18414 7528 18420 7540
rect 18375 7500 18420 7528
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 22554 7488 22560 7540
rect 22612 7528 22618 7540
rect 22649 7531 22707 7537
rect 22649 7528 22661 7531
rect 22612 7500 22661 7528
rect 22612 7488 22618 7500
rect 22649 7497 22661 7500
rect 22695 7497 22707 7531
rect 22649 7491 22707 7497
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 12986 7460 12992 7472
rect 10367 7432 12992 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 12986 7420 12992 7432
rect 13044 7420 13050 7472
rect 14826 7460 14832 7472
rect 14787 7432 14832 7460
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 18322 7420 18328 7472
rect 18380 7460 18386 7472
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 18380 7432 18797 7460
rect 18380 7420 18386 7432
rect 18785 7429 18797 7432
rect 18831 7429 18843 7463
rect 18785 7423 18843 7429
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2130 7392 2136 7404
rect 1903 7364 2136 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 3234 7392 3240 7404
rect 2639 7364 3240 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5626 7392 5632 7404
rect 5123 7364 5632 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 6270 7392 6276 7404
rect 5776 7364 6276 7392
rect 5776 7352 5782 7364
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 7006 7392 7012 7404
rect 6967 7364 7012 7392
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7466 7392 7472 7404
rect 7423 7364 7472 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 12124 7364 12173 7392
rect 12124 7352 12130 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12428 7395 12486 7401
rect 12428 7361 12440 7395
rect 12474 7392 12486 7395
rect 13538 7392 13544 7404
rect 12474 7364 13544 7392
rect 12474 7361 12486 7364
rect 12428 7355 12486 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 15930 7352 15936 7404
rect 15988 7352 15994 7404
rect 16942 7392 16948 7404
rect 16903 7364 16948 7392
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 17129 7355 17187 7361
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4212 7296 4813 7324
rect 4212 7284 4218 7296
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 6546 7324 6552 7336
rect 6507 7296 6552 7324
rect 4801 7287 4859 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7324 14611 7327
rect 15286 7324 15292 7336
rect 14599 7296 15292 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 17144 7324 17172 7355
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 19429 7395 19487 7401
rect 19429 7392 19441 7395
rect 18932 7364 19441 7392
rect 18932 7352 18938 7364
rect 19429 7361 19441 7364
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 19518 7352 19524 7404
rect 19576 7392 19582 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19576 7364 19625 7392
rect 19576 7352 19582 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 21174 7392 21180 7404
rect 21087 7364 21180 7392
rect 19613 7355 19671 7361
rect 21174 7352 21180 7364
rect 21232 7392 21238 7404
rect 21358 7392 21364 7404
rect 21232 7364 21364 7392
rect 21232 7352 21238 7364
rect 21358 7352 21364 7364
rect 21416 7352 21422 7404
rect 17954 7324 17960 7336
rect 16316 7296 17172 7324
rect 17867 7296 17960 7324
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 3510 7256 3516 7268
rect 2087 7228 3516 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6914 7256 6920 7268
rect 5951 7228 6920 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 4890 7188 4896 7200
rect 4851 7160 4896 7188
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 5258 7188 5264 7200
rect 5219 7160 5264 7188
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 9030 7188 9036 7200
rect 8991 7160 9036 7188
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11330 7188 11336 7200
rect 11011 7160 11336 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 16316 7197 16344 7296
rect 17954 7284 17960 7296
rect 18012 7324 18018 7336
rect 18966 7324 18972 7336
rect 18012 7296 18972 7324
rect 18012 7284 18018 7296
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7324 20499 7327
rect 20714 7324 20720 7336
rect 20487 7296 20720 7324
rect 20487 7293 20499 7296
rect 20441 7287 20499 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 22664 7324 22692 7491
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 24949 7531 25007 7537
rect 24949 7528 24961 7531
rect 23992 7500 24961 7528
rect 23992 7488 23998 7500
rect 24949 7497 24961 7500
rect 24995 7497 25007 7531
rect 24949 7491 25007 7497
rect 22830 7420 22836 7472
rect 22888 7460 22894 7472
rect 24121 7463 24179 7469
rect 22888 7432 22954 7460
rect 22888 7420 22894 7432
rect 24121 7429 24133 7463
rect 24167 7460 24179 7463
rect 25869 7463 25927 7469
rect 25869 7460 25881 7463
rect 24167 7432 25881 7460
rect 24167 7429 24179 7432
rect 24121 7423 24179 7429
rect 25869 7429 25881 7432
rect 25915 7429 25927 7463
rect 25869 7423 25927 7429
rect 24949 7395 25007 7401
rect 24949 7392 24961 7395
rect 24596 7364 24961 7392
rect 22664 7296 24348 7324
rect 24320 7256 24348 7296
rect 24394 7284 24400 7336
rect 24452 7324 24458 7336
rect 24452 7296 24497 7324
rect 24452 7284 24458 7296
rect 24596 7256 24624 7364
rect 24949 7361 24961 7364
rect 24995 7392 25007 7395
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 24995 7364 25605 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 25593 7361 25605 7364
rect 25639 7361 25651 7395
rect 25593 7355 25651 7361
rect 24320 7228 24624 7256
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 15068 7160 16313 7188
rect 15068 7148 15074 7160
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 20898 7148 20904 7200
rect 20956 7188 20962 7200
rect 20993 7191 21051 7197
rect 20993 7188 21005 7191
rect 20956 7160 21005 7188
rect 20956 7148 20962 7160
rect 20993 7157 21005 7160
rect 21039 7157 21051 7191
rect 20993 7151 21051 7157
rect 23474 7148 23480 7200
rect 23532 7188 23538 7200
rect 24394 7188 24400 7200
rect 23532 7160 24400 7188
rect 23532 7148 23538 7160
rect 24394 7148 24400 7160
rect 24452 7148 24458 7200
rect 1104 7098 27876 7120
rect 1104 7046 4296 7098
rect 4348 7046 4360 7098
rect 4412 7046 4424 7098
rect 4476 7046 4488 7098
rect 4540 7046 4552 7098
rect 4604 7046 10988 7098
rect 11040 7046 11052 7098
rect 11104 7046 11116 7098
rect 11168 7046 11180 7098
rect 11232 7046 11244 7098
rect 11296 7046 17680 7098
rect 17732 7046 17744 7098
rect 17796 7046 17808 7098
rect 17860 7046 17872 7098
rect 17924 7046 17936 7098
rect 17988 7046 24372 7098
rect 24424 7046 24436 7098
rect 24488 7046 24500 7098
rect 24552 7046 24564 7098
rect 24616 7046 24628 7098
rect 24680 7046 27876 7098
rect 1104 7024 27876 7046
rect 4154 6984 4160 6996
rect 4115 6956 4160 6984
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 6837 6987 6895 6993
rect 6837 6984 6849 6987
rect 5408 6956 6849 6984
rect 5408 6944 5414 6956
rect 6837 6953 6849 6956
rect 6883 6953 6895 6987
rect 6837 6947 6895 6953
rect 9572 6987 9630 6993
rect 9572 6953 9584 6987
rect 9618 6984 9630 6987
rect 14369 6987 14427 6993
rect 9618 6956 11928 6984
rect 9618 6953 9630 6956
rect 9572 6947 9630 6953
rect 3421 6919 3479 6925
rect 3421 6885 3433 6919
rect 3467 6914 3479 6919
rect 3467 6886 3501 6914
rect 3467 6885 3479 6886
rect 3421 6879 3479 6885
rect 3436 6848 3464 6879
rect 4172 6848 4200 6944
rect 11900 6916 11928 6956
rect 14369 6953 14381 6987
rect 14415 6984 14427 6987
rect 15194 6984 15200 6996
rect 14415 6956 15200 6984
rect 14415 6953 14427 6956
rect 14369 6947 14427 6953
rect 15194 6944 15200 6956
rect 15252 6984 15258 6996
rect 16482 6984 16488 6996
rect 15252 6956 16488 6984
rect 15252 6944 15258 6956
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 20162 6944 20168 6996
rect 20220 6984 20226 6996
rect 21158 6987 21216 6993
rect 21158 6984 21170 6987
rect 20220 6956 21170 6984
rect 20220 6944 20226 6956
rect 21158 6953 21170 6956
rect 21204 6953 21216 6987
rect 21158 6947 21216 6953
rect 12526 6916 12532 6928
rect 11900 6888 12532 6916
rect 12526 6876 12532 6888
rect 12584 6876 12590 6928
rect 8202 6848 8208 6860
rect 3436 6820 4200 6848
rect 8163 6820 8208 6848
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 10836 6820 11713 6848
rect 10836 6808 10842 6820
rect 11701 6817 11713 6820
rect 11747 6817 11759 6851
rect 13078 6848 13084 6860
rect 13039 6820 13084 6848
rect 11701 6811 11759 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13354 6848 13360 6860
rect 13315 6820 13360 6848
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 15105 6851 15163 6857
rect 15105 6817 15117 6851
rect 15151 6848 15163 6851
rect 17037 6851 17095 6857
rect 17037 6848 17049 6851
rect 15151 6820 17049 6848
rect 15151 6817 15163 6820
rect 15105 6811 15163 6817
rect 17037 6817 17049 6820
rect 17083 6817 17095 6851
rect 18506 6848 18512 6860
rect 17037 6811 17095 6817
rect 18064 6820 18512 6848
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2308 6783 2366 6789
rect 2308 6749 2320 6783
rect 2354 6780 2366 6783
rect 5258 6780 5264 6792
rect 2354 6752 5264 6780
rect 2354 6749 2366 6752
rect 2308 6743 2366 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7190 6780 7196 6792
rect 7147 6752 7196 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9180 6752 9321 6780
rect 9180 6740 9186 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 11977 6743 12035 6749
rect 3970 6712 3976 6724
rect 3931 6684 3976 6712
rect 3970 6672 3976 6684
rect 4028 6672 4034 6724
rect 4982 6712 4988 6724
rect 4356 6684 4988 6712
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4356 6653 4384 6684
rect 4982 6672 4988 6684
rect 5040 6672 5046 6724
rect 6546 6712 6552 6724
rect 6394 6684 6552 6712
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 10594 6672 10600 6724
rect 10652 6672 10658 6724
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 11992 6712 12020 6743
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 13780 6752 14841 6780
rect 13780 6740 13786 6752
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 17218 6780 17224 6792
rect 14829 6743 14887 6749
rect 16592 6752 17224 6780
rect 11020 6684 15516 6712
rect 11020 6672 11026 6684
rect 4173 6647 4231 6653
rect 4173 6644 4185 6647
rect 4120 6616 4185 6644
rect 4120 6604 4126 6616
rect 4173 6613 4185 6616
rect 4219 6613 4231 6647
rect 4173 6607 4231 6613
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6613 4399 6647
rect 4798 6644 4804 6656
rect 4759 6616 4804 6644
rect 4341 6607 4399 6613
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5350 6644 5356 6656
rect 5224 6616 5356 6644
rect 5224 6604 5230 6616
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 11422 6644 11428 6656
rect 11103 6616 11428 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11422 6604 11428 6616
rect 11480 6644 11486 6656
rect 11882 6644 11888 6656
rect 11480 6616 11888 6644
rect 11480 6604 11486 6616
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 12618 6644 12624 6656
rect 12579 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 15488 6644 15516 6684
rect 16114 6672 16120 6724
rect 16172 6672 16178 6724
rect 16482 6644 16488 6656
rect 15488 6616 16488 6644
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16592 6653 16620 6752
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 18064 6789 18092 6820
rect 18506 6808 18512 6820
rect 18564 6848 18570 6860
rect 19334 6848 19340 6860
rect 18564 6820 19340 6848
rect 18564 6808 18570 6820
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 22646 6848 22652 6860
rect 22607 6820 22652 6848
rect 22646 6808 22652 6820
rect 22704 6848 22710 6860
rect 23385 6851 23443 6857
rect 22704 6820 23152 6848
rect 22704 6808 22710 6820
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18656 6752 18797 6780
rect 18656 6740 18662 6752
rect 18785 6749 18797 6752
rect 18831 6780 18843 6783
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 18831 6752 19717 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 19705 6749 19717 6752
rect 19751 6780 19763 6783
rect 19978 6780 19984 6792
rect 19751 6752 19984 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 20456 6712 20484 6743
rect 22278 6740 22284 6792
rect 22336 6740 22342 6792
rect 23124 6789 23152 6820
rect 23385 6817 23397 6851
rect 23431 6848 23443 6851
rect 23474 6848 23480 6860
rect 23431 6820 23480 6848
rect 23431 6817 23443 6820
rect 23385 6811 23443 6817
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 20898 6712 20904 6724
rect 20456 6684 20904 6712
rect 20898 6672 20904 6684
rect 20956 6712 20962 6724
rect 21174 6712 21180 6724
rect 20956 6684 21180 6712
rect 20956 6672 20962 6684
rect 21174 6672 21180 6684
rect 21232 6672 21238 6724
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6613 16635 6647
rect 16577 6607 16635 6613
rect 17218 6604 17224 6656
rect 17276 6644 17282 6656
rect 17865 6647 17923 6653
rect 17865 6644 17877 6647
rect 17276 6616 17877 6644
rect 17276 6604 17282 6616
rect 17865 6613 17877 6616
rect 17911 6613 17923 6647
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 17865 6607 17923 6613
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 19392 6616 19533 6644
rect 19392 6604 19398 6616
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 19702 6604 19708 6656
rect 19760 6644 19766 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 19760 6616 20269 6644
rect 19760 6604 19766 6616
rect 20257 6613 20269 6616
rect 20303 6613 20315 6647
rect 20257 6607 20315 6613
rect 1104 6554 28032 6576
rect 1104 6502 7642 6554
rect 7694 6502 7706 6554
rect 7758 6502 7770 6554
rect 7822 6502 7834 6554
rect 7886 6502 7898 6554
rect 7950 6502 14334 6554
rect 14386 6502 14398 6554
rect 14450 6502 14462 6554
rect 14514 6502 14526 6554
rect 14578 6502 14590 6554
rect 14642 6502 21026 6554
rect 21078 6502 21090 6554
rect 21142 6502 21154 6554
rect 21206 6502 21218 6554
rect 21270 6502 21282 6554
rect 21334 6502 27718 6554
rect 27770 6502 27782 6554
rect 27834 6502 27846 6554
rect 27898 6502 27910 6554
rect 27962 6502 27974 6554
rect 28026 6502 28032 6554
rect 1104 6480 28032 6502
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3970 6440 3976 6452
rect 3467 6412 3976 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 7466 6440 7472 6452
rect 6886 6412 7472 6440
rect 6886 6372 6914 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8168 6412 8769 6440
rect 8168 6400 8174 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9309 6443 9367 6449
rect 9309 6440 9321 6443
rect 9272 6412 9321 6440
rect 9272 6400 9278 6412
rect 9309 6409 9321 6412
rect 9355 6409 9367 6443
rect 11698 6440 11704 6452
rect 9309 6403 9367 6409
rect 11440 6412 11704 6440
rect 5368 6344 6914 6372
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2308 6307 2366 6313
rect 2308 6273 2320 6307
rect 2354 6304 2366 6307
rect 2866 6304 2872 6316
rect 2354 6276 2872 6304
rect 2354 6273 2366 6276
rect 2308 6267 2366 6273
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 3970 6304 3976 6316
rect 3931 6276 3976 6304
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 5368 6313 5396 6344
rect 8294 6332 8300 6384
rect 8352 6332 8358 6384
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 10873 6375 10931 6381
rect 10873 6372 10885 6375
rect 10560 6344 10885 6372
rect 10560 6332 10566 6344
rect 10873 6341 10885 6344
rect 10919 6341 10931 6375
rect 10873 6335 10931 6341
rect 5353 6307 5411 6313
rect 4120 6276 4213 6304
rect 4120 6264 4126 6276
rect 5353 6273 5365 6307
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6972 6276 7021 6304
rect 6972 6264 6978 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 10008 6276 10149 6304
rect 10008 6264 10014 6276
rect 10137 6273 10149 6276
rect 10183 6304 10195 6307
rect 10962 6304 10968 6316
rect 10183 6276 10968 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11440 6304 11468 6412
rect 11698 6400 11704 6412
rect 11756 6440 11762 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 11756 6412 13461 6440
rect 11756 6400 11762 6412
rect 13449 6409 13461 6412
rect 13495 6440 13507 6443
rect 13906 6440 13912 6452
rect 13495 6412 13912 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 15930 6440 15936 6452
rect 15891 6412 15936 6440
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16482 6400 16488 6452
rect 16540 6440 16546 6452
rect 18966 6440 18972 6452
rect 16540 6412 18972 6440
rect 16540 6400 16546 6412
rect 18966 6400 18972 6412
rect 19024 6440 19030 6452
rect 19518 6440 19524 6452
rect 19024 6412 19524 6440
rect 19024 6400 19030 6412
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 20036 6412 20821 6440
rect 20036 6400 20042 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 22830 6440 22836 6452
rect 22791 6412 22836 6440
rect 20809 6403 20867 6409
rect 22830 6400 22836 6412
rect 22888 6400 22894 6452
rect 12618 6332 12624 6384
rect 12676 6332 12682 6384
rect 17129 6375 17187 6381
rect 17129 6341 17141 6375
rect 17175 6372 17187 6375
rect 17218 6372 17224 6384
rect 17175 6344 17224 6372
rect 17175 6341 17187 6344
rect 17129 6335 17187 6341
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 17586 6332 17592 6384
rect 17644 6332 17650 6384
rect 19334 6372 19340 6384
rect 19295 6344 19340 6372
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 19610 6332 19616 6384
rect 19668 6372 19674 6384
rect 25222 6372 25228 6384
rect 19668 6344 19826 6372
rect 23492 6344 25228 6372
rect 19668 6332 19674 6344
rect 11195 6276 11468 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11664 6276 11713 6304
rect 11664 6264 11670 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 13446 6264 13452 6316
rect 13504 6304 13510 6316
rect 14001 6307 14059 6313
rect 14001 6304 14013 6307
rect 13504 6276 14013 6304
rect 13504 6264 13510 6276
rect 14001 6273 14013 6276
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15562 6304 15568 6316
rect 15523 6276 15568 6304
rect 15289 6267 15347 6273
rect 3510 6196 3516 6248
rect 3568 6236 3574 6248
rect 4080 6236 4108 6264
rect 3568 6208 4108 6236
rect 5445 6239 5503 6245
rect 3568 6196 3574 6208
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5534 6236 5540 6248
rect 5491 6208 5540 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 5994 6236 6000 6248
rect 5955 6208 6000 6236
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 8018 6236 8024 6248
rect 7331 6208 8024 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10226 6236 10232 6248
rect 9916 6208 10232 6236
rect 9916 6196 9922 6208
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 11974 6236 11980 6248
rect 11935 6208 11980 6236
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15304 6236 15332 6267
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 23492 6313 23520 6344
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 23477 6307 23535 6313
rect 23477 6304 23489 6307
rect 22296 6276 23489 6304
rect 16850 6236 16856 6248
rect 15160 6208 15608 6236
rect 16811 6208 16856 6236
rect 15160 6196 15166 6208
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 4212 6072 4261 6100
rect 4212 6060 4218 6072
rect 4249 6069 4261 6072
rect 4295 6100 4307 6103
rect 4890 6100 4896 6112
rect 4295 6072 4896 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 13998 6100 14004 6112
rect 13959 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 15580 6100 15608 6208
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18472 6208 19073 6236
rect 18472 6196 18478 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 18156 6140 18736 6168
rect 18156 6100 18184 6140
rect 15580 6072 18184 6100
rect 18506 6060 18512 6112
rect 18564 6100 18570 6112
rect 18601 6103 18659 6109
rect 18601 6100 18613 6103
rect 18564 6072 18613 6100
rect 18564 6060 18570 6072
rect 18601 6069 18613 6072
rect 18647 6069 18659 6103
rect 18708 6100 18736 6140
rect 22296 6109 22324 6276
rect 23477 6273 23489 6276
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 23845 6307 23903 6313
rect 23845 6273 23857 6307
rect 23891 6304 23903 6307
rect 25130 6304 25136 6316
rect 23891 6276 25136 6304
rect 23891 6273 23903 6276
rect 23845 6267 23903 6273
rect 25130 6264 25136 6276
rect 25188 6264 25194 6316
rect 22281 6103 22339 6109
rect 22281 6100 22293 6103
rect 18708 6072 22293 6100
rect 18601 6063 18659 6069
rect 22281 6069 22293 6072
rect 22327 6069 22339 6103
rect 22281 6063 22339 6069
rect 1104 6010 27876 6032
rect 1104 5958 4296 6010
rect 4348 5958 4360 6010
rect 4412 5958 4424 6010
rect 4476 5958 4488 6010
rect 4540 5958 4552 6010
rect 4604 5958 10988 6010
rect 11040 5958 11052 6010
rect 11104 5958 11116 6010
rect 11168 5958 11180 6010
rect 11232 5958 11244 6010
rect 11296 5958 17680 6010
rect 17732 5958 17744 6010
rect 17796 5958 17808 6010
rect 17860 5958 17872 6010
rect 17924 5958 17936 6010
rect 17988 5958 24372 6010
rect 24424 5958 24436 6010
rect 24488 5958 24500 6010
rect 24552 5958 24564 6010
rect 24616 5958 24628 6010
rect 24680 5958 27876 6010
rect 1104 5936 27876 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 2372 5868 2421 5896
rect 2372 5856 2378 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2924 5868 2973 5896
rect 2924 5856 2930 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4764 5868 4813 5896
rect 4764 5856 4770 5868
rect 4801 5865 4813 5868
rect 4847 5865 4859 5899
rect 4801 5859 4859 5865
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 6328 5868 7389 5896
rect 6328 5856 6334 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 7377 5859 7435 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 11320 5899 11378 5905
rect 11320 5865 11332 5899
rect 11366 5896 11378 5899
rect 13998 5896 14004 5908
rect 11366 5868 14004 5896
rect 11366 5865 11378 5868
rect 11320 5859 11378 5865
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 18414 5896 18420 5908
rect 18375 5868 18420 5896
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 21177 5899 21235 5905
rect 21177 5896 21189 5899
rect 20956 5868 21189 5896
rect 20956 5856 20962 5868
rect 21177 5865 21189 5868
rect 21223 5865 21235 5899
rect 21177 5859 21235 5865
rect 2332 5828 2360 5856
rect 1596 5800 2360 5828
rect 1596 5701 1624 5800
rect 2774 5788 2780 5840
rect 2832 5828 2838 5840
rect 3973 5831 4031 5837
rect 3973 5828 3985 5831
rect 2832 5800 3985 5828
rect 2832 5788 2838 5800
rect 3973 5797 3985 5800
rect 4019 5797 4031 5831
rect 3973 5791 4031 5797
rect 12805 5831 12863 5837
rect 12805 5797 12817 5831
rect 12851 5828 12863 5831
rect 13446 5828 13452 5840
rect 12851 5800 13452 5828
rect 12851 5797 12863 5800
rect 12805 5791 12863 5797
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 13722 5828 13728 5840
rect 13683 5800 13728 5828
rect 13722 5788 13728 5800
rect 13780 5788 13786 5840
rect 3421 5763 3479 5769
rect 1780 5732 3372 5760
rect 1780 5701 1808 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2225 5695 2283 5701
rect 2225 5692 2237 5695
rect 2188 5664 2237 5692
rect 2188 5652 2194 5664
rect 2225 5661 2237 5664
rect 2271 5661 2283 5695
rect 3142 5692 3148 5704
rect 3103 5664 3148 5692
rect 2225 5655 2283 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3344 5701 3372 5732
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 3878 5760 3884 5772
rect 3467 5732 3884 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 5902 5760 5908 5772
rect 3988 5732 5028 5760
rect 5863 5732 5908 5760
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5692 3387 5695
rect 3510 5692 3516 5704
rect 3375 5664 3516 5692
rect 3375 5661 3387 5664
rect 3329 5655 3387 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3988 5701 4016 5732
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 1673 5627 1731 5633
rect 1673 5593 1685 5627
rect 1719 5624 1731 5627
rect 3050 5624 3056 5636
rect 1719 5596 3056 5624
rect 1719 5593 1731 5596
rect 1673 5587 1731 5593
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 3988 5556 4016 5655
rect 4264 5624 4292 5655
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 5000 5701 5028 5732
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 10594 5760 10600 5772
rect 10555 5732 10600 5760
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 11057 5763 11115 5769
rect 11057 5729 11069 5763
rect 11103 5760 11115 5763
rect 11330 5760 11336 5772
rect 11103 5732 11336 5760
rect 11103 5729 11115 5732
rect 11057 5723 11115 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 13648 5732 14565 5760
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4672 5664 4813 5692
rect 4672 5652 4678 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 5626 5692 5632 5704
rect 5587 5664 5632 5692
rect 4985 5655 5043 5661
rect 4706 5624 4712 5636
rect 4264 5596 4712 5624
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 2372 5528 4016 5556
rect 2372 5516 2378 5528
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 4120 5528 4169 5556
rect 4120 5516 4126 5528
rect 4157 5525 4169 5528
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5000 5556 5028 5655
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 8846 5692 8852 5704
rect 8168 5664 8852 5692
rect 8168 5652 8174 5664
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 9950 5692 9956 5704
rect 9911 5664 9956 5692
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10226 5692 10232 5704
rect 10139 5664 10232 5692
rect 10226 5652 10232 5664
rect 10284 5692 10290 5704
rect 10778 5692 10784 5704
rect 10284 5664 10784 5692
rect 10284 5652 10290 5664
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 5994 5584 6000 5636
rect 6052 5624 6058 5636
rect 6052 5596 6394 5624
rect 6052 5584 6058 5596
rect 11790 5584 11796 5636
rect 11848 5584 11854 5636
rect 6822 5556 6828 5568
rect 4948 5528 6828 5556
rect 4948 5516 4954 5528
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 13648 5556 13676 5732
rect 14553 5729 14565 5732
rect 14599 5760 14611 5763
rect 16114 5760 16120 5772
rect 14599 5732 15148 5760
rect 16075 5732 16120 5760
rect 14599 5729 14611 5732
rect 14553 5723 14611 5729
rect 15120 5704 15148 5732
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17681 5763 17739 5769
rect 17681 5760 17693 5763
rect 17644 5732 17693 5760
rect 17644 5720 17650 5732
rect 17681 5729 17693 5732
rect 17727 5729 17739 5763
rect 17681 5723 17739 5729
rect 18782 5720 18788 5772
rect 18840 5760 18846 5772
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 18840 5732 19441 5760
rect 18840 5720 18846 5732
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19702 5760 19708 5772
rect 19663 5732 19708 5760
rect 19429 5723 19487 5729
rect 19702 5720 19708 5732
rect 19760 5720 19766 5772
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 15010 5692 15016 5704
rect 13771 5664 15016 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 15160 5664 15301 5692
rect 15160 5652 15166 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 15620 5664 15761 5692
rect 15620 5652 15626 5664
rect 15749 5661 15761 5664
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 15764 5624 15792 5655
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 16945 5695 17003 5701
rect 16945 5692 16957 5695
rect 16540 5664 16957 5692
rect 16540 5652 16546 5664
rect 16945 5661 16957 5664
rect 16991 5661 17003 5695
rect 16945 5655 17003 5661
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 18506 5692 18512 5704
rect 18463 5664 18512 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 17420 5624 17448 5655
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 18874 5624 18880 5636
rect 15764 5596 18880 5624
rect 18874 5584 18880 5596
rect 18932 5584 18938 5636
rect 20714 5584 20720 5636
rect 20772 5584 20778 5636
rect 8260 5528 13676 5556
rect 8260 5516 8266 5528
rect 1104 5466 28032 5488
rect 1104 5414 7642 5466
rect 7694 5414 7706 5466
rect 7758 5414 7770 5466
rect 7822 5414 7834 5466
rect 7886 5414 7898 5466
rect 7950 5414 14334 5466
rect 14386 5414 14398 5466
rect 14450 5414 14462 5466
rect 14514 5414 14526 5466
rect 14578 5414 14590 5466
rect 14642 5414 21026 5466
rect 21078 5414 21090 5466
rect 21142 5414 21154 5466
rect 21206 5414 21218 5466
rect 21270 5414 21282 5466
rect 21334 5414 27718 5466
rect 27770 5414 27782 5466
rect 27834 5414 27846 5466
rect 27898 5414 27910 5466
rect 27962 5414 27974 5466
rect 28026 5414 28032 5466
rect 1104 5392 28032 5414
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5352 2099 5355
rect 3142 5352 3148 5364
rect 2087 5324 3148 5352
rect 2087 5321 2099 5324
rect 2041 5315 2099 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 6641 5355 6699 5361
rect 6641 5321 6653 5355
rect 6687 5352 6699 5355
rect 7190 5352 7196 5364
rect 6687 5324 7196 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8294 5352 8300 5364
rect 8255 5324 8300 5352
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 11790 5352 11796 5364
rect 11195 5324 11796 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12526 5352 12532 5364
rect 12487 5324 12532 5352
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 14921 5355 14979 5361
rect 14921 5321 14933 5355
rect 14967 5352 14979 5355
rect 15102 5352 15108 5364
rect 14967 5324 15108 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 18693 5355 18751 5361
rect 18693 5321 18705 5355
rect 18739 5352 18751 5355
rect 18874 5352 18880 5364
rect 18739 5324 18880 5352
rect 18739 5321 18751 5324
rect 18693 5315 18751 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 2314 5284 2320 5296
rect 1964 5256 2320 5284
rect 1964 5225 1992 5256
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 4154 5284 4160 5296
rect 2746 5256 4160 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2746 5216 2774 5256
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 4709 5287 4767 5293
rect 4709 5253 4721 5287
rect 4755 5284 4767 5287
rect 4890 5284 4896 5296
rect 4755 5256 4896 5284
rect 4755 5253 4767 5256
rect 4709 5247 4767 5253
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 9122 5284 9128 5296
rect 9083 5256 9128 5284
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 11974 5284 11980 5296
rect 11935 5256 11980 5284
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 16850 5284 16856 5296
rect 16811 5256 16856 5284
rect 16850 5244 16856 5256
rect 16908 5244 16914 5296
rect 19981 5287 20039 5293
rect 19981 5253 19993 5287
rect 20027 5284 20039 5287
rect 20806 5284 20812 5296
rect 20027 5256 20812 5284
rect 20027 5253 20039 5256
rect 19981 5247 20039 5253
rect 20806 5244 20812 5256
rect 20864 5244 20870 5296
rect 2866 5225 2872 5228
rect 2179 5188 2774 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2860 5179 2872 5225
rect 2924 5216 2930 5228
rect 4433 5219 4491 5225
rect 2924 5188 2960 5216
rect 2866 5176 2872 5179
rect 2924 5176 2930 5188
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4982 5216 4988 5228
rect 4479 5188 4988 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5408 5188 5641 5216
rect 5408 5176 5414 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 6236 5188 6745 5216
rect 6236 5176 6242 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7650 5216 7656 5228
rect 7524 5188 7656 5216
rect 7524 5176 7530 5188
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8846 5216 8852 5228
rect 8807 5188 8852 5216
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10008 5188 10333 5216
rect 10008 5176 10014 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10778 5216 10784 5228
rect 10739 5188 10784 5216
rect 10321 5179 10379 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 11940 5188 12449 5216
rect 11940 5176 11946 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 12437 5179 12495 5185
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2590 5148 2596 5160
rect 2096 5120 2596 5148
rect 2096 5108 2102 5120
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 7098 5148 7104 5160
rect 5592 5120 7104 5148
rect 5592 5108 5598 5120
rect 7098 5108 7104 5120
rect 7156 5148 7162 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 7156 5120 7389 5148
rect 7156 5108 7162 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 4525 5083 4583 5089
rect 4525 5049 4537 5083
rect 4571 5080 4583 5083
rect 4614 5080 4620 5092
rect 4571 5052 4620 5080
rect 4571 5049 4583 5052
rect 4525 5043 4583 5049
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 3970 5012 3976 5024
rect 3931 4984 3976 5012
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 4212 4984 4445 5012
rect 4212 4972 4218 4984
rect 4433 4981 4445 4984
rect 4479 4981 4491 5015
rect 4433 4975 4491 4981
rect 1104 4922 27876 4944
rect 1104 4870 4296 4922
rect 4348 4870 4360 4922
rect 4412 4870 4424 4922
rect 4476 4870 4488 4922
rect 4540 4870 4552 4922
rect 4604 4870 10988 4922
rect 11040 4870 11052 4922
rect 11104 4870 11116 4922
rect 11168 4870 11180 4922
rect 11232 4870 11244 4922
rect 11296 4870 17680 4922
rect 17732 4870 17744 4922
rect 17796 4870 17808 4922
rect 17860 4870 17872 4922
rect 17924 4870 17936 4922
rect 17988 4870 24372 4922
rect 24424 4870 24436 4922
rect 24488 4870 24500 4922
rect 24552 4870 24564 4922
rect 24616 4870 24628 4922
rect 24680 4870 27876 4922
rect 1104 4848 27876 4870
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3568 4780 3985 4808
rect 3568 4768 3574 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 3973 4771 4031 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 8628 4780 9137 4808
rect 8628 4768 8634 4780
rect 9125 4777 9137 4780
rect 9171 4777 9183 4811
rect 9125 4771 9183 4777
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 10836 4780 11713 4808
rect 10836 4768 10842 4780
rect 11701 4777 11713 4780
rect 11747 4777 11759 4811
rect 11701 4771 11759 4777
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 3418 4740 3424 4752
rect 2455 4712 3424 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 3418 4700 3424 4712
rect 3476 4700 3482 4752
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 4525 4743 4583 4749
rect 4525 4740 4537 4743
rect 4120 4712 4537 4740
rect 4120 4700 4126 4712
rect 4525 4709 4537 4712
rect 4571 4709 4583 4743
rect 4525 4703 4583 4709
rect 2774 4672 2780 4684
rect 2240 4644 2780 4672
rect 2240 4613 2268 4644
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3329 4675 3387 4681
rect 3108 4644 3188 4672
rect 3108 4632 3114 4644
rect 3160 4613 3188 4644
rect 3329 4641 3341 4675
rect 3375 4672 3387 4675
rect 4982 4672 4988 4684
rect 3375 4644 4988 4672
rect 3375 4641 3387 4644
rect 3329 4635 3387 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 8205 4675 8263 4681
rect 8205 4672 8217 4675
rect 7708 4644 8217 4672
rect 7708 4632 7714 4644
rect 8205 4641 8217 4644
rect 8251 4672 8263 4675
rect 9950 4672 9956 4684
rect 8251 4644 9956 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 3145 4607 3203 4613
rect 2547 4576 2820 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2792 4548 2820 4576
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3878 4604 3884 4616
rect 3467 4576 3884 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3878 4564 3884 4576
rect 3936 4604 3942 4616
rect 4157 4607 4215 4613
rect 4157 4604 4169 4607
rect 3936 4576 4169 4604
rect 3936 4564 3942 4576
rect 4157 4573 4169 4576
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 5166 4604 5172 4616
rect 4295 4576 5172 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 7558 4604 7564 4616
rect 7519 4576 7564 4604
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 9030 4604 9036 4616
rect 8312 4576 9036 4604
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 3970 4536 3976 4548
rect 2832 4508 3976 4536
rect 2832 4496 2838 4508
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 7009 4539 7067 4545
rect 7009 4505 7021 4539
rect 7055 4536 7067 4539
rect 8312 4536 8340 4576
rect 9030 4564 9036 4576
rect 9088 4604 9094 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 9088 4576 10425 4604
rect 9088 4564 9094 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 7055 4508 8340 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 2041 4471 2099 4477
rect 2041 4437 2053 4471
rect 2087 4468 2099 4471
rect 2314 4468 2320 4480
rect 2087 4440 2320 4468
rect 2087 4437 2099 4440
rect 2041 4431 2099 4437
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2958 4468 2964 4480
rect 2919 4440 2964 4468
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 4338 4468 4344 4480
rect 3476 4440 4344 4468
rect 3476 4428 3482 4440
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 9858 4468 9864 4480
rect 9819 4440 9864 4468
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 1104 4378 28032 4400
rect 1104 4326 7642 4378
rect 7694 4326 7706 4378
rect 7758 4326 7770 4378
rect 7822 4326 7834 4378
rect 7886 4326 7898 4378
rect 7950 4326 14334 4378
rect 14386 4326 14398 4378
rect 14450 4326 14462 4378
rect 14514 4326 14526 4378
rect 14578 4326 14590 4378
rect 14642 4326 21026 4378
rect 21078 4326 21090 4378
rect 21142 4326 21154 4378
rect 21206 4326 21218 4378
rect 21270 4326 21282 4378
rect 21334 4326 27718 4378
rect 27770 4326 27782 4378
rect 27834 4326 27846 4378
rect 27898 4326 27910 4378
rect 27962 4326 27974 4378
rect 28026 4326 28032 4378
rect 1104 4304 28032 4326
rect 3878 4224 3884 4276
rect 3936 4264 3942 4276
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 3936 4236 4261 4264
rect 3936 4224 3942 4236
rect 4249 4233 4261 4236
rect 4295 4233 4307 4267
rect 4982 4264 4988 4276
rect 4943 4236 4988 4264
rect 4249 4227 4307 4233
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 5092 4236 5396 4264
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3114 4199 3172 4205
rect 3114 4196 3126 4199
rect 3016 4168 3126 4196
rect 3016 4156 3022 4168
rect 3114 4165 3126 4168
rect 3160 4165 3172 4199
rect 3114 4159 3172 4165
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 5092 4196 5120 4236
rect 5166 4205 5172 4208
rect 4120 4168 5120 4196
rect 5153 4199 5172 4205
rect 4120 4156 4126 4168
rect 5153 4165 5165 4199
rect 5153 4159 5172 4165
rect 5166 4156 5172 4159
rect 5224 4156 5230 4208
rect 5368 4205 5396 4236
rect 5353 4199 5411 4205
rect 5353 4165 5365 4199
rect 5399 4165 5411 4199
rect 5353 4159 5411 4165
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1544 4100 1593 4128
rect 1544 4088 1550 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 1581 4091 1639 4097
rect 1596 3992 1624 4091
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2774 4128 2780 4140
rect 2455 4100 2780 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7374 4128 7380 4140
rect 7147 4100 7380 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7374 4088 7380 4100
rect 7432 4128 7438 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 7432 4100 7573 4128
rect 7432 4088 7438 4100
rect 7561 4097 7573 4100
rect 7607 4128 7619 4131
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 7607 4100 8953 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 18966 4128 18972 4140
rect 18927 4100 18972 4128
rect 8941 4091 8999 4097
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19610 4128 19616 4140
rect 19571 4100 19616 4128
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 2590 4020 2596 4072
rect 2648 4060 2654 4072
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2648 4032 2881 4060
rect 2648 4020 2654 4032
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 18874 4060 18880 4072
rect 18835 4032 18880 4060
rect 2869 4023 2927 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 2774 3992 2780 4004
rect 1596 3964 2780 3992
rect 2774 3952 2780 3964
rect 2832 3952 2838 4004
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 9858 3992 9864 4004
rect 5951 3964 9864 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 2130 3924 2136 3936
rect 1811 3896 2136 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 2866 3924 2872 3936
rect 2271 3896 2872 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4706 3924 4712 3936
rect 4396 3896 4712 3924
rect 4396 3884 4402 3896
rect 4706 3884 4712 3896
rect 4764 3924 4770 3936
rect 5169 3927 5227 3933
rect 5169 3924 5181 3927
rect 4764 3896 5181 3924
rect 4764 3884 4770 3896
rect 5169 3893 5181 3896
rect 5215 3893 5227 3927
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 5169 3887 5227 3893
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 1104 3834 27876 3856
rect 1104 3782 4296 3834
rect 4348 3782 4360 3834
rect 4412 3782 4424 3834
rect 4476 3782 4488 3834
rect 4540 3782 4552 3834
rect 4604 3782 10988 3834
rect 11040 3782 11052 3834
rect 11104 3782 11116 3834
rect 11168 3782 11180 3834
rect 11232 3782 11244 3834
rect 11296 3782 17680 3834
rect 17732 3782 17744 3834
rect 17796 3782 17808 3834
rect 17860 3782 17872 3834
rect 17924 3782 17936 3834
rect 17988 3782 24372 3834
rect 24424 3782 24436 3834
rect 24488 3782 24500 3834
rect 24552 3782 24564 3834
rect 24616 3782 24628 3834
rect 24680 3782 27876 3834
rect 1104 3760 27876 3782
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 4614 3720 4620 3732
rect 4295 3692 4620 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 4798 3720 4804 3732
rect 4759 3692 4804 3720
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5353 3723 5411 3729
rect 5353 3689 5365 3723
rect 5399 3720 5411 3723
rect 5442 3720 5448 3732
rect 5399 3692 5448 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5776 3692 5917 3720
rect 5776 3680 5782 3692
rect 5905 3689 5917 3692
rect 5951 3720 5963 3723
rect 6457 3723 6515 3729
rect 6457 3720 6469 3723
rect 5951 3692 6469 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 6457 3689 6469 3692
rect 6503 3720 6515 3723
rect 6822 3720 6828 3732
rect 6503 3692 6828 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6822 3680 6828 3692
rect 6880 3720 6886 3732
rect 6880 3680 6914 3720
rect 2038 3516 2044 3528
rect 1951 3488 2044 3516
rect 2038 3476 2044 3488
rect 2096 3516 2102 3528
rect 2590 3516 2596 3528
rect 2096 3488 2596 3516
rect 2096 3476 2102 3488
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 3436 3516 3464 3680
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3436 3488 3985 3516
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4249 3519 4307 3525
rect 4120 3488 4165 3516
rect 4120 3476 4126 3488
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 5166 3516 5172 3528
rect 4295 3488 5172 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 6886 3516 6914 3680
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6886 3488 7021 3516
rect 7009 3485 7021 3488
rect 7055 3516 7067 3519
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7055 3488 7941 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 2314 3457 2320 3460
rect 2308 3448 2320 3457
rect 2275 3420 2320 3448
rect 2308 3411 2320 3420
rect 2314 3408 2320 3411
rect 2372 3408 2378 3460
rect 1104 3290 28032 3312
rect 1104 3238 7642 3290
rect 7694 3238 7706 3290
rect 7758 3238 7770 3290
rect 7822 3238 7834 3290
rect 7886 3238 7898 3290
rect 7950 3238 14334 3290
rect 14386 3238 14398 3290
rect 14450 3238 14462 3290
rect 14514 3238 14526 3290
rect 14578 3238 14590 3290
rect 14642 3238 21026 3290
rect 21078 3238 21090 3290
rect 21142 3238 21154 3290
rect 21206 3238 21218 3290
rect 21270 3238 21282 3290
rect 21334 3238 27718 3290
rect 27770 3238 27782 3290
rect 27834 3238 27846 3290
rect 27898 3238 27910 3290
rect 27962 3238 27974 3290
rect 28026 3238 28032 3290
rect 1104 3216 28032 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5718 3176 5724 3188
rect 5679 3148 5724 3176
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 3326 3108 3332 3120
rect 3287 3080 3332 3108
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 4056 3111 4114 3117
rect 4056 3077 4068 3111
rect 4102 3108 4114 3111
rect 4154 3108 4160 3120
rect 4102 3080 4160 3108
rect 4102 3077 4114 3080
rect 4056 3071 4114 3077
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 2832 3012 6561 3040
rect 2832 3000 2838 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 2648 2944 3801 2972
rect 2648 2932 2654 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 1104 2746 27876 2768
rect 1104 2694 4296 2746
rect 4348 2694 4360 2746
rect 4412 2694 4424 2746
rect 4476 2694 4488 2746
rect 4540 2694 4552 2746
rect 4604 2694 10988 2746
rect 11040 2694 11052 2746
rect 11104 2694 11116 2746
rect 11168 2694 11180 2746
rect 11232 2694 11244 2746
rect 11296 2694 17680 2746
rect 17732 2694 17744 2746
rect 17796 2694 17808 2746
rect 17860 2694 17872 2746
rect 17924 2694 17936 2746
rect 17988 2694 24372 2746
rect 24424 2694 24436 2746
rect 24488 2694 24500 2746
rect 24552 2694 24564 2746
rect 24616 2694 24628 2746
rect 24680 2694 27876 2746
rect 1104 2672 27876 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 2225 2635 2283 2641
rect 2225 2601 2237 2635
rect 2271 2632 2283 2635
rect 3050 2632 3056 2644
rect 2271 2604 3056 2632
rect 2271 2601 2283 2604
rect 2225 2595 2283 2601
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3660 2604 3985 2632
rect 3660 2592 3666 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5718 2632 5724 2644
rect 5215 2604 5724 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 3786 2524 3792 2576
rect 3844 2564 3850 2576
rect 4525 2567 4583 2573
rect 4525 2564 4537 2567
rect 3844 2536 4537 2564
rect 3844 2524 3850 2536
rect 4525 2533 4537 2536
rect 4571 2564 4583 2567
rect 8110 2564 8116 2576
rect 4571 2536 8116 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2496 2835 2499
rect 5718 2496 5724 2508
rect 2823 2468 5724 2496
rect 2823 2465 2835 2468
rect 2777 2459 2835 2465
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 3234 2292 3240 2304
rect 3195 2264 3240 2292
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 1104 2202 28032 2224
rect 1104 2150 7642 2202
rect 7694 2150 7706 2202
rect 7758 2150 7770 2202
rect 7822 2150 7834 2202
rect 7886 2150 7898 2202
rect 7950 2150 14334 2202
rect 14386 2150 14398 2202
rect 14450 2150 14462 2202
rect 14514 2150 14526 2202
rect 14578 2150 14590 2202
rect 14642 2150 21026 2202
rect 21078 2150 21090 2202
rect 21142 2150 21154 2202
rect 21206 2150 21218 2202
rect 21270 2150 21282 2202
rect 21334 2150 27718 2202
rect 27770 2150 27782 2202
rect 27834 2150 27846 2202
rect 27898 2150 27910 2202
rect 27962 2150 27974 2202
rect 28026 2150 28032 2202
rect 1104 2128 28032 2150
<< via1 >>
rect 4296 26630 4348 26682
rect 4360 26630 4412 26682
rect 4424 26630 4476 26682
rect 4488 26630 4540 26682
rect 4552 26630 4604 26682
rect 10988 26630 11040 26682
rect 11052 26630 11104 26682
rect 11116 26630 11168 26682
rect 11180 26630 11232 26682
rect 11244 26630 11296 26682
rect 17680 26630 17732 26682
rect 17744 26630 17796 26682
rect 17808 26630 17860 26682
rect 17872 26630 17924 26682
rect 17936 26630 17988 26682
rect 24372 26630 24424 26682
rect 24436 26630 24488 26682
rect 24500 26630 24552 26682
rect 24564 26630 24616 26682
rect 24628 26630 24680 26682
rect 1860 26528 1912 26580
rect 5448 26528 5500 26580
rect 9036 26528 9088 26580
rect 19800 26528 19852 26580
rect 23480 26528 23532 26580
rect 26976 26528 27028 26580
rect 5724 26392 5776 26444
rect 15292 26435 15344 26444
rect 1676 26367 1728 26376
rect 1676 26333 1685 26367
rect 1685 26333 1719 26367
rect 1719 26333 1728 26367
rect 1676 26324 1728 26333
rect 4528 26324 4580 26376
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 15292 26392 15344 26401
rect 6552 26367 6604 26376
rect 6552 26333 6561 26367
rect 6561 26333 6595 26367
rect 6595 26333 6604 26367
rect 6552 26324 6604 26333
rect 9128 26367 9180 26376
rect 5080 26256 5132 26308
rect 5356 26256 5408 26308
rect 6368 26256 6420 26308
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 9404 26324 9456 26376
rect 9496 26256 9548 26308
rect 13636 26324 13688 26376
rect 13820 26324 13872 26376
rect 15752 26324 15804 26376
rect 16856 26367 16908 26376
rect 16856 26333 16865 26367
rect 16865 26333 16899 26367
rect 16899 26333 16908 26367
rect 16856 26324 16908 26333
rect 19340 26324 19392 26376
rect 20168 26367 20220 26376
rect 20168 26333 20177 26367
rect 20177 26333 20211 26367
rect 20211 26333 20220 26367
rect 20168 26324 20220 26333
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 12532 26256 12584 26308
rect 13268 26256 13320 26308
rect 16120 26299 16172 26308
rect 16120 26265 16129 26299
rect 16129 26265 16163 26299
rect 16163 26265 16172 26299
rect 16120 26256 16172 26265
rect 19432 26299 19484 26308
rect 19432 26265 19441 26299
rect 19441 26265 19475 26299
rect 19475 26265 19484 26299
rect 19432 26256 19484 26265
rect 5908 26188 5960 26240
rect 9864 26188 9916 26240
rect 12624 26188 12676 26240
rect 16212 26188 16264 26240
rect 7642 26086 7694 26138
rect 7706 26086 7758 26138
rect 7770 26086 7822 26138
rect 7834 26086 7886 26138
rect 7898 26086 7950 26138
rect 14334 26086 14386 26138
rect 14398 26086 14450 26138
rect 14462 26086 14514 26138
rect 14526 26086 14578 26138
rect 14590 26086 14642 26138
rect 21026 26086 21078 26138
rect 21090 26086 21142 26138
rect 21154 26086 21206 26138
rect 21218 26086 21270 26138
rect 21282 26086 21334 26138
rect 27718 26086 27770 26138
rect 27782 26086 27834 26138
rect 27846 26086 27898 26138
rect 27910 26086 27962 26138
rect 27974 26086 28026 26138
rect 1676 26027 1728 26036
rect 1676 25993 1685 26027
rect 1685 25993 1719 26027
rect 1719 25993 1728 26027
rect 1676 25984 1728 25993
rect 4528 26027 4580 26036
rect 4528 25993 4537 26027
rect 4537 25993 4571 26027
rect 4571 25993 4580 26027
rect 4528 25984 4580 25993
rect 4988 25984 5040 26036
rect 9128 25984 9180 26036
rect 13820 25916 13872 25968
rect 14096 25916 14148 25968
rect 2964 25848 3016 25900
rect 5448 25891 5500 25900
rect 2504 25823 2556 25832
rect 2504 25789 2513 25823
rect 2513 25789 2547 25823
rect 2547 25789 2556 25823
rect 2504 25780 2556 25789
rect 5448 25857 5457 25891
rect 5457 25857 5491 25891
rect 5491 25857 5500 25891
rect 5448 25848 5500 25857
rect 6736 25891 6788 25900
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 9772 25891 9824 25900
rect 4804 25780 4856 25832
rect 5908 25780 5960 25832
rect 7380 25780 7432 25832
rect 2228 25687 2280 25696
rect 2228 25653 2237 25687
rect 2237 25653 2271 25687
rect 2271 25653 2280 25687
rect 2228 25644 2280 25653
rect 7012 25644 7064 25696
rect 7104 25644 7156 25696
rect 9772 25857 9781 25891
rect 9781 25857 9815 25891
rect 9815 25857 9824 25891
rect 9772 25848 9824 25857
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 12072 25891 12124 25900
rect 12072 25857 12081 25891
rect 12081 25857 12115 25891
rect 12115 25857 12124 25891
rect 12072 25848 12124 25857
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 17316 25848 17368 25900
rect 19340 25848 19392 25900
rect 19892 25848 19944 25900
rect 9864 25823 9916 25832
rect 9864 25789 9873 25823
rect 9873 25789 9907 25823
rect 9907 25789 9916 25823
rect 9864 25780 9916 25789
rect 10692 25823 10744 25832
rect 10692 25789 10701 25823
rect 10701 25789 10735 25823
rect 10735 25789 10744 25823
rect 10692 25780 10744 25789
rect 14188 25780 14240 25832
rect 15016 25823 15068 25832
rect 15016 25789 15025 25823
rect 15025 25789 15059 25823
rect 15059 25789 15068 25823
rect 15016 25780 15068 25789
rect 15292 25780 15344 25832
rect 20076 25780 20128 25832
rect 20812 25780 20864 25832
rect 11336 25644 11388 25696
rect 11888 25687 11940 25696
rect 11888 25653 11897 25687
rect 11897 25653 11931 25687
rect 11931 25653 11940 25687
rect 11888 25644 11940 25653
rect 16856 25712 16908 25764
rect 15476 25687 15528 25696
rect 15476 25653 15485 25687
rect 15485 25653 15519 25687
rect 15519 25653 15528 25687
rect 15476 25644 15528 25653
rect 17132 25687 17184 25696
rect 17132 25653 17141 25687
rect 17141 25653 17175 25687
rect 17175 25653 17184 25687
rect 17132 25644 17184 25653
rect 18604 25687 18656 25696
rect 18604 25653 18613 25687
rect 18613 25653 18647 25687
rect 18647 25653 18656 25687
rect 18604 25644 18656 25653
rect 4296 25542 4348 25594
rect 4360 25542 4412 25594
rect 4424 25542 4476 25594
rect 4488 25542 4540 25594
rect 4552 25542 4604 25594
rect 10988 25542 11040 25594
rect 11052 25542 11104 25594
rect 11116 25542 11168 25594
rect 11180 25542 11232 25594
rect 11244 25542 11296 25594
rect 17680 25542 17732 25594
rect 17744 25542 17796 25594
rect 17808 25542 17860 25594
rect 17872 25542 17924 25594
rect 17936 25542 17988 25594
rect 24372 25542 24424 25594
rect 24436 25542 24488 25594
rect 24500 25542 24552 25594
rect 24564 25542 24616 25594
rect 24628 25542 24680 25594
rect 4804 25483 4856 25492
rect 4804 25449 4813 25483
rect 4813 25449 4847 25483
rect 4847 25449 4856 25483
rect 4804 25440 4856 25449
rect 4160 25372 4212 25424
rect 12716 25440 12768 25492
rect 5540 25372 5592 25424
rect 7380 25415 7432 25424
rect 7380 25381 7389 25415
rect 7389 25381 7423 25415
rect 7423 25381 7432 25415
rect 7380 25372 7432 25381
rect 9404 25415 9456 25424
rect 9404 25381 9413 25415
rect 9413 25381 9447 25415
rect 9447 25381 9456 25415
rect 9404 25372 9456 25381
rect 5448 25304 5500 25356
rect 7104 25304 7156 25356
rect 9588 25304 9640 25356
rect 11888 25347 11940 25356
rect 11888 25313 11897 25347
rect 11897 25313 11931 25347
rect 11931 25313 11940 25347
rect 11888 25304 11940 25313
rect 20168 25440 20220 25492
rect 19432 25347 19484 25356
rect 19432 25313 19441 25347
rect 19441 25313 19475 25347
rect 19475 25313 19484 25347
rect 19432 25304 19484 25313
rect 20720 25304 20772 25356
rect 20904 25304 20956 25356
rect 2044 25279 2096 25288
rect 2044 25245 2053 25279
rect 2053 25245 2087 25279
rect 2087 25245 2096 25279
rect 2044 25236 2096 25245
rect 4344 25279 4396 25288
rect 4344 25245 4353 25279
rect 4353 25245 4387 25279
rect 4387 25245 4396 25279
rect 4344 25236 4396 25245
rect 4712 25236 4764 25288
rect 1676 25168 1728 25220
rect 4804 25211 4856 25220
rect 4804 25177 4813 25211
rect 4813 25177 4847 25211
rect 4847 25177 4856 25211
rect 4804 25168 4856 25177
rect 5724 25236 5776 25288
rect 5908 25279 5960 25288
rect 5908 25245 5917 25279
rect 5917 25245 5951 25279
rect 5951 25245 5960 25279
rect 5908 25236 5960 25245
rect 6552 25236 6604 25288
rect 8484 25236 8536 25288
rect 9128 25236 9180 25288
rect 9496 25279 9548 25288
rect 5816 25168 5868 25220
rect 7380 25168 7432 25220
rect 8116 25211 8168 25220
rect 8116 25177 8125 25211
rect 8125 25177 8159 25211
rect 8159 25177 8168 25211
rect 8116 25168 8168 25177
rect 8300 25168 8352 25220
rect 8852 25168 8904 25220
rect 5632 25100 5684 25152
rect 6368 25143 6420 25152
rect 6368 25109 6377 25143
rect 6377 25109 6411 25143
rect 6411 25109 6420 25143
rect 6368 25100 6420 25109
rect 9220 25100 9272 25152
rect 9496 25245 9505 25279
rect 9505 25245 9539 25279
rect 9539 25245 9548 25279
rect 9496 25236 9548 25245
rect 10692 25236 10744 25288
rect 10876 25279 10928 25288
rect 10876 25245 10885 25279
rect 10885 25245 10919 25279
rect 10919 25245 10928 25279
rect 10876 25236 10928 25245
rect 13268 25236 13320 25288
rect 15568 25236 15620 25288
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 20812 25236 20864 25288
rect 12440 25168 12492 25220
rect 14924 25211 14976 25220
rect 14924 25177 14933 25211
rect 14933 25177 14967 25211
rect 14967 25177 14976 25211
rect 14924 25168 14976 25177
rect 16580 25168 16632 25220
rect 17592 25168 17644 25220
rect 18328 25168 18380 25220
rect 10692 25143 10744 25152
rect 10692 25109 10701 25143
rect 10701 25109 10735 25143
rect 10735 25109 10744 25143
rect 10692 25100 10744 25109
rect 14004 25100 14056 25152
rect 15108 25100 15160 25152
rect 15292 25100 15344 25152
rect 17316 25100 17368 25152
rect 18052 25100 18104 25152
rect 7642 24998 7694 25050
rect 7706 24998 7758 25050
rect 7770 24998 7822 25050
rect 7834 24998 7886 25050
rect 7898 24998 7950 25050
rect 14334 24998 14386 25050
rect 14398 24998 14450 25050
rect 14462 24998 14514 25050
rect 14526 24998 14578 25050
rect 14590 24998 14642 25050
rect 21026 24998 21078 25050
rect 21090 24998 21142 25050
rect 21154 24998 21206 25050
rect 21218 24998 21270 25050
rect 21282 24998 21334 25050
rect 27718 24998 27770 25050
rect 27782 24998 27834 25050
rect 27846 24998 27898 25050
rect 27910 24998 27962 25050
rect 27974 24998 28026 25050
rect 2504 24896 2556 24948
rect 4344 24896 4396 24948
rect 5448 24939 5500 24948
rect 4712 24871 4764 24880
rect 4712 24837 4721 24871
rect 4721 24837 4755 24871
rect 4755 24837 4764 24871
rect 4712 24828 4764 24837
rect 5448 24905 5457 24939
rect 5457 24905 5491 24939
rect 5491 24905 5500 24939
rect 5448 24896 5500 24905
rect 5724 24939 5776 24948
rect 5724 24905 5733 24939
rect 5733 24905 5767 24939
rect 5767 24905 5776 24939
rect 5724 24896 5776 24905
rect 6828 24896 6880 24948
rect 8484 24896 8536 24948
rect 9772 24896 9824 24948
rect 11336 24896 11388 24948
rect 13636 24896 13688 24948
rect 15752 24896 15804 24948
rect 20720 24939 20772 24948
rect 20720 24905 20729 24939
rect 20729 24905 20763 24939
rect 20763 24905 20772 24939
rect 20720 24896 20772 24905
rect 3976 24760 4028 24812
rect 6736 24828 6788 24880
rect 8392 24828 8444 24880
rect 9496 24828 9548 24880
rect 5632 24803 5684 24812
rect 3608 24735 3660 24744
rect 3608 24701 3617 24735
rect 3617 24701 3651 24735
rect 3651 24701 3660 24735
rect 3608 24692 3660 24701
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 5816 24803 5868 24812
rect 5816 24769 5825 24803
rect 5825 24769 5859 24803
rect 5859 24769 5868 24803
rect 5816 24760 5868 24769
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 7104 24760 7156 24812
rect 8116 24760 8168 24812
rect 9588 24760 9640 24812
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 12164 24760 12216 24812
rect 12532 24760 12584 24812
rect 14924 24828 14976 24880
rect 16120 24828 16172 24880
rect 17408 24828 17460 24880
rect 17592 24871 17644 24880
rect 17592 24837 17601 24871
rect 17601 24837 17635 24871
rect 17635 24837 17644 24871
rect 17592 24828 17644 24837
rect 18604 24871 18656 24880
rect 18604 24837 18613 24871
rect 18613 24837 18647 24871
rect 18647 24837 18656 24871
rect 18604 24828 18656 24837
rect 14096 24803 14148 24812
rect 5724 24692 5776 24744
rect 4804 24624 4856 24676
rect 6276 24624 6328 24676
rect 8852 24667 8904 24676
rect 8852 24633 8861 24667
rect 8861 24633 8895 24667
rect 8895 24633 8904 24667
rect 8852 24624 8904 24633
rect 9496 24624 9548 24676
rect 5908 24556 5960 24608
rect 8300 24556 8352 24608
rect 8484 24556 8536 24608
rect 9220 24556 9272 24608
rect 14096 24769 14105 24803
rect 14105 24769 14139 24803
rect 14139 24769 14148 24803
rect 14096 24760 14148 24769
rect 15476 24692 15528 24744
rect 15568 24692 15620 24744
rect 17316 24760 17368 24812
rect 18328 24803 18380 24812
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 19708 24760 19760 24812
rect 20904 24803 20956 24812
rect 20904 24769 20913 24803
rect 20913 24769 20947 24803
rect 20947 24769 20956 24803
rect 20904 24760 20956 24769
rect 14004 24624 14056 24676
rect 11888 24556 11940 24608
rect 19340 24556 19392 24608
rect 4296 24454 4348 24506
rect 4360 24454 4412 24506
rect 4424 24454 4476 24506
rect 4488 24454 4540 24506
rect 4552 24454 4604 24506
rect 10988 24454 11040 24506
rect 11052 24454 11104 24506
rect 11116 24454 11168 24506
rect 11180 24454 11232 24506
rect 11244 24454 11296 24506
rect 17680 24454 17732 24506
rect 17744 24454 17796 24506
rect 17808 24454 17860 24506
rect 17872 24454 17924 24506
rect 17936 24454 17988 24506
rect 24372 24454 24424 24506
rect 24436 24454 24488 24506
rect 24500 24454 24552 24506
rect 24564 24454 24616 24506
rect 24628 24454 24680 24506
rect 3976 24395 4028 24404
rect 3976 24361 3985 24395
rect 3985 24361 4019 24395
rect 4019 24361 4028 24395
rect 3976 24352 4028 24361
rect 6368 24352 6420 24404
rect 9128 24352 9180 24404
rect 9496 24352 9548 24404
rect 10692 24352 10744 24404
rect 12072 24352 12124 24404
rect 14188 24352 14240 24404
rect 15108 24395 15160 24404
rect 15108 24361 15117 24395
rect 15117 24361 15151 24395
rect 15151 24361 15160 24395
rect 15108 24352 15160 24361
rect 6736 24327 6788 24336
rect 6736 24293 6745 24327
rect 6745 24293 6779 24327
rect 6779 24293 6788 24327
rect 6736 24284 6788 24293
rect 4160 24216 4212 24268
rect 5356 24259 5408 24268
rect 5356 24225 5365 24259
rect 5365 24225 5399 24259
rect 5399 24225 5408 24259
rect 5356 24216 5408 24225
rect 2228 24191 2280 24200
rect 2228 24157 2262 24191
rect 2262 24157 2280 24191
rect 2228 24148 2280 24157
rect 4712 24148 4764 24200
rect 6368 24148 6420 24200
rect 2044 24080 2096 24132
rect 3056 24080 3108 24132
rect 3608 24080 3660 24132
rect 3240 24012 3292 24064
rect 5540 24012 5592 24064
rect 5724 24080 5776 24132
rect 7380 24191 7432 24200
rect 8852 24284 8904 24336
rect 8116 24216 8168 24268
rect 11888 24259 11940 24268
rect 11888 24225 11897 24259
rect 11897 24225 11931 24259
rect 11931 24225 11940 24259
rect 11888 24216 11940 24225
rect 16580 24259 16632 24268
rect 16580 24225 16589 24259
rect 16589 24225 16623 24259
rect 16623 24225 16632 24259
rect 16580 24216 16632 24225
rect 17132 24259 17184 24268
rect 17132 24225 17141 24259
rect 17141 24225 17175 24259
rect 17175 24225 17184 24259
rect 17132 24216 17184 24225
rect 18052 24216 18104 24268
rect 20076 24216 20128 24268
rect 7380 24157 7408 24191
rect 7408 24157 7432 24191
rect 7380 24148 7432 24157
rect 8208 24123 8260 24132
rect 8208 24089 8217 24123
rect 8217 24089 8251 24123
rect 8251 24089 8260 24123
rect 8208 24080 8260 24089
rect 6736 24012 6788 24064
rect 7472 24012 7524 24064
rect 8024 24012 8076 24064
rect 10600 24148 10652 24200
rect 10876 24148 10928 24200
rect 11612 24191 11664 24200
rect 9404 24123 9456 24132
rect 9404 24089 9438 24123
rect 9438 24089 9456 24123
rect 9404 24080 9456 24089
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 15016 24148 15068 24200
rect 15108 24148 15160 24200
rect 15752 24148 15804 24200
rect 18512 24148 18564 24200
rect 19892 24148 19944 24200
rect 20904 24148 20956 24200
rect 11520 24080 11572 24132
rect 13176 24080 13228 24132
rect 19708 24123 19760 24132
rect 19708 24089 19717 24123
rect 19717 24089 19751 24123
rect 19751 24089 19760 24123
rect 19708 24080 19760 24089
rect 21456 24080 21508 24132
rect 9588 24012 9640 24064
rect 18880 24055 18932 24064
rect 18880 24021 18889 24055
rect 18889 24021 18923 24055
rect 18923 24021 18932 24055
rect 18880 24012 18932 24021
rect 7642 23910 7694 23962
rect 7706 23910 7758 23962
rect 7770 23910 7822 23962
rect 7834 23910 7886 23962
rect 7898 23910 7950 23962
rect 14334 23910 14386 23962
rect 14398 23910 14450 23962
rect 14462 23910 14514 23962
rect 14526 23910 14578 23962
rect 14590 23910 14642 23962
rect 21026 23910 21078 23962
rect 21090 23910 21142 23962
rect 21154 23910 21206 23962
rect 21218 23910 21270 23962
rect 21282 23910 21334 23962
rect 27718 23910 27770 23962
rect 27782 23910 27834 23962
rect 27846 23910 27898 23962
rect 27910 23910 27962 23962
rect 27974 23910 28026 23962
rect 1676 23851 1728 23860
rect 1676 23817 1685 23851
rect 1685 23817 1719 23851
rect 1719 23817 1728 23851
rect 1676 23808 1728 23817
rect 5632 23808 5684 23860
rect 7104 23808 7156 23860
rect 8116 23808 8168 23860
rect 8208 23808 8260 23860
rect 9220 23808 9272 23860
rect 9404 23851 9456 23860
rect 9404 23817 9413 23851
rect 9413 23817 9447 23851
rect 9447 23817 9456 23851
rect 9404 23808 9456 23817
rect 13636 23808 13688 23860
rect 8024 23740 8076 23792
rect 19892 23808 19944 23860
rect 20168 23808 20220 23860
rect 2964 23672 3016 23724
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 4712 23715 4764 23724
rect 4712 23681 4746 23715
rect 4746 23681 4764 23715
rect 4712 23672 4764 23681
rect 8300 23672 8352 23724
rect 9588 23715 9640 23724
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 3056 23647 3108 23656
rect 3056 23613 3065 23647
rect 3065 23613 3099 23647
rect 3099 23613 3108 23647
rect 3056 23604 3108 23613
rect 3332 23604 3384 23656
rect 4160 23604 4212 23656
rect 11980 23647 12032 23656
rect 11980 23613 11989 23647
rect 11989 23613 12023 23647
rect 12023 23613 12032 23647
rect 11980 23604 12032 23613
rect 6276 23536 6328 23588
rect 8484 23468 8536 23520
rect 9496 23468 9548 23520
rect 9772 23468 9824 23520
rect 12164 23536 12216 23588
rect 12256 23468 12308 23520
rect 15384 23468 15436 23520
rect 4296 23366 4348 23418
rect 4360 23366 4412 23418
rect 4424 23366 4476 23418
rect 4488 23366 4540 23418
rect 4552 23366 4604 23418
rect 10988 23366 11040 23418
rect 11052 23366 11104 23418
rect 11116 23366 11168 23418
rect 11180 23366 11232 23418
rect 11244 23366 11296 23418
rect 17680 23366 17732 23418
rect 17744 23366 17796 23418
rect 17808 23366 17860 23418
rect 17872 23366 17924 23418
rect 17936 23366 17988 23418
rect 24372 23366 24424 23418
rect 24436 23366 24488 23418
rect 24500 23366 24552 23418
rect 24564 23366 24616 23418
rect 24628 23366 24680 23418
rect 5724 23264 5776 23316
rect 8208 23264 8260 23316
rect 9496 23307 9548 23316
rect 9496 23273 9505 23307
rect 9505 23273 9539 23307
rect 9539 23273 9548 23307
rect 9496 23264 9548 23273
rect 4160 23128 4212 23180
rect 3240 23060 3292 23112
rect 3332 23103 3384 23112
rect 3332 23069 3341 23103
rect 3341 23069 3375 23103
rect 3375 23069 3384 23103
rect 3332 23060 3384 23069
rect 3884 23060 3936 23112
rect 6368 23103 6420 23112
rect 6368 23069 6377 23103
rect 6377 23069 6411 23103
rect 6411 23069 6420 23103
rect 6368 23060 6420 23069
rect 18696 23196 18748 23248
rect 11428 23128 11480 23180
rect 13176 23171 13228 23180
rect 13176 23137 13185 23171
rect 13185 23137 13219 23171
rect 13219 23137 13228 23171
rect 13176 23128 13228 23137
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 11980 23060 12032 23112
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 13636 23060 13688 23112
rect 15476 23128 15528 23180
rect 18512 23171 18564 23180
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 4620 22992 4672 23044
rect 5724 22992 5776 23044
rect 6828 22992 6880 23044
rect 9496 22992 9548 23044
rect 12624 22992 12676 23044
rect 15200 23060 15252 23112
rect 15292 23060 15344 23112
rect 17224 23060 17276 23112
rect 15016 22992 15068 23044
rect 16304 22992 16356 23044
rect 2044 22924 2096 22976
rect 8300 22924 8352 22976
rect 10048 22967 10100 22976
rect 10048 22933 10057 22967
rect 10057 22933 10091 22967
rect 10091 22933 10100 22967
rect 10048 22924 10100 22933
rect 13728 22967 13780 22976
rect 13728 22933 13737 22967
rect 13737 22933 13771 22967
rect 13771 22933 13780 22967
rect 13728 22924 13780 22933
rect 17040 22967 17092 22976
rect 17040 22933 17049 22967
rect 17049 22933 17083 22967
rect 17083 22933 17092 22967
rect 17040 22924 17092 22933
rect 18236 23060 18288 23112
rect 20168 23128 20220 23180
rect 21456 23171 21508 23180
rect 21456 23137 21465 23171
rect 21465 23137 21499 23171
rect 21499 23137 21508 23171
rect 21456 23128 21508 23137
rect 20720 22992 20772 23044
rect 18420 22924 18472 22976
rect 19248 22924 19300 22976
rect 20444 22924 20496 22976
rect 7642 22822 7694 22874
rect 7706 22822 7758 22874
rect 7770 22822 7822 22874
rect 7834 22822 7886 22874
rect 7898 22822 7950 22874
rect 14334 22822 14386 22874
rect 14398 22822 14450 22874
rect 14462 22822 14514 22874
rect 14526 22822 14578 22874
rect 14590 22822 14642 22874
rect 21026 22822 21078 22874
rect 21090 22822 21142 22874
rect 21154 22822 21206 22874
rect 21218 22822 21270 22874
rect 21282 22822 21334 22874
rect 27718 22822 27770 22874
rect 27782 22822 27834 22874
rect 27846 22822 27898 22874
rect 27910 22822 27962 22874
rect 27974 22822 28026 22874
rect 3516 22720 3568 22772
rect 8392 22720 8444 22772
rect 11152 22763 11204 22772
rect 11152 22729 11161 22763
rect 11161 22729 11195 22763
rect 11195 22729 11204 22763
rect 11152 22720 11204 22729
rect 11612 22720 11664 22772
rect 15200 22720 15252 22772
rect 10048 22695 10100 22704
rect 10048 22661 10082 22695
rect 10082 22661 10100 22695
rect 10048 22652 10100 22661
rect 12440 22652 12492 22704
rect 13728 22652 13780 22704
rect 18972 22652 19024 22704
rect 2964 22584 3016 22636
rect 4712 22584 4764 22636
rect 6368 22584 6420 22636
rect 6644 22584 6696 22636
rect 8208 22584 8260 22636
rect 12164 22584 12216 22636
rect 12716 22584 12768 22636
rect 2044 22559 2096 22568
rect 2044 22525 2053 22559
rect 2053 22525 2087 22559
rect 2087 22525 2096 22559
rect 2044 22516 2096 22525
rect 9220 22516 9272 22568
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 15292 22584 15344 22636
rect 15568 22584 15620 22636
rect 18880 22584 18932 22636
rect 20904 22720 20956 22772
rect 19248 22652 19300 22704
rect 20720 22652 20772 22704
rect 19800 22627 19852 22636
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 20168 22584 20220 22636
rect 15844 22559 15896 22568
rect 14924 22448 14976 22500
rect 15844 22525 15853 22559
rect 15853 22525 15887 22559
rect 15887 22525 15896 22559
rect 15844 22516 15896 22525
rect 16304 22559 16356 22568
rect 16304 22525 16313 22559
rect 16313 22525 16347 22559
rect 16347 22525 16356 22559
rect 16304 22516 16356 22525
rect 17224 22559 17276 22568
rect 17224 22525 17233 22559
rect 17233 22525 17267 22559
rect 17267 22525 17276 22559
rect 17224 22516 17276 22525
rect 17500 22559 17552 22568
rect 17500 22525 17509 22559
rect 17509 22525 17543 22559
rect 17543 22525 17552 22559
rect 17500 22516 17552 22525
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 19248 22516 19300 22568
rect 19432 22448 19484 22500
rect 1860 22380 1912 22432
rect 3516 22380 3568 22432
rect 13820 22380 13872 22432
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 4296 22278 4348 22330
rect 4360 22278 4412 22330
rect 4424 22278 4476 22330
rect 4488 22278 4540 22330
rect 4552 22278 4604 22330
rect 10988 22278 11040 22330
rect 11052 22278 11104 22330
rect 11116 22278 11168 22330
rect 11180 22278 11232 22330
rect 11244 22278 11296 22330
rect 17680 22278 17732 22330
rect 17744 22278 17796 22330
rect 17808 22278 17860 22330
rect 17872 22278 17924 22330
rect 17936 22278 17988 22330
rect 24372 22278 24424 22330
rect 24436 22278 24488 22330
rect 24500 22278 24552 22330
rect 24564 22278 24616 22330
rect 24628 22278 24680 22330
rect 4712 22176 4764 22228
rect 6828 22176 6880 22228
rect 11336 22176 11388 22228
rect 4620 22040 4672 22092
rect 3884 21972 3936 22024
rect 5356 21972 5408 22024
rect 8300 22015 8352 22024
rect 8300 21981 8318 22015
rect 8318 21981 8352 22015
rect 8300 21972 8352 21981
rect 9312 21972 9364 22024
rect 9220 21904 9272 21956
rect 1676 21879 1728 21888
rect 1676 21845 1685 21879
rect 1685 21845 1719 21879
rect 1719 21845 1728 21879
rect 1676 21836 1728 21845
rect 3516 21836 3568 21888
rect 6552 21836 6604 21888
rect 15200 22176 15252 22228
rect 19432 22176 19484 22228
rect 20812 22176 20864 22228
rect 13820 21972 13872 22024
rect 20352 22083 20404 22092
rect 16212 22015 16264 22024
rect 12440 21904 12492 21956
rect 13728 21904 13780 21956
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 17408 21972 17460 22024
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 20444 22015 20496 22024
rect 20444 21981 20453 22015
rect 20453 21981 20487 22015
rect 20487 21981 20496 22015
rect 20444 21972 20496 21981
rect 20904 21972 20956 22024
rect 21732 22015 21784 22024
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 22008 22015 22060 22024
rect 22008 21981 22042 22015
rect 22042 21981 22060 22015
rect 22008 21972 22060 21981
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 16304 21836 16356 21888
rect 17500 21836 17552 21888
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 19524 21879 19576 21888
rect 19524 21845 19533 21879
rect 19533 21845 19567 21879
rect 19567 21845 19576 21879
rect 19524 21836 19576 21845
rect 21364 21836 21416 21888
rect 23480 21836 23532 21888
rect 7642 21734 7694 21786
rect 7706 21734 7758 21786
rect 7770 21734 7822 21786
rect 7834 21734 7886 21786
rect 7898 21734 7950 21786
rect 14334 21734 14386 21786
rect 14398 21734 14450 21786
rect 14462 21734 14514 21786
rect 14526 21734 14578 21786
rect 14590 21734 14642 21786
rect 21026 21734 21078 21786
rect 21090 21734 21142 21786
rect 21154 21734 21206 21786
rect 21218 21734 21270 21786
rect 21282 21734 21334 21786
rect 27718 21734 27770 21786
rect 27782 21734 27834 21786
rect 27846 21734 27898 21786
rect 27910 21734 27962 21786
rect 27974 21734 28026 21786
rect 3516 21632 3568 21684
rect 3424 21564 3476 21616
rect 4620 21632 4672 21684
rect 5356 21675 5408 21684
rect 5356 21641 5365 21675
rect 5365 21641 5399 21675
rect 5399 21641 5408 21675
rect 5356 21632 5408 21641
rect 15200 21632 15252 21684
rect 15844 21632 15896 21684
rect 16212 21632 16264 21684
rect 17500 21632 17552 21684
rect 20352 21632 20404 21684
rect 22008 21632 22060 21684
rect 26332 21632 26384 21684
rect 3976 21496 4028 21548
rect 4988 21496 5040 21548
rect 5356 21539 5408 21548
rect 5356 21505 5365 21539
rect 5365 21505 5399 21539
rect 5399 21505 5408 21539
rect 5356 21496 5408 21505
rect 6552 21564 6604 21616
rect 7472 21564 7524 21616
rect 10048 21539 10100 21548
rect 10048 21505 10082 21539
rect 10082 21505 10100 21539
rect 12164 21539 12216 21548
rect 10048 21496 10100 21505
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 1492 21428 1544 21480
rect 2688 21471 2740 21480
rect 2688 21437 2697 21471
rect 2697 21437 2731 21471
rect 2731 21437 2740 21471
rect 2688 21428 2740 21437
rect 3884 21428 3936 21480
rect 6828 21471 6880 21480
rect 6828 21437 6837 21471
rect 6837 21437 6871 21471
rect 6871 21437 6880 21471
rect 6828 21428 6880 21437
rect 7380 21428 7432 21480
rect 11336 21428 11388 21480
rect 13084 21496 13136 21548
rect 16304 21564 16356 21616
rect 18696 21564 18748 21616
rect 15476 21471 15528 21480
rect 12348 21360 12400 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 8208 21292 8260 21344
rect 9220 21335 9272 21344
rect 9220 21301 9229 21335
rect 9229 21301 9263 21335
rect 9263 21301 9272 21335
rect 9220 21292 9272 21301
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 18144 21539 18196 21548
rect 18144 21505 18153 21539
rect 18153 21505 18187 21539
rect 18187 21505 18196 21539
rect 18144 21496 18196 21505
rect 19800 21496 19852 21548
rect 21272 21496 21324 21548
rect 21364 21496 21416 21548
rect 17408 21428 17460 21480
rect 14924 21360 14976 21412
rect 21916 21428 21968 21480
rect 13728 21292 13780 21344
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 18328 21335 18380 21344
rect 18328 21301 18337 21335
rect 18337 21301 18371 21335
rect 18371 21301 18380 21335
rect 18328 21292 18380 21301
rect 19064 21335 19116 21344
rect 19064 21301 19073 21335
rect 19073 21301 19107 21335
rect 19107 21301 19116 21335
rect 19064 21292 19116 21301
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 4296 21190 4348 21242
rect 4360 21190 4412 21242
rect 4424 21190 4476 21242
rect 4488 21190 4540 21242
rect 4552 21190 4604 21242
rect 10988 21190 11040 21242
rect 11052 21190 11104 21242
rect 11116 21190 11168 21242
rect 11180 21190 11232 21242
rect 11244 21190 11296 21242
rect 17680 21190 17732 21242
rect 17744 21190 17796 21242
rect 17808 21190 17860 21242
rect 17872 21190 17924 21242
rect 17936 21190 17988 21242
rect 24372 21190 24424 21242
rect 24436 21190 24488 21242
rect 24500 21190 24552 21242
rect 24564 21190 24616 21242
rect 24628 21190 24680 21242
rect 2688 21088 2740 21140
rect 6828 21088 6880 21140
rect 7472 21131 7524 21140
rect 7472 21097 7481 21131
rect 7481 21097 7515 21131
rect 7515 21097 7524 21131
rect 7472 21088 7524 21097
rect 10048 21088 10100 21140
rect 11336 21088 11388 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 1492 20952 1544 21004
rect 3884 20952 3936 21004
rect 8208 20952 8260 21004
rect 3516 20816 3568 20868
rect 4804 20884 4856 20936
rect 4988 20884 5040 20936
rect 5540 20884 5592 20936
rect 6920 20884 6972 20936
rect 7472 20884 7524 20936
rect 12164 21020 12216 21072
rect 18144 21088 18196 21140
rect 20812 21088 20864 21140
rect 21272 21088 21324 21140
rect 11428 20995 11480 21004
rect 11428 20961 11437 20995
rect 11437 20961 11471 20995
rect 11471 20961 11480 20995
rect 11428 20952 11480 20961
rect 14924 20995 14976 21004
rect 12348 20927 12400 20936
rect 6460 20816 6512 20868
rect 9220 20816 9272 20868
rect 11060 20816 11112 20868
rect 12348 20893 12357 20927
rect 12357 20893 12391 20927
rect 12391 20893 12400 20927
rect 12348 20884 12400 20893
rect 14924 20961 14933 20995
rect 14933 20961 14967 20995
rect 14967 20961 14976 20995
rect 14924 20952 14976 20961
rect 15844 20995 15896 21004
rect 15844 20961 15853 20995
rect 15853 20961 15887 20995
rect 15887 20961 15896 20995
rect 15844 20952 15896 20961
rect 18328 20995 18380 21004
rect 18328 20961 18337 20995
rect 18337 20961 18371 20995
rect 18371 20961 18380 20995
rect 18328 20952 18380 20961
rect 19064 20952 19116 21004
rect 14188 20884 14240 20936
rect 15200 20884 15252 20936
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 17040 20884 17092 20936
rect 18604 20927 18656 20936
rect 18604 20893 18613 20927
rect 18613 20893 18647 20927
rect 18647 20893 18656 20927
rect 18604 20884 18656 20893
rect 21548 20927 21600 20936
rect 17316 20816 17368 20868
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 21916 20884 21968 20936
rect 23480 20816 23532 20868
rect 2780 20748 2832 20800
rect 4712 20748 4764 20800
rect 4804 20748 4856 20800
rect 5356 20748 5408 20800
rect 7012 20748 7064 20800
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 11796 20748 11848 20800
rect 14096 20748 14148 20800
rect 16120 20791 16172 20800
rect 16120 20757 16129 20791
rect 16129 20757 16163 20791
rect 16163 20757 16172 20791
rect 16120 20748 16172 20757
rect 23664 20748 23716 20800
rect 7642 20646 7694 20698
rect 7706 20646 7758 20698
rect 7770 20646 7822 20698
rect 7834 20646 7886 20698
rect 7898 20646 7950 20698
rect 14334 20646 14386 20698
rect 14398 20646 14450 20698
rect 14462 20646 14514 20698
rect 14526 20646 14578 20698
rect 14590 20646 14642 20698
rect 21026 20646 21078 20698
rect 21090 20646 21142 20698
rect 21154 20646 21206 20698
rect 21218 20646 21270 20698
rect 21282 20646 21334 20698
rect 27718 20646 27770 20698
rect 27782 20646 27834 20698
rect 27846 20646 27898 20698
rect 27910 20646 27962 20698
rect 27974 20646 28026 20698
rect 2780 20587 2832 20596
rect 2780 20553 2789 20587
rect 2789 20553 2823 20587
rect 2823 20553 2832 20587
rect 3424 20587 3476 20596
rect 2780 20544 2832 20553
rect 3424 20553 3433 20587
rect 3433 20553 3467 20587
rect 3467 20553 3476 20587
rect 3424 20544 3476 20553
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 3240 20476 3292 20528
rect 4896 20544 4948 20596
rect 5540 20544 5592 20596
rect 6460 20544 6512 20596
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 11704 20544 11756 20596
rect 12624 20544 12676 20596
rect 4712 20476 4764 20528
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 3884 20408 3936 20460
rect 7472 20476 7524 20528
rect 5540 20340 5592 20392
rect 5356 20272 5408 20324
rect 6920 20408 6972 20460
rect 9588 20408 9640 20460
rect 4896 20204 4948 20256
rect 9680 20340 9732 20392
rect 11612 20476 11664 20528
rect 11796 20519 11848 20528
rect 11796 20485 11805 20519
rect 11805 20485 11839 20519
rect 11839 20485 11848 20519
rect 11796 20476 11848 20485
rect 14188 20544 14240 20596
rect 16028 20544 16080 20596
rect 20352 20544 20404 20596
rect 21548 20544 21600 20596
rect 23480 20587 23532 20596
rect 23480 20553 23489 20587
rect 23489 20553 23523 20587
rect 23523 20553 23532 20587
rect 23480 20544 23532 20553
rect 23664 20544 23716 20596
rect 16948 20476 17000 20528
rect 17316 20519 17368 20528
rect 17316 20485 17325 20519
rect 17325 20485 17359 20519
rect 17359 20485 17368 20519
rect 17316 20476 17368 20485
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 10416 20408 10468 20460
rect 11520 20408 11572 20460
rect 13176 20408 13228 20460
rect 13544 20408 13596 20460
rect 15568 20408 15620 20460
rect 16028 20451 16080 20460
rect 13084 20340 13136 20392
rect 14924 20383 14976 20392
rect 14924 20349 14933 20383
rect 14933 20349 14967 20383
rect 14967 20349 14976 20383
rect 14924 20340 14976 20349
rect 8484 20272 8536 20324
rect 8760 20272 8812 20324
rect 8116 20204 8168 20256
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 8852 20247 8904 20256
rect 8852 20213 8861 20247
rect 8861 20213 8895 20247
rect 8895 20213 8904 20247
rect 8852 20204 8904 20213
rect 10324 20272 10376 20324
rect 12164 20272 12216 20324
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 17592 20408 17644 20460
rect 18236 20408 18288 20460
rect 18420 20408 18472 20460
rect 18788 20408 18840 20460
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 20628 20408 20680 20460
rect 18052 20340 18104 20392
rect 19248 20340 19300 20392
rect 22100 20340 22152 20392
rect 11520 20204 11572 20256
rect 13636 20204 13688 20256
rect 18604 20272 18656 20324
rect 21732 20272 21784 20324
rect 15936 20204 15988 20256
rect 18144 20204 18196 20256
rect 18512 20204 18564 20256
rect 19064 20204 19116 20256
rect 21364 20204 21416 20256
rect 4296 20102 4348 20154
rect 4360 20102 4412 20154
rect 4424 20102 4476 20154
rect 4488 20102 4540 20154
rect 4552 20102 4604 20154
rect 10988 20102 11040 20154
rect 11052 20102 11104 20154
rect 11116 20102 11168 20154
rect 11180 20102 11232 20154
rect 11244 20102 11296 20154
rect 17680 20102 17732 20154
rect 17744 20102 17796 20154
rect 17808 20102 17860 20154
rect 17872 20102 17924 20154
rect 17936 20102 17988 20154
rect 24372 20102 24424 20154
rect 24436 20102 24488 20154
rect 24500 20102 24552 20154
rect 24564 20102 24616 20154
rect 24628 20102 24680 20154
rect 10600 20043 10652 20052
rect 10600 20009 10609 20043
rect 10609 20009 10643 20043
rect 10643 20009 10652 20043
rect 10600 20000 10652 20009
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 15568 20000 15620 20052
rect 5264 19932 5316 19984
rect 1492 19864 1544 19916
rect 7288 19864 7340 19916
rect 1860 19839 1912 19848
rect 1860 19805 1894 19839
rect 1894 19805 1912 19839
rect 1860 19796 1912 19805
rect 6920 19796 6972 19848
rect 7472 19796 7524 19848
rect 2964 19703 3016 19712
rect 2964 19669 2973 19703
rect 2973 19669 3007 19703
rect 3007 19669 3016 19703
rect 2964 19660 3016 19669
rect 3516 19660 3568 19712
rect 5908 19728 5960 19780
rect 5080 19703 5132 19712
rect 5080 19669 5089 19703
rect 5089 19669 5123 19703
rect 5123 19669 5132 19703
rect 6368 19728 6420 19780
rect 12256 19932 12308 19984
rect 11428 19864 11480 19916
rect 9956 19796 10008 19848
rect 10324 19796 10376 19848
rect 13084 19796 13136 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 13728 19796 13780 19848
rect 16028 20000 16080 20052
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 17592 20000 17644 20052
rect 18052 20000 18104 20052
rect 19800 20043 19852 20052
rect 19800 20009 19809 20043
rect 19809 20009 19843 20043
rect 19843 20009 19852 20043
rect 19800 20000 19852 20009
rect 24860 20000 24912 20052
rect 17132 19932 17184 19984
rect 5080 19660 5132 19669
rect 10140 19728 10192 19780
rect 11336 19771 11388 19780
rect 11336 19737 11345 19771
rect 11345 19737 11379 19771
rect 11379 19737 11388 19771
rect 11336 19728 11388 19737
rect 12164 19771 12216 19780
rect 12164 19737 12173 19771
rect 12173 19737 12207 19771
rect 12207 19737 12216 19771
rect 12164 19728 12216 19737
rect 13452 19728 13504 19780
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 9588 19660 9640 19712
rect 10416 19660 10468 19712
rect 10508 19660 10560 19712
rect 13268 19660 13320 19712
rect 14096 19728 14148 19780
rect 17408 19796 17460 19848
rect 19248 19864 19300 19916
rect 23664 19864 23716 19916
rect 17132 19771 17184 19780
rect 17132 19737 17141 19771
rect 17141 19737 17175 19771
rect 17175 19737 17184 19771
rect 17132 19728 17184 19737
rect 19340 19796 19392 19848
rect 20812 19796 20864 19848
rect 21456 19796 21508 19848
rect 21916 19796 21968 19848
rect 23572 19839 23624 19848
rect 23572 19805 23581 19839
rect 23581 19805 23615 19839
rect 23615 19805 23624 19839
rect 23572 19796 23624 19805
rect 25872 19796 25924 19848
rect 15200 19660 15252 19712
rect 15844 19660 15896 19712
rect 18696 19728 18748 19780
rect 20904 19728 20956 19780
rect 19340 19660 19392 19712
rect 19524 19660 19576 19712
rect 20536 19660 20588 19712
rect 20720 19660 20772 19712
rect 22284 19660 22336 19712
rect 25412 19660 25464 19712
rect 7642 19558 7694 19610
rect 7706 19558 7758 19610
rect 7770 19558 7822 19610
rect 7834 19558 7886 19610
rect 7898 19558 7950 19610
rect 14334 19558 14386 19610
rect 14398 19558 14450 19610
rect 14462 19558 14514 19610
rect 14526 19558 14578 19610
rect 14590 19558 14642 19610
rect 21026 19558 21078 19610
rect 21090 19558 21142 19610
rect 21154 19558 21206 19610
rect 21218 19558 21270 19610
rect 21282 19558 21334 19610
rect 27718 19558 27770 19610
rect 27782 19558 27834 19610
rect 27846 19558 27898 19610
rect 27910 19558 27962 19610
rect 27974 19558 28026 19610
rect 3332 19456 3384 19508
rect 4804 19456 4856 19508
rect 5908 19499 5960 19508
rect 5908 19465 5917 19499
rect 5917 19465 5951 19499
rect 5951 19465 5960 19499
rect 5908 19456 5960 19465
rect 7104 19499 7156 19508
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 8484 19456 8536 19508
rect 2964 19388 3016 19440
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 7012 19363 7064 19372
rect 7012 19329 7021 19363
rect 7021 19329 7055 19363
rect 7055 19329 7064 19363
rect 7012 19320 7064 19329
rect 7564 19388 7616 19440
rect 9956 19456 10008 19508
rect 11428 19456 11480 19508
rect 16856 19456 16908 19508
rect 18696 19456 18748 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 22284 19499 22336 19508
rect 22284 19465 22293 19499
rect 22293 19465 22327 19499
rect 22327 19465 22336 19499
rect 22284 19456 22336 19465
rect 23572 19456 23624 19508
rect 25872 19499 25924 19508
rect 25872 19465 25881 19499
rect 25881 19465 25915 19499
rect 25915 19465 25924 19499
rect 25872 19456 25924 19465
rect 10140 19388 10192 19440
rect 11520 19320 11572 19372
rect 12624 19388 12676 19440
rect 13176 19388 13228 19440
rect 15844 19431 15896 19440
rect 12072 19320 12124 19372
rect 2964 19295 3016 19304
rect 2964 19261 2973 19295
rect 2973 19261 3007 19295
rect 3007 19261 3016 19295
rect 2964 19252 3016 19261
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 7380 19252 7432 19304
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9128 19252 9180 19304
rect 11428 19252 11480 19304
rect 14188 19320 14240 19372
rect 15844 19397 15853 19431
rect 15853 19397 15887 19431
rect 15887 19397 15896 19431
rect 15844 19388 15896 19397
rect 15936 19431 15988 19440
rect 15936 19397 15945 19431
rect 15945 19397 15979 19431
rect 15979 19397 15988 19431
rect 15936 19388 15988 19397
rect 19340 19388 19392 19440
rect 20812 19388 20864 19440
rect 15384 19252 15436 19304
rect 4804 19116 4856 19168
rect 5724 19116 5776 19168
rect 6736 19116 6788 19168
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19064 19320 19116 19372
rect 20444 19363 20496 19372
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 20444 19329 20453 19363
rect 20453 19329 20487 19363
rect 20487 19329 20496 19363
rect 20444 19320 20496 19329
rect 20536 19320 20588 19372
rect 18236 19252 18288 19261
rect 20904 19320 20956 19372
rect 21640 19388 21692 19440
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 23572 19320 23624 19372
rect 25504 19320 25556 19372
rect 26332 19363 26384 19372
rect 26332 19329 26341 19363
rect 26341 19329 26375 19363
rect 26375 19329 26384 19363
rect 26332 19320 26384 19329
rect 9220 19116 9272 19168
rect 12164 19116 12216 19168
rect 16120 19116 16172 19168
rect 19248 19184 19300 19236
rect 19616 19184 19668 19236
rect 21824 19252 21876 19304
rect 22100 19295 22152 19304
rect 22100 19261 22109 19295
rect 22109 19261 22143 19295
rect 22143 19261 22152 19295
rect 22100 19252 22152 19261
rect 25412 19252 25464 19304
rect 16856 19159 16908 19168
rect 16856 19125 16865 19159
rect 16865 19125 16899 19159
rect 16899 19125 16908 19159
rect 16856 19116 16908 19125
rect 17408 19116 17460 19168
rect 18696 19116 18748 19168
rect 21548 19116 21600 19168
rect 27068 19116 27120 19168
rect 4296 19014 4348 19066
rect 4360 19014 4412 19066
rect 4424 19014 4476 19066
rect 4488 19014 4540 19066
rect 4552 19014 4604 19066
rect 10988 19014 11040 19066
rect 11052 19014 11104 19066
rect 11116 19014 11168 19066
rect 11180 19014 11232 19066
rect 11244 19014 11296 19066
rect 17680 19014 17732 19066
rect 17744 19014 17796 19066
rect 17808 19014 17860 19066
rect 17872 19014 17924 19066
rect 17936 19014 17988 19066
rect 24372 19014 24424 19066
rect 24436 19014 24488 19066
rect 24500 19014 24552 19066
rect 24564 19014 24616 19066
rect 24628 19014 24680 19066
rect 7104 18912 7156 18964
rect 10324 18912 10376 18964
rect 13084 18955 13136 18964
rect 13084 18921 13093 18955
rect 13093 18921 13127 18955
rect 13127 18921 13136 18955
rect 13084 18912 13136 18921
rect 15844 18912 15896 18964
rect 7380 18844 7432 18896
rect 7288 18776 7340 18828
rect 4160 18708 4212 18760
rect 4712 18708 4764 18760
rect 8208 18751 8260 18760
rect 6552 18640 6604 18692
rect 2228 18572 2280 18624
rect 2596 18572 2648 18624
rect 3516 18572 3568 18624
rect 7380 18615 7432 18624
rect 7380 18581 7389 18615
rect 7389 18581 7423 18615
rect 7423 18581 7432 18615
rect 7380 18572 7432 18581
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 9680 18708 9732 18760
rect 11428 18776 11480 18828
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 15108 18844 15160 18896
rect 18420 18912 18472 18964
rect 17408 18844 17460 18896
rect 20168 18912 20220 18964
rect 20812 18955 20864 18964
rect 20812 18921 20821 18955
rect 20821 18921 20855 18955
rect 20855 18921 20864 18955
rect 20812 18912 20864 18921
rect 9588 18640 9640 18692
rect 11336 18640 11388 18692
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 14004 18708 14056 18760
rect 14924 18776 14976 18828
rect 11796 18640 11848 18692
rect 12624 18640 12676 18692
rect 16856 18708 16908 18760
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 25504 18776 25556 18828
rect 16396 18640 16448 18692
rect 17500 18708 17552 18760
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 12164 18572 12216 18624
rect 13636 18615 13688 18624
rect 13636 18581 13645 18615
rect 13645 18581 13679 18615
rect 13679 18581 13688 18615
rect 13636 18572 13688 18581
rect 18420 18572 18472 18624
rect 22836 18640 22888 18692
rect 22100 18572 22152 18624
rect 23480 18708 23532 18760
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 25320 18708 25372 18760
rect 26608 18708 26660 18760
rect 25780 18640 25832 18692
rect 27344 18640 27396 18692
rect 7642 18470 7694 18522
rect 7706 18470 7758 18522
rect 7770 18470 7822 18522
rect 7834 18470 7886 18522
rect 7898 18470 7950 18522
rect 14334 18470 14386 18522
rect 14398 18470 14450 18522
rect 14462 18470 14514 18522
rect 14526 18470 14578 18522
rect 14590 18470 14642 18522
rect 21026 18470 21078 18522
rect 21090 18470 21142 18522
rect 21154 18470 21206 18522
rect 21218 18470 21270 18522
rect 21282 18470 21334 18522
rect 27718 18470 27770 18522
rect 27782 18470 27834 18522
rect 27846 18470 27898 18522
rect 27910 18470 27962 18522
rect 27974 18470 28026 18522
rect 6368 18368 6420 18420
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 9588 18368 9640 18420
rect 9680 18368 9732 18420
rect 10416 18368 10468 18420
rect 13728 18368 13780 18420
rect 2596 18300 2648 18352
rect 5724 18343 5776 18352
rect 5724 18309 5733 18343
rect 5733 18309 5767 18343
rect 5767 18309 5776 18343
rect 5724 18300 5776 18309
rect 7380 18300 7432 18352
rect 8300 18300 8352 18352
rect 9220 18300 9272 18352
rect 14188 18368 14240 18420
rect 20628 18368 20680 18420
rect 20904 18368 20956 18420
rect 23572 18411 23624 18420
rect 23572 18377 23581 18411
rect 23581 18377 23615 18411
rect 23615 18377 23624 18411
rect 23572 18368 23624 18377
rect 16396 18300 16448 18352
rect 19340 18300 19392 18352
rect 22836 18343 22888 18352
rect 22836 18309 22845 18343
rect 22845 18309 22879 18343
rect 22879 18309 22888 18343
rect 22836 18300 22888 18309
rect 1952 18028 2004 18080
rect 3332 18275 3384 18284
rect 3332 18241 3341 18275
rect 3341 18241 3375 18275
rect 3375 18241 3384 18275
rect 3332 18232 3384 18241
rect 4620 18232 4672 18284
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 13636 18232 13688 18284
rect 15936 18232 15988 18284
rect 3976 18164 4028 18216
rect 6000 18207 6052 18216
rect 6000 18173 6009 18207
rect 6009 18173 6043 18207
rect 6043 18173 6052 18207
rect 6000 18164 6052 18173
rect 8024 18164 8076 18216
rect 8668 18164 8720 18216
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 12532 18164 12584 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 15200 18164 15252 18216
rect 17500 18232 17552 18284
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 21916 18232 21968 18284
rect 22376 18232 22428 18284
rect 25320 18232 25372 18284
rect 17592 18164 17644 18216
rect 26516 18207 26568 18216
rect 26516 18173 26525 18207
rect 26525 18173 26559 18207
rect 26559 18173 26568 18207
rect 26516 18164 26568 18173
rect 13820 18096 13872 18148
rect 26240 18096 26292 18148
rect 9496 18028 9548 18080
rect 9772 18028 9824 18080
rect 14740 18028 14792 18080
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 17040 18028 17092 18080
rect 20904 18028 20956 18080
rect 4296 17926 4348 17978
rect 4360 17926 4412 17978
rect 4424 17926 4476 17978
rect 4488 17926 4540 17978
rect 4552 17926 4604 17978
rect 10988 17926 11040 17978
rect 11052 17926 11104 17978
rect 11116 17926 11168 17978
rect 11180 17926 11232 17978
rect 11244 17926 11296 17978
rect 17680 17926 17732 17978
rect 17744 17926 17796 17978
rect 17808 17926 17860 17978
rect 17872 17926 17924 17978
rect 17936 17926 17988 17978
rect 24372 17926 24424 17978
rect 24436 17926 24488 17978
rect 24500 17926 24552 17978
rect 24564 17926 24616 17978
rect 24628 17926 24680 17978
rect 2964 17824 3016 17876
rect 3976 17824 4028 17876
rect 5540 17824 5592 17876
rect 8300 17824 8352 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 11796 17824 11848 17876
rect 13084 17824 13136 17876
rect 15384 17867 15436 17876
rect 9404 17756 9456 17808
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 9496 17731 9548 17740
rect 9496 17697 9505 17731
rect 9505 17697 9539 17731
rect 9539 17697 9548 17731
rect 9496 17688 9548 17697
rect 3056 17620 3108 17672
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 6920 17620 6972 17672
rect 7472 17620 7524 17672
rect 8852 17620 8904 17672
rect 9680 17620 9732 17672
rect 4068 17484 4120 17536
rect 9956 17688 10008 17740
rect 10508 17663 10560 17672
rect 10508 17629 10517 17663
rect 10517 17629 10551 17663
rect 10551 17629 10560 17663
rect 10508 17620 10560 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 11704 17552 11756 17604
rect 12716 17756 12768 17808
rect 13268 17688 13320 17740
rect 12808 17620 12860 17672
rect 12716 17552 12768 17604
rect 13452 17595 13504 17604
rect 13452 17561 13461 17595
rect 13461 17561 13495 17595
rect 13495 17561 13504 17595
rect 13452 17552 13504 17561
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 8852 17484 8904 17536
rect 10876 17484 10928 17536
rect 12348 17484 12400 17536
rect 14004 17620 14056 17672
rect 15384 17833 15393 17867
rect 15393 17833 15427 17867
rect 15427 17833 15436 17867
rect 15384 17824 15436 17833
rect 13728 17552 13780 17604
rect 14096 17484 14148 17536
rect 14924 17552 14976 17604
rect 16948 17688 17000 17740
rect 19616 17824 19668 17876
rect 21824 17824 21876 17876
rect 17684 17756 17736 17808
rect 18236 17688 18288 17740
rect 20812 17688 20864 17740
rect 22284 17756 22336 17808
rect 22468 17731 22520 17740
rect 22468 17697 22477 17731
rect 22477 17697 22511 17731
rect 22511 17697 22520 17731
rect 22468 17688 22520 17697
rect 20628 17663 20680 17672
rect 17592 17552 17644 17604
rect 17040 17484 17092 17536
rect 17500 17484 17552 17536
rect 18144 17527 18196 17536
rect 18144 17493 18153 17527
rect 18153 17493 18187 17527
rect 18187 17493 18196 17527
rect 18144 17484 18196 17493
rect 20628 17629 20637 17663
rect 20637 17629 20671 17663
rect 20671 17629 20680 17663
rect 20628 17620 20680 17629
rect 22100 17663 22152 17672
rect 22100 17629 22109 17663
rect 22109 17629 22143 17663
rect 22143 17629 22152 17663
rect 22100 17620 22152 17629
rect 22284 17620 22336 17672
rect 23572 17620 23624 17672
rect 23756 17620 23808 17672
rect 24584 17620 24636 17672
rect 20812 17552 20864 17604
rect 19708 17484 19760 17536
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 20536 17527 20588 17536
rect 20536 17493 20545 17527
rect 20545 17493 20579 17527
rect 20579 17493 20588 17527
rect 20536 17484 20588 17493
rect 22008 17484 22060 17536
rect 22928 17527 22980 17536
rect 22928 17493 22937 17527
rect 22937 17493 22971 17527
rect 22971 17493 22980 17527
rect 22928 17484 22980 17493
rect 23940 17484 23992 17536
rect 24216 17484 24268 17536
rect 27068 17731 27120 17740
rect 27068 17697 27077 17731
rect 27077 17697 27111 17731
rect 27111 17697 27120 17731
rect 27068 17688 27120 17697
rect 27344 17731 27396 17740
rect 27344 17697 27353 17731
rect 27353 17697 27387 17731
rect 27387 17697 27396 17731
rect 27344 17688 27396 17697
rect 26516 17552 26568 17604
rect 26332 17484 26384 17536
rect 7642 17382 7694 17434
rect 7706 17382 7758 17434
rect 7770 17382 7822 17434
rect 7834 17382 7886 17434
rect 7898 17382 7950 17434
rect 14334 17382 14386 17434
rect 14398 17382 14450 17434
rect 14462 17382 14514 17434
rect 14526 17382 14578 17434
rect 14590 17382 14642 17434
rect 21026 17382 21078 17434
rect 21090 17382 21142 17434
rect 21154 17382 21206 17434
rect 21218 17382 21270 17434
rect 21282 17382 21334 17434
rect 27718 17382 27770 17434
rect 27782 17382 27834 17434
rect 27846 17382 27898 17434
rect 27910 17382 27962 17434
rect 27974 17382 28026 17434
rect 2228 17280 2280 17332
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 6644 17280 6696 17332
rect 5080 17212 5132 17264
rect 10048 17280 10100 17332
rect 10784 17280 10836 17332
rect 10692 17212 10744 17264
rect 11428 17212 11480 17264
rect 1584 17187 1636 17196
rect 1584 17153 1593 17187
rect 1593 17153 1627 17187
rect 1627 17153 1636 17187
rect 1584 17144 1636 17153
rect 3516 17144 3568 17196
rect 4160 17144 4212 17196
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 6736 17144 6788 17196
rect 8944 17144 8996 17196
rect 9404 17144 9456 17196
rect 10600 17144 10652 17196
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 9956 17119 10008 17128
rect 9956 17085 9965 17119
rect 9965 17085 9999 17119
rect 9999 17085 10008 17119
rect 9956 17076 10008 17085
rect 13728 17280 13780 17332
rect 15200 17280 15252 17332
rect 12900 17212 12952 17264
rect 13084 17212 13136 17264
rect 13452 17212 13504 17264
rect 14556 17144 14608 17196
rect 18144 17212 18196 17264
rect 15200 17144 15252 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 1768 17051 1820 17060
rect 1768 17017 1777 17051
rect 1777 17017 1811 17051
rect 1811 17017 1820 17051
rect 1768 17008 1820 17017
rect 4160 17008 4212 17060
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 8300 17008 8352 17060
rect 10508 17008 10560 17060
rect 13820 17076 13872 17128
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 17316 17076 17368 17128
rect 19340 17255 19392 17264
rect 19340 17221 19349 17255
rect 19349 17221 19383 17255
rect 19383 17221 19392 17255
rect 19340 17212 19392 17221
rect 24584 17280 24636 17332
rect 19984 17212 20036 17264
rect 18788 17119 18840 17128
rect 18788 17085 18797 17119
rect 18797 17085 18831 17119
rect 18831 17085 18840 17119
rect 18788 17076 18840 17085
rect 19156 17076 19208 17128
rect 20168 17187 20220 17196
rect 20168 17153 20178 17187
rect 20178 17153 20212 17187
rect 20212 17153 20220 17187
rect 20168 17144 20220 17153
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 20536 17187 20588 17196
rect 22192 17212 22244 17264
rect 24216 17255 24268 17264
rect 24216 17221 24225 17255
rect 24225 17221 24259 17255
rect 24259 17221 24268 17255
rect 24216 17212 24268 17221
rect 20536 17153 20550 17187
rect 20550 17153 20584 17187
rect 20584 17153 20588 17187
rect 20536 17144 20588 17153
rect 22376 17144 22428 17196
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 22100 17076 22152 17128
rect 23296 17119 23348 17128
rect 7196 16940 7248 16992
rect 8852 16983 8904 16992
rect 8852 16949 8861 16983
rect 8861 16949 8895 16983
rect 8895 16949 8904 16983
rect 8852 16940 8904 16949
rect 9496 16940 9548 16992
rect 13912 17008 13964 17060
rect 11704 16940 11756 16992
rect 14648 16940 14700 16992
rect 21088 17008 21140 17060
rect 17408 16940 17460 16992
rect 21916 17008 21968 17060
rect 23296 17085 23305 17119
rect 23305 17085 23339 17119
rect 23339 17085 23348 17119
rect 23296 17076 23348 17085
rect 25412 17076 25464 17128
rect 21364 16983 21416 16992
rect 21364 16949 21373 16983
rect 21373 16949 21407 16983
rect 21407 16949 21416 16983
rect 21364 16940 21416 16949
rect 26332 16983 26384 16992
rect 26332 16949 26341 16983
rect 26341 16949 26375 16983
rect 26375 16949 26384 16983
rect 26332 16940 26384 16949
rect 4296 16838 4348 16890
rect 4360 16838 4412 16890
rect 4424 16838 4476 16890
rect 4488 16838 4540 16890
rect 4552 16838 4604 16890
rect 10988 16838 11040 16890
rect 11052 16838 11104 16890
rect 11116 16838 11168 16890
rect 11180 16838 11232 16890
rect 11244 16838 11296 16890
rect 17680 16838 17732 16890
rect 17744 16838 17796 16890
rect 17808 16838 17860 16890
rect 17872 16838 17924 16890
rect 17936 16838 17988 16890
rect 24372 16838 24424 16890
rect 24436 16838 24488 16890
rect 24500 16838 24552 16890
rect 24564 16838 24616 16890
rect 24628 16838 24680 16890
rect 4068 16736 4120 16788
rect 6000 16736 6052 16788
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 7196 16736 7248 16788
rect 8760 16736 8812 16788
rect 8852 16736 8904 16788
rect 10600 16736 10652 16788
rect 13268 16736 13320 16788
rect 14556 16736 14608 16788
rect 14648 16736 14700 16788
rect 7932 16668 7984 16720
rect 14832 16668 14884 16720
rect 18788 16736 18840 16788
rect 19616 16736 19668 16788
rect 21916 16736 21968 16788
rect 5080 16600 5132 16652
rect 6920 16600 6972 16652
rect 8944 16600 8996 16652
rect 9680 16600 9732 16652
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10692 16600 10744 16652
rect 17592 16643 17644 16652
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 20904 16668 20956 16720
rect 22468 16736 22520 16788
rect 23480 16643 23532 16652
rect 23480 16609 23489 16643
rect 23489 16609 23523 16643
rect 23523 16609 23532 16643
rect 23480 16600 23532 16609
rect 24676 16600 24728 16652
rect 26240 16600 26292 16652
rect 27160 16600 27212 16652
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 3792 16532 3844 16584
rect 3884 16532 3936 16584
rect 4804 16532 4856 16584
rect 6644 16575 6696 16584
rect 6644 16541 6653 16575
rect 6653 16541 6687 16575
rect 6687 16541 6696 16575
rect 6644 16532 6696 16541
rect 9496 16532 9548 16584
rect 10048 16532 10100 16584
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 15016 16532 15068 16584
rect 18696 16532 18748 16584
rect 19156 16532 19208 16584
rect 19616 16575 19668 16584
rect 19616 16541 19625 16575
rect 19625 16541 19659 16575
rect 19659 16541 19668 16575
rect 19616 16532 19668 16541
rect 20536 16532 20588 16584
rect 20720 16532 20772 16584
rect 21088 16532 21140 16584
rect 8116 16464 8168 16516
rect 11336 16464 11388 16516
rect 2044 16439 2096 16448
rect 2044 16405 2053 16439
rect 2053 16405 2087 16439
rect 2087 16405 2096 16439
rect 2044 16396 2096 16405
rect 2780 16439 2832 16448
rect 2780 16405 2789 16439
rect 2789 16405 2823 16439
rect 2823 16405 2832 16439
rect 2780 16396 2832 16405
rect 6000 16396 6052 16448
rect 8024 16396 8076 16448
rect 10784 16396 10836 16448
rect 10968 16396 11020 16448
rect 15384 16507 15436 16516
rect 11796 16396 11848 16448
rect 13452 16396 13504 16448
rect 13636 16396 13688 16448
rect 15384 16473 15393 16507
rect 15393 16473 15427 16507
rect 15427 16473 15436 16507
rect 15384 16464 15436 16473
rect 19708 16464 19760 16516
rect 25320 16532 25372 16584
rect 25596 16532 25648 16584
rect 22192 16464 22244 16516
rect 23388 16507 23440 16516
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 15660 16396 15712 16448
rect 22376 16396 22428 16448
rect 23388 16473 23397 16507
rect 23397 16473 23431 16507
rect 23431 16473 23440 16507
rect 23388 16464 23440 16473
rect 23572 16464 23624 16516
rect 23940 16464 23992 16516
rect 25504 16464 25556 16516
rect 26976 16507 27028 16516
rect 26976 16473 26985 16507
rect 26985 16473 27019 16507
rect 27019 16473 27028 16507
rect 26976 16464 27028 16473
rect 7642 16294 7694 16346
rect 7706 16294 7758 16346
rect 7770 16294 7822 16346
rect 7834 16294 7886 16346
rect 7898 16294 7950 16346
rect 14334 16294 14386 16346
rect 14398 16294 14450 16346
rect 14462 16294 14514 16346
rect 14526 16294 14578 16346
rect 14590 16294 14642 16346
rect 21026 16294 21078 16346
rect 21090 16294 21142 16346
rect 21154 16294 21206 16346
rect 21218 16294 21270 16346
rect 21282 16294 21334 16346
rect 27718 16294 27770 16346
rect 27782 16294 27834 16346
rect 27846 16294 27898 16346
rect 27910 16294 27962 16346
rect 27974 16294 28026 16346
rect 2228 16192 2280 16244
rect 3792 16192 3844 16244
rect 2044 16124 2096 16176
rect 3700 16124 3752 16176
rect 5724 16124 5776 16176
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 10600 16192 10652 16244
rect 10968 16192 11020 16244
rect 12808 16192 12860 16244
rect 15936 16235 15988 16244
rect 15936 16201 15945 16235
rect 15945 16201 15979 16235
rect 15979 16201 15988 16235
rect 15936 16192 15988 16201
rect 17316 16235 17368 16244
rect 17316 16201 17325 16235
rect 17325 16201 17359 16235
rect 17359 16201 17368 16235
rect 17316 16192 17368 16201
rect 17408 16235 17460 16244
rect 17408 16201 17417 16235
rect 17417 16201 17451 16235
rect 17451 16201 17460 16235
rect 18696 16235 18748 16244
rect 17408 16192 17460 16201
rect 18696 16201 18705 16235
rect 18705 16201 18739 16235
rect 18739 16201 18748 16235
rect 18696 16192 18748 16201
rect 10692 16124 10744 16176
rect 14188 16124 14240 16176
rect 14740 16124 14792 16176
rect 15752 16124 15804 16176
rect 20812 16192 20864 16244
rect 22284 16192 22336 16244
rect 27160 16235 27212 16244
rect 19524 16124 19576 16176
rect 22376 16124 22428 16176
rect 23296 16124 23348 16176
rect 27160 16201 27169 16235
rect 27169 16201 27203 16235
rect 27203 16201 27212 16235
rect 27160 16192 27212 16201
rect 6000 16056 6052 16065
rect 8024 16099 8076 16108
rect 2780 15988 2832 16040
rect 8024 16065 8033 16099
rect 8033 16065 8067 16099
rect 8067 16065 8076 16099
rect 8024 16056 8076 16065
rect 8760 16056 8812 16108
rect 10968 16056 11020 16108
rect 21640 16056 21692 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 8300 15988 8352 16040
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 10508 15988 10560 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 17224 16031 17276 16040
rect 17224 15997 17233 16031
rect 17233 15997 17267 16031
rect 17267 15997 17276 16031
rect 17224 15988 17276 15997
rect 20812 16031 20864 16040
rect 10048 15920 10100 15972
rect 9036 15852 9088 15904
rect 10508 15895 10560 15904
rect 10508 15861 10517 15895
rect 10517 15861 10551 15895
rect 10551 15861 10560 15895
rect 10508 15852 10560 15861
rect 10784 15920 10836 15972
rect 13544 15920 13596 15972
rect 17408 15920 17460 15972
rect 20812 15997 20821 16031
rect 20821 15997 20855 16031
rect 20855 15997 20864 16031
rect 20812 15988 20864 15997
rect 19616 15852 19668 15904
rect 20904 15920 20956 15972
rect 22008 15920 22060 15972
rect 23480 15920 23532 15972
rect 23940 15920 23992 15972
rect 23296 15852 23348 15904
rect 25596 15852 25648 15904
rect 4296 15750 4348 15802
rect 4360 15750 4412 15802
rect 4424 15750 4476 15802
rect 4488 15750 4540 15802
rect 4552 15750 4604 15802
rect 10988 15750 11040 15802
rect 11052 15750 11104 15802
rect 11116 15750 11168 15802
rect 11180 15750 11232 15802
rect 11244 15750 11296 15802
rect 17680 15750 17732 15802
rect 17744 15750 17796 15802
rect 17808 15750 17860 15802
rect 17872 15750 17924 15802
rect 17936 15750 17988 15802
rect 24372 15750 24424 15802
rect 24436 15750 24488 15802
rect 24500 15750 24552 15802
rect 24564 15750 24616 15802
rect 24628 15750 24680 15802
rect 4160 15691 4212 15700
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 4160 15648 4212 15657
rect 8300 15648 8352 15700
rect 8852 15648 8904 15700
rect 6828 15580 6880 15632
rect 12532 15648 12584 15700
rect 10692 15555 10744 15564
rect 10692 15521 10701 15555
rect 10701 15521 10735 15555
rect 10735 15521 10744 15555
rect 10692 15512 10744 15521
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 4160 15444 4212 15496
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 7104 15444 7156 15496
rect 9220 15444 9272 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 10784 15444 10836 15496
rect 12624 15580 12676 15632
rect 15384 15648 15436 15700
rect 16856 15648 16908 15700
rect 19708 15648 19760 15700
rect 20812 15648 20864 15700
rect 3332 15376 3384 15428
rect 4068 15419 4120 15428
rect 4068 15385 4077 15419
rect 4077 15385 4111 15419
rect 4111 15385 4120 15419
rect 4068 15376 4120 15385
rect 5816 15419 5868 15428
rect 5816 15385 5825 15419
rect 5825 15385 5859 15419
rect 5859 15385 5868 15419
rect 5816 15376 5868 15385
rect 11888 15444 11940 15496
rect 17592 15512 17644 15564
rect 23388 15648 23440 15700
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 22100 15580 22152 15632
rect 23388 15555 23440 15564
rect 23388 15521 23397 15555
rect 23397 15521 23431 15555
rect 23431 15521 23440 15555
rect 23388 15512 23440 15521
rect 26332 15648 26384 15700
rect 25780 15555 25832 15564
rect 2872 15308 2924 15360
rect 3424 15351 3476 15360
rect 3424 15317 3433 15351
rect 3433 15317 3467 15351
rect 3467 15317 3476 15351
rect 3424 15308 3476 15317
rect 11428 15376 11480 15428
rect 11796 15376 11848 15428
rect 13452 15376 13504 15428
rect 14832 15444 14884 15496
rect 15660 15487 15712 15496
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 8300 15308 8352 15360
rect 9680 15308 9732 15360
rect 14096 15376 14148 15428
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 17500 15444 17552 15496
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 21364 15444 21416 15496
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 23480 15444 23532 15496
rect 25780 15521 25789 15555
rect 25789 15521 25823 15555
rect 25823 15521 25832 15555
rect 25780 15512 25832 15521
rect 26976 15512 27028 15564
rect 24860 15487 24912 15496
rect 24860 15453 24869 15487
rect 24869 15453 24903 15487
rect 24903 15453 24912 15487
rect 24860 15444 24912 15453
rect 25044 15419 25096 15428
rect 16396 15308 16448 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 22928 15308 22980 15360
rect 25044 15385 25053 15419
rect 25053 15385 25087 15419
rect 25087 15385 25096 15419
rect 25044 15376 25096 15385
rect 26608 15308 26660 15360
rect 7642 15206 7694 15258
rect 7706 15206 7758 15258
rect 7770 15206 7822 15258
rect 7834 15206 7886 15258
rect 7898 15206 7950 15258
rect 14334 15206 14386 15258
rect 14398 15206 14450 15258
rect 14462 15206 14514 15258
rect 14526 15206 14578 15258
rect 14590 15206 14642 15258
rect 21026 15206 21078 15258
rect 21090 15206 21142 15258
rect 21154 15206 21206 15258
rect 21218 15206 21270 15258
rect 21282 15206 21334 15258
rect 27718 15206 27770 15258
rect 27782 15206 27834 15258
rect 27846 15206 27898 15258
rect 27910 15206 27962 15258
rect 27974 15206 28026 15258
rect 3700 15147 3752 15156
rect 3700 15113 3709 15147
rect 3709 15113 3743 15147
rect 3743 15113 3752 15147
rect 3700 15104 3752 15113
rect 5816 15104 5868 15156
rect 8208 15104 8260 15156
rect 10692 15104 10744 15156
rect 10784 15104 10836 15156
rect 1676 15036 1728 15088
rect 2872 15079 2924 15088
rect 2872 15045 2881 15079
rect 2881 15045 2915 15079
rect 2915 15045 2924 15079
rect 2872 15036 2924 15045
rect 4160 15036 4212 15088
rect 4988 15036 5040 15088
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 2780 14968 2832 15020
rect 3424 14968 3476 15020
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 9036 14968 9088 15020
rect 9680 15036 9732 15088
rect 10784 14968 10836 15020
rect 10876 14968 10928 15020
rect 4160 14900 4212 14952
rect 6828 14900 6880 14952
rect 8668 14900 8720 14952
rect 12164 14943 12216 14952
rect 5816 14832 5868 14884
rect 7104 14832 7156 14884
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 7472 14764 7524 14816
rect 9036 14764 9088 14816
rect 12164 14909 12173 14943
rect 12173 14909 12207 14943
rect 12207 14909 12216 14943
rect 12164 14900 12216 14909
rect 15200 15104 15252 15156
rect 15660 15036 15712 15088
rect 13544 14968 13596 15020
rect 17132 15104 17184 15156
rect 17316 15104 17368 15156
rect 20168 15104 20220 15156
rect 17592 15036 17644 15088
rect 19432 15036 19484 15088
rect 19524 15079 19576 15088
rect 19524 15045 19533 15079
rect 19533 15045 19567 15079
rect 19567 15045 19576 15079
rect 22468 15079 22520 15088
rect 19524 15036 19576 15045
rect 22468 15045 22477 15079
rect 22477 15045 22511 15079
rect 22511 15045 22520 15079
rect 22468 15036 22520 15045
rect 15660 14900 15712 14952
rect 10416 14764 10468 14816
rect 11612 14764 11664 14816
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 16396 14900 16448 14952
rect 19340 15011 19392 15020
rect 19340 14977 19349 15011
rect 19349 14977 19383 15011
rect 19383 14977 19392 15011
rect 19340 14968 19392 14977
rect 21456 14968 21508 15020
rect 22652 14968 22704 15020
rect 23480 14968 23532 15020
rect 23756 14968 23808 15020
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 20904 14900 20956 14952
rect 23204 14900 23256 14952
rect 26424 15104 26476 15156
rect 27160 15147 27212 15156
rect 27160 15113 27169 15147
rect 27169 15113 27203 15147
rect 27203 15113 27212 15147
rect 27160 15104 27212 15113
rect 25320 14968 25372 15020
rect 25596 14968 25648 15020
rect 24860 14900 24912 14952
rect 26608 14900 26660 14952
rect 16856 14807 16908 14816
rect 11704 14764 11756 14773
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 17224 14764 17276 14816
rect 25044 14832 25096 14884
rect 21456 14764 21508 14816
rect 4296 14662 4348 14714
rect 4360 14662 4412 14714
rect 4424 14662 4476 14714
rect 4488 14662 4540 14714
rect 4552 14662 4604 14714
rect 10988 14662 11040 14714
rect 11052 14662 11104 14714
rect 11116 14662 11168 14714
rect 11180 14662 11232 14714
rect 11244 14662 11296 14714
rect 17680 14662 17732 14714
rect 17744 14662 17796 14714
rect 17808 14662 17860 14714
rect 17872 14662 17924 14714
rect 17936 14662 17988 14714
rect 24372 14662 24424 14714
rect 24436 14662 24488 14714
rect 24500 14662 24552 14714
rect 24564 14662 24616 14714
rect 24628 14662 24680 14714
rect 4160 14560 4212 14612
rect 4988 14603 5040 14612
rect 4988 14569 4997 14603
rect 4997 14569 5031 14603
rect 5031 14569 5040 14603
rect 4988 14560 5040 14569
rect 5540 14560 5592 14612
rect 1676 14424 1728 14476
rect 8300 14424 8352 14476
rect 1860 14288 1912 14340
rect 3056 14288 3108 14340
rect 2136 14220 2188 14272
rect 2228 14220 2280 14272
rect 3976 14356 4028 14408
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 8024 14288 8076 14340
rect 11704 14560 11756 14612
rect 12348 14560 12400 14612
rect 9496 14356 9548 14408
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 11612 14424 11664 14476
rect 10416 14356 10468 14408
rect 10508 14288 10560 14340
rect 10600 14288 10652 14340
rect 12072 14288 12124 14340
rect 12992 14288 13044 14340
rect 13544 14560 13596 14612
rect 14004 14560 14056 14612
rect 17592 14603 17644 14612
rect 17592 14569 17601 14603
rect 17601 14569 17635 14603
rect 17635 14569 17644 14603
rect 17592 14560 17644 14569
rect 20352 14560 20404 14612
rect 22468 14603 22520 14612
rect 13452 14424 13504 14476
rect 13636 14356 13688 14408
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 15752 14288 15804 14340
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 18972 14492 19024 14544
rect 22468 14569 22477 14603
rect 22477 14569 22511 14603
rect 22511 14569 22520 14603
rect 22468 14560 22520 14569
rect 22652 14560 22704 14612
rect 16304 14356 16356 14408
rect 16856 14356 16908 14408
rect 19340 14356 19392 14408
rect 19524 14356 19576 14408
rect 19800 14288 19852 14340
rect 22652 14424 22704 14476
rect 20904 14356 20956 14408
rect 23296 14399 23348 14408
rect 23296 14365 23305 14399
rect 23305 14365 23339 14399
rect 23339 14365 23348 14399
rect 23296 14356 23348 14365
rect 25044 14356 25096 14408
rect 25320 14399 25372 14408
rect 25320 14365 25329 14399
rect 25329 14365 25363 14399
rect 25363 14365 25372 14399
rect 25320 14356 25372 14365
rect 25596 14356 25648 14408
rect 26424 14356 26476 14408
rect 27068 14356 27120 14408
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 7564 14220 7616 14272
rect 10048 14220 10100 14272
rect 12164 14220 12216 14272
rect 13084 14263 13136 14272
rect 13084 14229 13093 14263
rect 13093 14229 13127 14263
rect 13127 14229 13136 14263
rect 13084 14220 13136 14229
rect 15660 14220 15712 14272
rect 19064 14220 19116 14272
rect 21364 14331 21416 14340
rect 21364 14297 21398 14331
rect 21398 14297 21416 14331
rect 26332 14331 26384 14340
rect 21364 14288 21416 14297
rect 26332 14297 26341 14331
rect 26341 14297 26375 14331
rect 26375 14297 26384 14331
rect 26332 14288 26384 14297
rect 26792 14331 26844 14340
rect 26792 14297 26801 14331
rect 26801 14297 26835 14331
rect 26835 14297 26844 14331
rect 26792 14288 26844 14297
rect 23204 14263 23256 14272
rect 23204 14229 23213 14263
rect 23213 14229 23247 14263
rect 23247 14229 23256 14263
rect 23204 14220 23256 14229
rect 24032 14220 24084 14272
rect 7642 14118 7694 14170
rect 7706 14118 7758 14170
rect 7770 14118 7822 14170
rect 7834 14118 7886 14170
rect 7898 14118 7950 14170
rect 14334 14118 14386 14170
rect 14398 14118 14450 14170
rect 14462 14118 14514 14170
rect 14526 14118 14578 14170
rect 14590 14118 14642 14170
rect 21026 14118 21078 14170
rect 21090 14118 21142 14170
rect 21154 14118 21206 14170
rect 21218 14118 21270 14170
rect 21282 14118 21334 14170
rect 27718 14118 27770 14170
rect 27782 14118 27834 14170
rect 27846 14118 27898 14170
rect 27910 14118 27962 14170
rect 27974 14118 28026 14170
rect 1768 14016 1820 14068
rect 2228 14059 2280 14068
rect 2228 14025 2237 14059
rect 2237 14025 2271 14059
rect 2271 14025 2280 14059
rect 2228 14016 2280 14025
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 3332 14016 3384 14068
rect 7288 14016 7340 14068
rect 7564 14016 7616 14068
rect 9128 14016 9180 14068
rect 9496 14016 9548 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 13452 14016 13504 14068
rect 14280 14016 14332 14068
rect 2136 13948 2188 14000
rect 2504 13948 2556 14000
rect 2780 13880 2832 13932
rect 1768 13744 1820 13796
rect 4896 13880 4948 13932
rect 7380 13948 7432 14000
rect 9036 13948 9088 14000
rect 6368 13880 6420 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10600 13880 10652 13932
rect 4160 13812 4212 13864
rect 6736 13812 6788 13864
rect 9956 13855 10008 13864
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 10876 13812 10928 13864
rect 11428 13880 11480 13932
rect 12072 13923 12124 13932
rect 12072 13889 12081 13923
rect 12081 13889 12115 13923
rect 12115 13889 12124 13923
rect 12072 13880 12124 13889
rect 12348 13880 12400 13932
rect 12808 13880 12860 13932
rect 12900 13880 12952 13932
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 5356 13744 5408 13796
rect 6276 13676 6328 13728
rect 11520 13744 11572 13796
rect 11980 13744 12032 13796
rect 13820 13812 13872 13864
rect 14004 13812 14056 13864
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 19340 14016 19392 14068
rect 18972 13948 19024 14000
rect 15752 13880 15804 13932
rect 17592 13880 17644 13932
rect 20904 14016 20956 14068
rect 25044 14016 25096 14068
rect 27160 14059 27212 14068
rect 27160 14025 27169 14059
rect 27169 14025 27203 14059
rect 27203 14025 27212 14059
rect 27160 14016 27212 14025
rect 26332 13948 26384 14000
rect 19616 13923 19668 13932
rect 19616 13889 19650 13923
rect 19650 13889 19668 13923
rect 19616 13880 19668 13889
rect 21916 13880 21968 13932
rect 23480 13880 23532 13932
rect 14096 13744 14148 13796
rect 14648 13744 14700 13796
rect 15108 13744 15160 13796
rect 17316 13812 17368 13864
rect 20904 13812 20956 13864
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 25136 13812 25188 13864
rect 17408 13744 17460 13796
rect 9128 13676 9180 13728
rect 12164 13676 12216 13728
rect 12440 13676 12492 13728
rect 12624 13676 12676 13728
rect 12992 13676 13044 13728
rect 15292 13676 15344 13728
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 23388 13719 23440 13728
rect 23388 13685 23397 13719
rect 23397 13685 23431 13719
rect 23431 13685 23440 13719
rect 23388 13676 23440 13685
rect 24768 13676 24820 13728
rect 4296 13574 4348 13626
rect 4360 13574 4412 13626
rect 4424 13574 4476 13626
rect 4488 13574 4540 13626
rect 4552 13574 4604 13626
rect 10988 13574 11040 13626
rect 11052 13574 11104 13626
rect 11116 13574 11168 13626
rect 11180 13574 11232 13626
rect 11244 13574 11296 13626
rect 17680 13574 17732 13626
rect 17744 13574 17796 13626
rect 17808 13574 17860 13626
rect 17872 13574 17924 13626
rect 17936 13574 17988 13626
rect 24372 13574 24424 13626
rect 24436 13574 24488 13626
rect 24500 13574 24552 13626
rect 24564 13574 24616 13626
rect 24628 13574 24680 13626
rect 5540 13472 5592 13524
rect 8300 13472 8352 13524
rect 8576 13472 8628 13524
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 9864 13472 9916 13524
rect 12440 13472 12492 13524
rect 12624 13472 12676 13524
rect 12716 13472 12768 13524
rect 15200 13472 15252 13524
rect 15292 13472 15344 13524
rect 13728 13447 13780 13456
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 7288 13336 7340 13388
rect 1952 13311 2004 13320
rect 1952 13277 1961 13311
rect 1961 13277 1995 13311
rect 1995 13277 2004 13311
rect 1952 13268 2004 13277
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2780 13200 2832 13252
rect 4712 13268 4764 13320
rect 5264 13268 5316 13320
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 8300 13311 8352 13320
rect 5540 13268 5592 13277
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 10508 13379 10560 13388
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 12072 13336 12124 13388
rect 13728 13413 13737 13447
rect 13737 13413 13771 13447
rect 13771 13413 13780 13447
rect 13728 13404 13780 13413
rect 14096 13404 14148 13456
rect 17224 13472 17276 13524
rect 18328 13472 18380 13524
rect 13912 13336 13964 13388
rect 12164 13268 12216 13320
rect 6552 13200 6604 13252
rect 6736 13200 6788 13252
rect 9404 13200 9456 13252
rect 14188 13268 14240 13320
rect 15200 13336 15252 13388
rect 17316 13336 17368 13388
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 17408 13311 17460 13320
rect 2228 13132 2280 13184
rect 4160 13132 4212 13184
rect 5356 13132 5408 13184
rect 7564 13132 7616 13184
rect 8024 13132 8076 13184
rect 13084 13200 13136 13252
rect 13452 13200 13504 13252
rect 13544 13200 13596 13252
rect 14280 13200 14332 13252
rect 15292 13200 15344 13252
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 23204 13472 23256 13524
rect 24768 13515 24820 13524
rect 24768 13481 24777 13515
rect 24777 13481 24811 13515
rect 24811 13481 24820 13515
rect 24768 13472 24820 13481
rect 27068 13515 27120 13524
rect 27068 13481 27077 13515
rect 27077 13481 27111 13515
rect 27111 13481 27120 13515
rect 27068 13472 27120 13481
rect 23664 13404 23716 13456
rect 19984 13336 20036 13388
rect 20076 13379 20128 13388
rect 20076 13345 20085 13379
rect 20085 13345 20119 13379
rect 20119 13345 20128 13379
rect 20720 13379 20772 13388
rect 20076 13336 20128 13345
rect 20720 13345 20729 13379
rect 20729 13345 20763 13379
rect 20763 13345 20772 13379
rect 20720 13336 20772 13345
rect 22008 13379 22060 13388
rect 22008 13345 22017 13379
rect 22017 13345 22051 13379
rect 22051 13345 22060 13379
rect 22008 13336 22060 13345
rect 18880 13311 18932 13320
rect 17500 13243 17552 13252
rect 10232 13132 10284 13184
rect 11704 13132 11756 13184
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 11980 13132 12032 13184
rect 14188 13132 14240 13184
rect 14648 13132 14700 13184
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 17500 13209 17509 13243
rect 17509 13209 17543 13243
rect 17543 13209 17552 13243
rect 17500 13200 17552 13209
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 19432 13268 19484 13320
rect 24032 13311 24084 13320
rect 19524 13200 19576 13252
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 26792 13336 26844 13388
rect 25136 13268 25188 13320
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 18512 13132 18564 13184
rect 19340 13132 19392 13184
rect 20076 13132 20128 13184
rect 22652 13132 22704 13184
rect 26608 13200 26660 13252
rect 7642 13030 7694 13082
rect 7706 13030 7758 13082
rect 7770 13030 7822 13082
rect 7834 13030 7886 13082
rect 7898 13030 7950 13082
rect 14334 13030 14386 13082
rect 14398 13030 14450 13082
rect 14462 13030 14514 13082
rect 14526 13030 14578 13082
rect 14590 13030 14642 13082
rect 21026 13030 21078 13082
rect 21090 13030 21142 13082
rect 21154 13030 21206 13082
rect 21218 13030 21270 13082
rect 21282 13030 21334 13082
rect 27718 13030 27770 13082
rect 27782 13030 27834 13082
rect 27846 13030 27898 13082
rect 27910 13030 27962 13082
rect 27974 13030 28026 13082
rect 1860 12928 1912 12980
rect 1952 12928 2004 12980
rect 2780 12860 2832 12912
rect 4252 12928 4304 12980
rect 4712 12928 4764 12980
rect 6644 12928 6696 12980
rect 7104 12928 7156 12980
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 10508 12928 10560 12980
rect 11520 12928 11572 12980
rect 13544 12928 13596 12980
rect 14004 12928 14056 12980
rect 16948 12928 17000 12980
rect 17132 12928 17184 12980
rect 17316 12928 17368 12980
rect 19616 12928 19668 12980
rect 19984 12928 20036 12980
rect 21364 12928 21416 12980
rect 21916 12928 21968 12980
rect 23388 12928 23440 12980
rect 25320 12928 25372 12980
rect 4160 12860 4212 12912
rect 5264 12860 5316 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 4712 12792 4764 12844
rect 7288 12792 7340 12844
rect 7656 12724 7708 12776
rect 6920 12656 6972 12708
rect 10232 12792 10284 12844
rect 9312 12724 9364 12776
rect 9680 12724 9732 12776
rect 12440 12792 12492 12844
rect 12532 12792 12584 12844
rect 13176 12792 13228 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 12716 12724 12768 12776
rect 13452 12724 13504 12776
rect 14188 12860 14240 12912
rect 15016 12860 15068 12912
rect 15844 12860 15896 12912
rect 17408 12860 17460 12912
rect 18144 12860 18196 12912
rect 18512 12903 18564 12912
rect 18512 12869 18521 12903
rect 18521 12869 18555 12903
rect 18555 12869 18564 12903
rect 18512 12860 18564 12869
rect 19708 12860 19760 12912
rect 23296 12903 23348 12912
rect 13728 12792 13780 12844
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 18696 12835 18748 12844
rect 18696 12801 18741 12835
rect 18741 12801 18748 12835
rect 18696 12792 18748 12801
rect 19340 12835 19392 12844
rect 19340 12801 19349 12835
rect 19349 12801 19383 12835
rect 19383 12801 19392 12835
rect 19340 12792 19392 12801
rect 19800 12792 19852 12844
rect 20444 12792 20496 12844
rect 23296 12869 23305 12903
rect 23305 12869 23339 12903
rect 23339 12869 23348 12903
rect 23296 12860 23348 12869
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 22100 12792 22152 12844
rect 23388 12792 23440 12844
rect 25136 12792 25188 12844
rect 22468 12724 22520 12776
rect 22652 12767 22704 12776
rect 22652 12733 22661 12767
rect 22661 12733 22695 12767
rect 22695 12733 22704 12767
rect 22652 12724 22704 12733
rect 19064 12656 19116 12708
rect 6000 12631 6052 12640
rect 6000 12597 6009 12631
rect 6009 12597 6043 12631
rect 6043 12597 6052 12631
rect 6000 12588 6052 12597
rect 9772 12588 9824 12640
rect 10232 12588 10284 12640
rect 10876 12588 10928 12640
rect 12348 12588 12400 12640
rect 12440 12588 12492 12640
rect 12992 12588 13044 12640
rect 16672 12588 16724 12640
rect 17316 12588 17368 12640
rect 18880 12588 18932 12640
rect 18972 12588 19024 12640
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 23388 12588 23440 12640
rect 4296 12486 4348 12538
rect 4360 12486 4412 12538
rect 4424 12486 4476 12538
rect 4488 12486 4540 12538
rect 4552 12486 4604 12538
rect 10988 12486 11040 12538
rect 11052 12486 11104 12538
rect 11116 12486 11168 12538
rect 11180 12486 11232 12538
rect 11244 12486 11296 12538
rect 17680 12486 17732 12538
rect 17744 12486 17796 12538
rect 17808 12486 17860 12538
rect 17872 12486 17924 12538
rect 17936 12486 17988 12538
rect 24372 12486 24424 12538
rect 24436 12486 24488 12538
rect 24500 12486 24552 12538
rect 24564 12486 24616 12538
rect 24628 12486 24680 12538
rect 5172 12316 5224 12368
rect 6920 12384 6972 12436
rect 7104 12384 7156 12436
rect 8208 12384 8260 12436
rect 8392 12384 8444 12436
rect 9956 12384 10008 12436
rect 9128 12316 9180 12368
rect 10600 12316 10652 12368
rect 4620 12291 4672 12300
rect 2780 12180 2832 12232
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 6920 12248 6972 12300
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 8116 12248 8168 12300
rect 1584 12112 1636 12164
rect 2044 12112 2096 12164
rect 4712 12180 4764 12232
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 11336 12248 11388 12300
rect 11612 12248 11664 12300
rect 5448 12155 5500 12164
rect 5448 12121 5482 12155
rect 5482 12121 5500 12155
rect 5448 12112 5500 12121
rect 6000 12112 6052 12164
rect 6644 12112 6696 12164
rect 6920 12112 6972 12164
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4436 12087 4488 12096
rect 4436 12053 4445 12087
rect 4445 12053 4479 12087
rect 4479 12053 4488 12087
rect 4436 12044 4488 12053
rect 4896 12044 4948 12096
rect 8300 12112 8352 12164
rect 8576 12155 8628 12164
rect 7472 12044 7524 12096
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 9036 12112 9088 12164
rect 10692 12180 10744 12232
rect 13820 12316 13872 12368
rect 16764 12384 16816 12436
rect 17316 12384 17368 12436
rect 19064 12384 19116 12436
rect 22468 12384 22520 12436
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 13912 12180 13964 12232
rect 15936 12180 15988 12232
rect 18512 12248 18564 12300
rect 18972 12248 19024 12300
rect 9404 12155 9456 12164
rect 9404 12121 9413 12155
rect 9413 12121 9447 12155
rect 9447 12121 9456 12155
rect 9404 12112 9456 12121
rect 10416 12112 10468 12164
rect 11796 12112 11848 12164
rect 12624 12112 12676 12164
rect 18880 12180 18932 12232
rect 19524 12180 19576 12232
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 21732 12223 21784 12232
rect 16120 12155 16172 12164
rect 16120 12121 16154 12155
rect 16154 12121 16172 12155
rect 16120 12112 16172 12121
rect 17132 12112 17184 12164
rect 19340 12112 19392 12164
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 10784 12044 10836 12096
rect 11704 12044 11756 12096
rect 12532 12044 12584 12096
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13636 12044 13688 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 18972 12044 19024 12096
rect 20444 12044 20496 12096
rect 21916 12087 21968 12096
rect 21916 12053 21925 12087
rect 21925 12053 21959 12087
rect 21959 12053 21968 12087
rect 21916 12044 21968 12053
rect 7642 11942 7694 11994
rect 7706 11942 7758 11994
rect 7770 11942 7822 11994
rect 7834 11942 7886 11994
rect 7898 11942 7950 11994
rect 14334 11942 14386 11994
rect 14398 11942 14450 11994
rect 14462 11942 14514 11994
rect 14526 11942 14578 11994
rect 14590 11942 14642 11994
rect 21026 11942 21078 11994
rect 21090 11942 21142 11994
rect 21154 11942 21206 11994
rect 21218 11942 21270 11994
rect 21282 11942 21334 11994
rect 27718 11942 27770 11994
rect 27782 11942 27834 11994
rect 27846 11942 27898 11994
rect 27910 11942 27962 11994
rect 27974 11942 28026 11994
rect 4436 11840 4488 11892
rect 4620 11772 4672 11824
rect 3976 11704 4028 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 4988 11679 5040 11688
rect 4988 11645 4997 11679
rect 4997 11645 5031 11679
rect 5031 11645 5040 11679
rect 4988 11636 5040 11645
rect 5448 11772 5500 11824
rect 7932 11840 7984 11892
rect 10416 11883 10468 11892
rect 6368 11704 6420 11756
rect 6460 11704 6512 11756
rect 2872 11500 2924 11552
rect 4712 11568 4764 11620
rect 4160 11500 4212 11552
rect 6552 11636 6604 11688
rect 7012 11772 7064 11824
rect 7472 11772 7524 11824
rect 7840 11772 7892 11824
rect 8852 11815 8904 11824
rect 8852 11781 8861 11815
rect 8861 11781 8895 11815
rect 8895 11781 8904 11815
rect 8852 11772 8904 11781
rect 9956 11772 10008 11824
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 11796 11840 11848 11892
rect 15016 11840 15068 11892
rect 15200 11883 15252 11892
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 16120 11840 16172 11892
rect 18972 11883 19024 11892
rect 18972 11849 18981 11883
rect 18981 11849 19015 11883
rect 19015 11849 19024 11883
rect 18972 11840 19024 11849
rect 10692 11772 10744 11824
rect 7564 11636 7616 11688
rect 10232 11704 10284 11756
rect 10600 11704 10652 11756
rect 10876 11704 10928 11756
rect 12440 11772 12492 11824
rect 14924 11772 14976 11824
rect 17592 11772 17644 11824
rect 19708 11840 19760 11892
rect 20168 11840 20220 11892
rect 20444 11840 20496 11892
rect 22744 11840 22796 11892
rect 21916 11772 21968 11824
rect 11980 11747 12032 11756
rect 11980 11713 12014 11747
rect 12014 11713 12032 11747
rect 11980 11704 12032 11713
rect 12348 11704 12400 11756
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 16028 11704 16080 11756
rect 16672 11704 16724 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 17316 11704 17368 11756
rect 17684 11704 17736 11756
rect 8300 11636 8352 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 11520 11636 11572 11688
rect 14004 11636 14056 11688
rect 15292 11636 15344 11688
rect 17500 11636 17552 11688
rect 18788 11704 18840 11756
rect 22560 11704 22612 11756
rect 23204 11704 23256 11756
rect 26332 11704 26384 11756
rect 11612 11568 11664 11620
rect 9220 11500 9272 11552
rect 19708 11568 19760 11620
rect 20444 11568 20496 11620
rect 20628 11500 20680 11552
rect 22192 11500 22244 11552
rect 23112 11500 23164 11552
rect 24860 11500 24912 11552
rect 4296 11398 4348 11450
rect 4360 11398 4412 11450
rect 4424 11398 4476 11450
rect 4488 11398 4540 11450
rect 4552 11398 4604 11450
rect 10988 11398 11040 11450
rect 11052 11398 11104 11450
rect 11116 11398 11168 11450
rect 11180 11398 11232 11450
rect 11244 11398 11296 11450
rect 17680 11398 17732 11450
rect 17744 11398 17796 11450
rect 17808 11398 17860 11450
rect 17872 11398 17924 11450
rect 17936 11398 17988 11450
rect 24372 11398 24424 11450
rect 24436 11398 24488 11450
rect 24500 11398 24552 11450
rect 24564 11398 24616 11450
rect 24628 11398 24680 11450
rect 4988 11296 5040 11348
rect 5172 11296 5224 11348
rect 4620 11160 4672 11212
rect 4804 11228 4856 11280
rect 6368 11228 6420 11280
rect 2872 11092 2924 11144
rect 5080 11092 5132 11144
rect 2136 11024 2188 11076
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 6828 11092 6880 11144
rect 6552 11024 6604 11076
rect 7748 11296 7800 11348
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 17592 11296 17644 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19340 11296 19392 11348
rect 20628 11296 20680 11348
rect 21732 11339 21784 11348
rect 21732 11305 21741 11339
rect 21741 11305 21775 11339
rect 21775 11305 21784 11339
rect 21732 11296 21784 11305
rect 22744 11296 22796 11348
rect 23296 11296 23348 11348
rect 26332 11339 26384 11348
rect 26332 11305 26341 11339
rect 26341 11305 26375 11339
rect 26375 11305 26384 11339
rect 26332 11296 26384 11305
rect 7380 11228 7432 11280
rect 9220 11271 9272 11280
rect 9220 11237 9229 11271
rect 9229 11237 9263 11271
rect 9263 11237 9272 11271
rect 9220 11228 9272 11237
rect 9496 11228 9548 11280
rect 8392 11160 8444 11212
rect 10140 11160 10192 11212
rect 8576 11092 8628 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 8484 11024 8536 11076
rect 9496 11092 9548 11144
rect 10324 11092 10376 11144
rect 16672 11135 16724 11144
rect 7012 10956 7064 11008
rect 11336 10999 11388 11008
rect 11336 10965 11345 10999
rect 11345 10965 11379 10999
rect 11379 10965 11388 10999
rect 11336 10956 11388 10965
rect 12440 10956 12492 11008
rect 12716 11024 12768 11076
rect 13636 10999 13688 11008
rect 13636 10965 13645 10999
rect 13645 10965 13679 10999
rect 13679 10965 13688 10999
rect 13636 10956 13688 10965
rect 14096 10956 14148 11008
rect 14832 10956 14884 11008
rect 15936 11024 15988 11076
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18972 11160 19024 11212
rect 20720 11203 20772 11212
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 22192 11203 22244 11212
rect 20720 11160 20772 11169
rect 22192 11169 22201 11203
rect 22201 11169 22235 11203
rect 22235 11169 22244 11203
rect 22192 11160 22244 11169
rect 23112 11160 23164 11212
rect 24860 11203 24912 11212
rect 24860 11169 24869 11203
rect 24869 11169 24903 11203
rect 24903 11169 24912 11203
rect 24860 11160 24912 11169
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 17316 11024 17368 11076
rect 20168 11092 20220 11144
rect 22100 11092 22152 11144
rect 19616 11024 19668 11076
rect 20444 11024 20496 11076
rect 19800 10956 19852 11008
rect 21364 10956 21416 11008
rect 23296 11024 23348 11076
rect 24768 11024 24820 11076
rect 24952 11024 25004 11076
rect 7642 10854 7694 10906
rect 7706 10854 7758 10906
rect 7770 10854 7822 10906
rect 7834 10854 7886 10906
rect 7898 10854 7950 10906
rect 14334 10854 14386 10906
rect 14398 10854 14450 10906
rect 14462 10854 14514 10906
rect 14526 10854 14578 10906
rect 14590 10854 14642 10906
rect 21026 10854 21078 10906
rect 21090 10854 21142 10906
rect 21154 10854 21206 10906
rect 21218 10854 21270 10906
rect 21282 10854 21334 10906
rect 27718 10854 27770 10906
rect 27782 10854 27834 10906
rect 27846 10854 27898 10906
rect 27910 10854 27962 10906
rect 27974 10854 28026 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 9680 10752 9732 10804
rect 11980 10752 12032 10804
rect 12440 10752 12492 10804
rect 13912 10795 13964 10804
rect 13912 10761 13921 10795
rect 13921 10761 13955 10795
rect 13955 10761 13964 10795
rect 13912 10752 13964 10761
rect 16672 10752 16724 10804
rect 4804 10684 4856 10736
rect 4160 10616 4212 10668
rect 6920 10684 6972 10736
rect 10324 10684 10376 10736
rect 11336 10684 11388 10736
rect 14096 10684 14148 10736
rect 19616 10684 19668 10736
rect 20536 10752 20588 10804
rect 24952 10795 25004 10804
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 8116 10616 8168 10668
rect 4988 10548 5040 10600
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 9772 10616 9824 10668
rect 9680 10548 9732 10600
rect 10048 10616 10100 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 12532 10659 12584 10668
rect 12532 10625 12541 10659
rect 12541 10625 12575 10659
rect 12575 10625 12584 10659
rect 12532 10616 12584 10625
rect 10140 10591 10192 10600
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 8208 10480 8260 10532
rect 9772 10480 9824 10532
rect 12164 10548 12216 10600
rect 14832 10616 14884 10668
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 17316 10659 17368 10668
rect 15476 10616 15528 10625
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 21364 10616 21416 10668
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 25320 10684 25372 10736
rect 25136 10616 25188 10668
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 17500 10591 17552 10600
rect 17500 10557 17509 10591
rect 17509 10557 17543 10591
rect 17543 10557 17552 10591
rect 17500 10548 17552 10557
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 2872 10412 2924 10464
rect 4252 10412 4304 10464
rect 4620 10412 4672 10464
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 7656 10412 7708 10464
rect 10048 10412 10100 10464
rect 14096 10480 14148 10532
rect 15200 10480 15252 10532
rect 15936 10480 15988 10532
rect 16764 10480 16816 10532
rect 11336 10412 11388 10464
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 19432 10412 19484 10464
rect 20996 10412 21048 10464
rect 23296 10412 23348 10464
rect 4296 10310 4348 10362
rect 4360 10310 4412 10362
rect 4424 10310 4476 10362
rect 4488 10310 4540 10362
rect 4552 10310 4604 10362
rect 10988 10310 11040 10362
rect 11052 10310 11104 10362
rect 11116 10310 11168 10362
rect 11180 10310 11232 10362
rect 11244 10310 11296 10362
rect 17680 10310 17732 10362
rect 17744 10310 17796 10362
rect 17808 10310 17860 10362
rect 17872 10310 17924 10362
rect 17936 10310 17988 10362
rect 24372 10310 24424 10362
rect 24436 10310 24488 10362
rect 24500 10310 24552 10362
rect 24564 10310 24616 10362
rect 24628 10310 24680 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 5540 10208 5592 10260
rect 9128 10208 9180 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 12808 10208 12860 10260
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 18328 10208 18380 10260
rect 19524 10208 19576 10260
rect 20260 10208 20312 10260
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 11520 10140 11572 10192
rect 4712 10072 4764 10124
rect 5540 10072 5592 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 13636 10140 13688 10192
rect 22100 10183 22152 10192
rect 22100 10149 22109 10183
rect 22109 10149 22143 10183
rect 22143 10149 22152 10183
rect 22100 10140 22152 10149
rect 14832 10115 14884 10124
rect 14832 10081 14841 10115
rect 14841 10081 14875 10115
rect 14875 10081 14884 10115
rect 14832 10072 14884 10081
rect 15292 10072 15344 10124
rect 17316 10072 17368 10124
rect 18512 10072 18564 10124
rect 23112 10115 23164 10124
rect 23112 10081 23121 10115
rect 23121 10081 23155 10115
rect 23155 10081 23164 10115
rect 23112 10072 23164 10081
rect 2136 10004 2188 10056
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 6552 10004 6604 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 9864 10047 9916 10056
rect 7380 9979 7432 9988
rect 7380 9945 7389 9979
rect 7389 9945 7423 9979
rect 7423 9945 7432 9979
rect 7380 9936 7432 9945
rect 8392 9979 8444 9988
rect 8392 9945 8401 9979
rect 8401 9945 8435 9979
rect 8435 9945 8444 9979
rect 8392 9936 8444 9945
rect 8484 9936 8536 9988
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 13084 10004 13136 10056
rect 15384 10004 15436 10056
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 17500 10004 17552 10056
rect 19524 10004 19576 10056
rect 19800 10047 19852 10056
rect 19800 10013 19809 10047
rect 19809 10013 19843 10047
rect 19843 10013 19852 10047
rect 19800 10004 19852 10013
rect 20996 10047 21048 10056
rect 20996 10013 21030 10047
rect 21030 10013 21048 10047
rect 10692 9979 10744 9988
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 2504 9868 2556 9877
rect 2964 9868 3016 9920
rect 4160 9868 4212 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 10232 9911 10284 9920
rect 6920 9868 6972 9877
rect 10232 9877 10241 9911
rect 10241 9877 10275 9911
rect 10275 9877 10284 9911
rect 10232 9868 10284 9877
rect 10692 9945 10701 9979
rect 10701 9945 10735 9979
rect 10735 9945 10744 9979
rect 10692 9936 10744 9945
rect 14188 9936 14240 9988
rect 14832 9936 14884 9988
rect 16580 9936 16632 9988
rect 13268 9868 13320 9920
rect 15844 9911 15896 9920
rect 15844 9877 15853 9911
rect 15853 9877 15887 9911
rect 15887 9877 15896 9911
rect 15844 9868 15896 9877
rect 16120 9868 16172 9920
rect 19248 9936 19300 9988
rect 20996 10004 21048 10013
rect 23756 10047 23808 10056
rect 23756 10013 23765 10047
rect 23765 10013 23799 10047
rect 23799 10013 23808 10047
rect 23756 10004 23808 10013
rect 20812 9936 20864 9988
rect 22008 9936 22060 9988
rect 23388 9936 23440 9988
rect 25228 9936 25280 9988
rect 18420 9868 18472 9920
rect 20536 9868 20588 9920
rect 22928 9911 22980 9920
rect 22928 9877 22937 9911
rect 22937 9877 22971 9911
rect 22971 9877 22980 9911
rect 22928 9868 22980 9877
rect 23296 9868 23348 9920
rect 7642 9766 7694 9818
rect 7706 9766 7758 9818
rect 7770 9766 7822 9818
rect 7834 9766 7886 9818
rect 7898 9766 7950 9818
rect 14334 9766 14386 9818
rect 14398 9766 14450 9818
rect 14462 9766 14514 9818
rect 14526 9766 14578 9818
rect 14590 9766 14642 9818
rect 21026 9766 21078 9818
rect 21090 9766 21142 9818
rect 21154 9766 21206 9818
rect 21218 9766 21270 9818
rect 21282 9766 21334 9818
rect 27718 9766 27770 9818
rect 27782 9766 27834 9818
rect 27846 9766 27898 9818
rect 27910 9766 27962 9818
rect 27974 9766 28026 9818
rect 4528 9664 4580 9716
rect 10048 9664 10100 9716
rect 10140 9664 10192 9716
rect 11428 9664 11480 9716
rect 12716 9664 12768 9716
rect 15844 9664 15896 9716
rect 16304 9707 16356 9716
rect 16304 9673 16313 9707
rect 16313 9673 16347 9707
rect 16347 9673 16356 9707
rect 16304 9664 16356 9673
rect 20536 9707 20588 9716
rect 20536 9673 20545 9707
rect 20545 9673 20579 9707
rect 20579 9673 20588 9707
rect 20536 9664 20588 9673
rect 2504 9596 2556 9648
rect 3884 9596 3936 9648
rect 4160 9639 4212 9648
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 4160 9605 4169 9639
rect 4169 9605 4203 9639
rect 4203 9605 4212 9639
rect 4160 9596 4212 9605
rect 6552 9639 6604 9648
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 6552 9605 6561 9639
rect 6561 9605 6595 9639
rect 6595 9605 6604 9639
rect 6552 9596 6604 9605
rect 8392 9596 8444 9648
rect 13820 9596 13872 9648
rect 15476 9596 15528 9648
rect 17500 9596 17552 9648
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 7012 9528 7064 9537
rect 7196 9528 7248 9580
rect 4620 9460 4672 9512
rect 4528 9392 4580 9444
rect 7472 9392 7524 9444
rect 8760 9528 8812 9580
rect 10232 9528 10284 9580
rect 10692 9460 10744 9512
rect 8484 9392 8536 9444
rect 13728 9571 13780 9580
rect 13728 9537 13737 9571
rect 13737 9537 13771 9571
rect 13771 9537 13780 9571
rect 13728 9528 13780 9537
rect 15016 9528 15068 9580
rect 15936 9528 15988 9580
rect 12716 9392 12768 9444
rect 14832 9460 14884 9512
rect 3608 9324 3660 9376
rect 10140 9324 10192 9376
rect 10784 9324 10836 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 14556 9324 14608 9376
rect 17592 9528 17644 9580
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 18328 9503 18380 9512
rect 17408 9460 17460 9469
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 23020 9596 23072 9648
rect 24768 9596 24820 9648
rect 25228 9639 25280 9648
rect 25228 9605 25237 9639
rect 25237 9605 25271 9639
rect 25271 9605 25280 9639
rect 25228 9596 25280 9605
rect 19248 9528 19300 9580
rect 19432 9571 19484 9580
rect 19432 9537 19466 9571
rect 19466 9537 19484 9571
rect 19432 9528 19484 9537
rect 19800 9528 19852 9580
rect 22652 9528 22704 9580
rect 23204 9571 23256 9580
rect 23204 9537 23213 9571
rect 23213 9537 23247 9571
rect 23247 9537 23256 9571
rect 23204 9528 23256 9537
rect 20536 9460 20588 9512
rect 25504 9503 25556 9512
rect 25504 9469 25513 9503
rect 25513 9469 25547 9503
rect 25547 9469 25556 9503
rect 25504 9460 25556 9469
rect 18052 9392 18104 9444
rect 18880 9324 18932 9376
rect 22836 9392 22888 9444
rect 20720 9324 20772 9376
rect 21088 9324 21140 9376
rect 23572 9324 23624 9376
rect 23756 9367 23808 9376
rect 23756 9333 23765 9367
rect 23765 9333 23799 9367
rect 23799 9333 23808 9367
rect 23756 9324 23808 9333
rect 4296 9222 4348 9274
rect 4360 9222 4412 9274
rect 4424 9222 4476 9274
rect 4488 9222 4540 9274
rect 4552 9222 4604 9274
rect 10988 9222 11040 9274
rect 11052 9222 11104 9274
rect 11116 9222 11168 9274
rect 11180 9222 11232 9274
rect 11244 9222 11296 9274
rect 17680 9222 17732 9274
rect 17744 9222 17796 9274
rect 17808 9222 17860 9274
rect 17872 9222 17924 9274
rect 17936 9222 17988 9274
rect 24372 9222 24424 9274
rect 24436 9222 24488 9274
rect 24500 9222 24552 9274
rect 24564 9222 24616 9274
rect 24628 9222 24680 9274
rect 2044 9120 2096 9172
rect 5172 9120 5224 9172
rect 3148 8984 3200 9036
rect 4988 9052 5040 9104
rect 7288 9120 7340 9172
rect 7380 9120 7432 9172
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 2688 8848 2740 8900
rect 5816 8891 5868 8900
rect 5816 8857 5825 8891
rect 5825 8857 5859 8891
rect 5859 8857 5868 8891
rect 5816 8848 5868 8857
rect 6552 8848 6604 8900
rect 9772 9120 9824 9172
rect 12808 9120 12860 9172
rect 13268 9120 13320 9172
rect 16948 9120 17000 9172
rect 17316 9120 17368 9172
rect 17592 9163 17644 9172
rect 17592 9129 17601 9163
rect 17601 9129 17635 9163
rect 17635 9129 17644 9163
rect 17592 9120 17644 9129
rect 18144 9120 18196 9172
rect 21088 9120 21140 9172
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 11796 8984 11848 9036
rect 11888 8984 11940 9036
rect 15200 9027 15252 9036
rect 8760 8916 8812 8968
rect 10140 8848 10192 8900
rect 10968 8848 11020 8900
rect 11428 8916 11480 8968
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 15200 8993 15209 9027
rect 15209 8993 15243 9027
rect 15243 8993 15252 9027
rect 15200 8984 15252 8993
rect 16304 8984 16356 9036
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 17224 8959 17276 8968
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17224 8916 17276 8925
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18880 8959 18932 8968
rect 18696 8916 18748 8925
rect 18880 8925 18889 8959
rect 18889 8925 18923 8959
rect 18923 8925 18932 8959
rect 18880 8916 18932 8925
rect 20812 9027 20864 9036
rect 20812 8993 20821 9027
rect 20821 8993 20855 9027
rect 20855 8993 20864 9027
rect 20812 8984 20864 8993
rect 11520 8848 11572 8900
rect 4620 8780 4672 8832
rect 6828 8780 6880 8832
rect 13820 8780 13872 8832
rect 19432 8823 19484 8832
rect 19432 8789 19441 8823
rect 19441 8789 19475 8823
rect 19475 8789 19484 8823
rect 19432 8780 19484 8789
rect 20720 8916 20772 8968
rect 24952 9052 25004 9104
rect 22100 8984 22152 9036
rect 24768 8984 24820 9036
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 23204 8959 23256 8968
rect 22008 8916 22060 8925
rect 23204 8925 23213 8959
rect 23213 8925 23247 8959
rect 23247 8925 23256 8959
rect 23204 8916 23256 8925
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 25136 8916 25188 8925
rect 25320 8959 25372 8968
rect 25320 8925 25329 8959
rect 25329 8925 25363 8959
rect 25363 8925 25372 8959
rect 26148 8959 26200 8968
rect 25320 8916 25372 8925
rect 26148 8925 26157 8959
rect 26157 8925 26191 8959
rect 26191 8925 26200 8959
rect 26148 8916 26200 8925
rect 22284 8780 22336 8832
rect 7642 8678 7694 8730
rect 7706 8678 7758 8730
rect 7770 8678 7822 8730
rect 7834 8678 7886 8730
rect 7898 8678 7950 8730
rect 14334 8678 14386 8730
rect 14398 8678 14450 8730
rect 14462 8678 14514 8730
rect 14526 8678 14578 8730
rect 14590 8678 14642 8730
rect 21026 8678 21078 8730
rect 21090 8678 21142 8730
rect 21154 8678 21206 8730
rect 21218 8678 21270 8730
rect 21282 8678 21334 8730
rect 27718 8678 27770 8730
rect 27782 8678 27834 8730
rect 27846 8678 27898 8730
rect 27910 8678 27962 8730
rect 27974 8678 28026 8730
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 2780 8576 2832 8628
rect 4068 8576 4120 8628
rect 5540 8576 5592 8628
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 13176 8576 13228 8628
rect 15936 8619 15988 8628
rect 15936 8585 15945 8619
rect 15945 8585 15979 8619
rect 15979 8585 15988 8619
rect 15936 8576 15988 8585
rect 16580 8576 16632 8628
rect 2320 8508 2372 8560
rect 4620 8508 4672 8560
rect 3148 8483 3200 8492
rect 2780 8372 2832 8424
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 5724 8508 5776 8560
rect 6460 8508 6512 8560
rect 6828 8508 6880 8560
rect 6920 8440 6972 8492
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7196 8483 7248 8492
rect 7012 8440 7064 8449
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 7288 8440 7340 8492
rect 9220 8508 9272 8560
rect 12900 8508 12952 8560
rect 16856 8508 16908 8560
rect 19800 8576 19852 8628
rect 23204 8576 23256 8628
rect 19524 8508 19576 8560
rect 19708 8551 19760 8560
rect 19708 8517 19717 8551
rect 19717 8517 19751 8551
rect 19751 8517 19760 8551
rect 19708 8508 19760 8517
rect 11336 8440 11388 8492
rect 13452 8440 13504 8492
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 4712 8372 4764 8424
rect 2136 8304 2188 8356
rect 4160 8304 4212 8356
rect 5908 8372 5960 8424
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11612 8372 11664 8424
rect 18512 8440 18564 8492
rect 18972 8440 19024 8492
rect 22928 8508 22980 8560
rect 23572 8551 23624 8560
rect 23572 8517 23581 8551
rect 23581 8517 23615 8551
rect 23615 8517 23624 8551
rect 23572 8508 23624 8517
rect 21364 8440 21416 8492
rect 25504 8576 25556 8628
rect 18328 8372 18380 8424
rect 18420 8372 18472 8424
rect 19432 8372 19484 8424
rect 23940 8372 23992 8424
rect 24768 8372 24820 8424
rect 5632 8304 5684 8356
rect 8760 8347 8812 8356
rect 8760 8313 8769 8347
rect 8769 8313 8803 8347
rect 8803 8313 8812 8347
rect 8760 8304 8812 8313
rect 18696 8304 18748 8356
rect 15292 8279 15344 8288
rect 15292 8245 15301 8279
rect 15301 8245 15335 8279
rect 15335 8245 15344 8279
rect 15292 8236 15344 8245
rect 18236 8236 18288 8288
rect 20812 8236 20864 8288
rect 4296 8134 4348 8186
rect 4360 8134 4412 8186
rect 4424 8134 4476 8186
rect 4488 8134 4540 8186
rect 4552 8134 4604 8186
rect 10988 8134 11040 8186
rect 11052 8134 11104 8186
rect 11116 8134 11168 8186
rect 11180 8134 11232 8186
rect 11244 8134 11296 8186
rect 17680 8134 17732 8186
rect 17744 8134 17796 8186
rect 17808 8134 17860 8186
rect 17872 8134 17924 8186
rect 17936 8134 17988 8186
rect 24372 8134 24424 8186
rect 24436 8134 24488 8186
rect 24500 8134 24552 8186
rect 24564 8134 24616 8186
rect 24628 8134 24680 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 5816 8032 5868 8084
rect 7196 8032 7248 8084
rect 7380 8032 7432 8084
rect 8944 8032 8996 8084
rect 10232 8032 10284 8084
rect 13728 8032 13780 8084
rect 14188 8032 14240 8084
rect 18604 8032 18656 8084
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 22008 8032 22060 8084
rect 23020 8075 23072 8084
rect 23020 8041 23029 8075
rect 23029 8041 23063 8075
rect 23063 8041 23072 8075
rect 23020 8032 23072 8041
rect 26148 8075 26200 8084
rect 26148 8041 26157 8075
rect 26157 8041 26191 8075
rect 26191 8041 26200 8075
rect 26148 8032 26200 8041
rect 6736 7896 6788 7948
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 12716 7939 12768 7948
rect 12716 7905 12725 7939
rect 12725 7905 12759 7939
rect 12759 7905 12768 7939
rect 12716 7896 12768 7905
rect 13820 7896 13872 7948
rect 23296 7939 23348 7948
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 24768 7896 24820 7948
rect 2136 7828 2188 7880
rect 4068 7828 4120 7880
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 8760 7828 8812 7880
rect 10324 7828 10376 7880
rect 13912 7828 13964 7880
rect 15016 7828 15068 7880
rect 16948 7871 17000 7880
rect 3332 7803 3384 7812
rect 3332 7769 3341 7803
rect 3341 7769 3375 7803
rect 3375 7769 3384 7803
rect 3332 7760 3384 7769
rect 7564 7760 7616 7812
rect 15200 7760 15252 7812
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 18420 7828 18472 7880
rect 18144 7803 18196 7812
rect 18144 7769 18153 7803
rect 18153 7769 18187 7803
rect 18187 7769 18196 7803
rect 18144 7760 18196 7769
rect 20812 7803 20864 7812
rect 20812 7769 20821 7803
rect 20821 7769 20855 7803
rect 20855 7769 20864 7803
rect 20812 7760 20864 7769
rect 23756 7828 23808 7880
rect 25136 7871 25188 7880
rect 25136 7837 25145 7871
rect 25145 7837 25179 7871
rect 25179 7837 25188 7871
rect 25136 7828 25188 7837
rect 25228 7828 25280 7880
rect 26148 7828 26200 7880
rect 22652 7760 22704 7812
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 14832 7692 14884 7744
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 17960 7692 18012 7744
rect 20168 7735 20220 7744
rect 20168 7701 20177 7735
rect 20177 7701 20211 7735
rect 20211 7701 20220 7735
rect 20168 7692 20220 7701
rect 7642 7590 7694 7642
rect 7706 7590 7758 7642
rect 7770 7590 7822 7642
rect 7834 7590 7886 7642
rect 7898 7590 7950 7642
rect 14334 7590 14386 7642
rect 14398 7590 14450 7642
rect 14462 7590 14514 7642
rect 14526 7590 14578 7642
rect 14590 7590 14642 7642
rect 21026 7590 21078 7642
rect 21090 7590 21142 7642
rect 21154 7590 21206 7642
rect 21218 7590 21270 7642
rect 21282 7590 21334 7642
rect 27718 7590 27770 7642
rect 27782 7590 27834 7642
rect 27846 7590 27898 7642
rect 27910 7590 27962 7642
rect 27974 7590 28026 7642
rect 3332 7488 3384 7540
rect 12900 7488 12952 7540
rect 13360 7488 13412 7540
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 18144 7488 18196 7540
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 22560 7488 22612 7540
rect 12992 7420 13044 7472
rect 14832 7463 14884 7472
rect 14832 7429 14841 7463
rect 14841 7429 14875 7463
rect 14875 7429 14884 7463
rect 14832 7420 14884 7429
rect 18328 7420 18380 7472
rect 2136 7352 2188 7404
rect 3240 7352 3292 7404
rect 5632 7352 5684 7404
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 6276 7352 6328 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 7472 7352 7524 7404
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 12072 7352 12124 7404
rect 13544 7352 13596 7404
rect 15936 7352 15988 7404
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 18604 7395 18656 7404
rect 4160 7284 4212 7336
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 15292 7284 15344 7336
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 18880 7352 18932 7404
rect 19524 7352 19576 7404
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 21364 7352 21416 7404
rect 17960 7327 18012 7336
rect 3516 7216 3568 7268
rect 6920 7216 6972 7268
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 11336 7148 11388 7200
rect 15016 7148 15068 7200
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18972 7284 19024 7336
rect 20720 7284 20772 7336
rect 23940 7488 23992 7540
rect 22836 7420 22888 7472
rect 24400 7327 24452 7336
rect 24400 7293 24409 7327
rect 24409 7293 24443 7327
rect 24443 7293 24452 7327
rect 24400 7284 24452 7293
rect 20904 7148 20956 7200
rect 23480 7148 23532 7200
rect 24400 7148 24452 7200
rect 4296 7046 4348 7098
rect 4360 7046 4412 7098
rect 4424 7046 4476 7098
rect 4488 7046 4540 7098
rect 4552 7046 4604 7098
rect 10988 7046 11040 7098
rect 11052 7046 11104 7098
rect 11116 7046 11168 7098
rect 11180 7046 11232 7098
rect 11244 7046 11296 7098
rect 17680 7046 17732 7098
rect 17744 7046 17796 7098
rect 17808 7046 17860 7098
rect 17872 7046 17924 7098
rect 17936 7046 17988 7098
rect 24372 7046 24424 7098
rect 24436 7046 24488 7098
rect 24500 7046 24552 7098
rect 24564 7046 24616 7098
rect 24628 7046 24680 7098
rect 4160 6987 4212 6996
rect 4160 6953 4169 6987
rect 4169 6953 4203 6987
rect 4203 6953 4212 6987
rect 4160 6944 4212 6953
rect 5356 6944 5408 6996
rect 15200 6944 15252 6996
rect 16488 6944 16540 6996
rect 20168 6944 20220 6996
rect 12532 6876 12584 6928
rect 8208 6851 8260 6860
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 8208 6808 8260 6817
rect 10784 6808 10836 6860
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 5264 6740 5316 6792
rect 7196 6740 7248 6792
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 9128 6740 9180 6792
rect 13452 6783 13504 6792
rect 3976 6715 4028 6724
rect 3976 6681 3985 6715
rect 3985 6681 4019 6715
rect 4019 6681 4028 6715
rect 3976 6672 4028 6681
rect 4068 6604 4120 6656
rect 4988 6672 5040 6724
rect 6552 6672 6604 6724
rect 10600 6672 10652 6724
rect 10968 6672 11020 6724
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 13728 6740 13780 6792
rect 17224 6783 17276 6792
rect 4804 6647 4856 6656
rect 4804 6613 4813 6647
rect 4813 6613 4847 6647
rect 4847 6613 4856 6647
rect 4804 6604 4856 6613
rect 5172 6604 5224 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 11428 6604 11480 6656
rect 11888 6604 11940 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 16120 6672 16172 6724
rect 16488 6604 16540 6656
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 18512 6808 18564 6860
rect 19340 6808 19392 6860
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 22652 6851 22704 6860
rect 22652 6817 22661 6851
rect 22661 6817 22695 6851
rect 22695 6817 22704 6851
rect 22652 6808 22704 6817
rect 18604 6740 18656 6792
rect 19984 6740 20036 6792
rect 22284 6740 22336 6792
rect 23480 6808 23532 6860
rect 20904 6672 20956 6724
rect 21180 6672 21232 6724
rect 17224 6604 17276 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 19340 6604 19392 6656
rect 19708 6604 19760 6656
rect 7642 6502 7694 6554
rect 7706 6502 7758 6554
rect 7770 6502 7822 6554
rect 7834 6502 7886 6554
rect 7898 6502 7950 6554
rect 14334 6502 14386 6554
rect 14398 6502 14450 6554
rect 14462 6502 14514 6554
rect 14526 6502 14578 6554
rect 14590 6502 14642 6554
rect 21026 6502 21078 6554
rect 21090 6502 21142 6554
rect 21154 6502 21206 6554
rect 21218 6502 21270 6554
rect 21282 6502 21334 6554
rect 27718 6502 27770 6554
rect 27782 6502 27834 6554
rect 27846 6502 27898 6554
rect 27910 6502 27962 6554
rect 27974 6502 28026 6554
rect 3976 6400 4028 6452
rect 7472 6400 7524 6452
rect 8116 6400 8168 6452
rect 9220 6400 9272 6452
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2872 6264 2924 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 8300 6332 8352 6384
rect 10508 6332 10560 6384
rect 4068 6264 4120 6273
rect 6920 6264 6972 6316
rect 9956 6264 10008 6316
rect 10968 6264 11020 6316
rect 11704 6400 11756 6452
rect 13912 6400 13964 6452
rect 15936 6443 15988 6452
rect 15936 6409 15945 6443
rect 15945 6409 15979 6443
rect 15979 6409 15988 6443
rect 15936 6400 15988 6409
rect 16488 6400 16540 6452
rect 18972 6400 19024 6452
rect 19524 6400 19576 6452
rect 19984 6400 20036 6452
rect 22836 6443 22888 6452
rect 22836 6409 22845 6443
rect 22845 6409 22879 6443
rect 22879 6409 22888 6443
rect 22836 6400 22888 6409
rect 12624 6332 12676 6384
rect 17224 6332 17276 6384
rect 17592 6332 17644 6384
rect 19340 6375 19392 6384
rect 19340 6341 19349 6375
rect 19349 6341 19383 6375
rect 19383 6341 19392 6375
rect 19340 6332 19392 6341
rect 19616 6332 19668 6384
rect 11612 6264 11664 6316
rect 13452 6264 13504 6316
rect 15568 6307 15620 6316
rect 3516 6196 3568 6248
rect 5540 6196 5592 6248
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 8024 6196 8076 6248
rect 9864 6196 9916 6248
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 15108 6196 15160 6248
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 25228 6332 25280 6384
rect 16856 6239 16908 6248
rect 4160 6060 4212 6112
rect 4896 6060 4948 6112
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 18420 6196 18472 6248
rect 18512 6060 18564 6112
rect 25136 6264 25188 6316
rect 4296 5958 4348 6010
rect 4360 5958 4412 6010
rect 4424 5958 4476 6010
rect 4488 5958 4540 6010
rect 4552 5958 4604 6010
rect 10988 5958 11040 6010
rect 11052 5958 11104 6010
rect 11116 5958 11168 6010
rect 11180 5958 11232 6010
rect 11244 5958 11296 6010
rect 17680 5958 17732 6010
rect 17744 5958 17796 6010
rect 17808 5958 17860 6010
rect 17872 5958 17924 6010
rect 17936 5958 17988 6010
rect 24372 5958 24424 6010
rect 24436 5958 24488 6010
rect 24500 5958 24552 6010
rect 24564 5958 24616 6010
rect 24628 5958 24680 6010
rect 2320 5856 2372 5908
rect 2872 5856 2924 5908
rect 4712 5856 4764 5908
rect 6276 5856 6328 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 14004 5856 14056 5908
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 20904 5856 20956 5908
rect 2780 5788 2832 5840
rect 13452 5788 13504 5840
rect 13728 5831 13780 5840
rect 13728 5797 13737 5831
rect 13737 5797 13771 5831
rect 13771 5797 13780 5831
rect 13728 5788 13780 5797
rect 2136 5652 2188 5704
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 3884 5720 3936 5772
rect 5908 5763 5960 5772
rect 3516 5652 3568 5704
rect 3056 5584 3108 5636
rect 2320 5516 2372 5568
rect 4620 5652 4672 5704
rect 5908 5729 5917 5763
rect 5917 5729 5951 5763
rect 5951 5729 5960 5763
rect 5908 5720 5960 5729
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 11336 5720 11388 5772
rect 5632 5695 5684 5704
rect 4712 5584 4764 5636
rect 4068 5516 4120 5568
rect 4896 5516 4948 5568
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8852 5652 8904 5704
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10784 5652 10836 5704
rect 6000 5584 6052 5636
rect 11796 5584 11848 5636
rect 6828 5516 6880 5568
rect 8208 5516 8260 5568
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 17592 5720 17644 5772
rect 18788 5720 18840 5772
rect 19708 5763 19760 5772
rect 19708 5729 19717 5763
rect 19717 5729 19751 5763
rect 19751 5729 19760 5763
rect 19708 5720 19760 5729
rect 15016 5652 15068 5704
rect 15108 5652 15160 5704
rect 15568 5652 15620 5704
rect 16488 5652 16540 5704
rect 18512 5652 18564 5704
rect 18880 5584 18932 5636
rect 20720 5584 20772 5636
rect 7642 5414 7694 5466
rect 7706 5414 7758 5466
rect 7770 5414 7822 5466
rect 7834 5414 7886 5466
rect 7898 5414 7950 5466
rect 14334 5414 14386 5466
rect 14398 5414 14450 5466
rect 14462 5414 14514 5466
rect 14526 5414 14578 5466
rect 14590 5414 14642 5466
rect 21026 5414 21078 5466
rect 21090 5414 21142 5466
rect 21154 5414 21206 5466
rect 21218 5414 21270 5466
rect 21282 5414 21334 5466
rect 27718 5414 27770 5466
rect 27782 5414 27834 5466
rect 27846 5414 27898 5466
rect 27910 5414 27962 5466
rect 27974 5414 28026 5466
rect 3148 5312 3200 5364
rect 5632 5312 5684 5364
rect 7196 5312 7248 5364
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 11796 5312 11848 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 15108 5312 15160 5364
rect 18880 5312 18932 5364
rect 2320 5244 2372 5296
rect 4160 5244 4212 5296
rect 4896 5244 4948 5296
rect 9128 5287 9180 5296
rect 9128 5253 9137 5287
rect 9137 5253 9171 5287
rect 9171 5253 9180 5287
rect 9128 5244 9180 5253
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 16856 5287 16908 5296
rect 16856 5253 16865 5287
rect 16865 5253 16899 5287
rect 16899 5253 16908 5287
rect 16856 5244 16908 5253
rect 20812 5244 20864 5296
rect 2872 5219 2924 5228
rect 2872 5185 2906 5219
rect 2906 5185 2924 5219
rect 2872 5176 2924 5185
rect 4988 5176 5040 5228
rect 5356 5176 5408 5228
rect 6184 5176 6236 5228
rect 7472 5176 7524 5228
rect 7656 5219 7708 5228
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 8852 5219 8904 5228
rect 8852 5185 8861 5219
rect 8861 5185 8895 5219
rect 8895 5185 8904 5219
rect 8852 5176 8904 5185
rect 9956 5176 10008 5228
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11888 5176 11940 5228
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 2044 5108 2096 5160
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 5540 5108 5592 5160
rect 7104 5108 7156 5160
rect 4620 5040 4672 5092
rect 3976 5015 4028 5024
rect 3976 4981 3985 5015
rect 3985 4981 4019 5015
rect 4019 4981 4028 5015
rect 3976 4972 4028 4981
rect 4160 4972 4212 5024
rect 4296 4870 4348 4922
rect 4360 4870 4412 4922
rect 4424 4870 4476 4922
rect 4488 4870 4540 4922
rect 4552 4870 4604 4922
rect 10988 4870 11040 4922
rect 11052 4870 11104 4922
rect 11116 4870 11168 4922
rect 11180 4870 11232 4922
rect 11244 4870 11296 4922
rect 17680 4870 17732 4922
rect 17744 4870 17796 4922
rect 17808 4870 17860 4922
rect 17872 4870 17924 4922
rect 17936 4870 17988 4922
rect 24372 4870 24424 4922
rect 24436 4870 24488 4922
rect 24500 4870 24552 4922
rect 24564 4870 24616 4922
rect 24628 4870 24680 4922
rect 3516 4768 3568 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 8576 4768 8628 4820
rect 10784 4768 10836 4820
rect 3424 4700 3476 4752
rect 4068 4700 4120 4752
rect 2780 4632 2832 4684
rect 3056 4632 3108 4684
rect 4988 4632 5040 4684
rect 7656 4632 7708 4684
rect 9956 4632 10008 4684
rect 3884 4564 3936 4616
rect 5172 4564 5224 4616
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 2780 4496 2832 4548
rect 3976 4496 4028 4548
rect 9036 4564 9088 4616
rect 2320 4428 2372 4480
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3424 4428 3476 4480
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 9864 4471 9916 4480
rect 9864 4437 9873 4471
rect 9873 4437 9907 4471
rect 9907 4437 9916 4471
rect 9864 4428 9916 4437
rect 7642 4326 7694 4378
rect 7706 4326 7758 4378
rect 7770 4326 7822 4378
rect 7834 4326 7886 4378
rect 7898 4326 7950 4378
rect 14334 4326 14386 4378
rect 14398 4326 14450 4378
rect 14462 4326 14514 4378
rect 14526 4326 14578 4378
rect 14590 4326 14642 4378
rect 21026 4326 21078 4378
rect 21090 4326 21142 4378
rect 21154 4326 21206 4378
rect 21218 4326 21270 4378
rect 21282 4326 21334 4378
rect 27718 4326 27770 4378
rect 27782 4326 27834 4378
rect 27846 4326 27898 4378
rect 27910 4326 27962 4378
rect 27974 4326 28026 4378
rect 3884 4224 3936 4276
rect 4988 4267 5040 4276
rect 4988 4233 4997 4267
rect 4997 4233 5031 4267
rect 5031 4233 5040 4267
rect 4988 4224 5040 4233
rect 2964 4156 3016 4208
rect 4068 4156 4120 4208
rect 5172 4199 5224 4208
rect 5172 4165 5199 4199
rect 5199 4165 5224 4199
rect 5172 4156 5224 4165
rect 1492 4088 1544 4140
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 2780 4088 2832 4140
rect 7380 4088 7432 4140
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19616 4131 19668 4140
rect 19616 4097 19625 4131
rect 19625 4097 19659 4131
rect 19659 4097 19668 4131
rect 19616 4088 19668 4097
rect 2596 4020 2648 4072
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 2780 3952 2832 4004
rect 9864 3952 9916 4004
rect 2136 3884 2188 3936
rect 2872 3884 2924 3936
rect 4344 3884 4396 3936
rect 4712 3884 4764 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 4296 3782 4348 3834
rect 4360 3782 4412 3834
rect 4424 3782 4476 3834
rect 4488 3782 4540 3834
rect 4552 3782 4604 3834
rect 10988 3782 11040 3834
rect 11052 3782 11104 3834
rect 11116 3782 11168 3834
rect 11180 3782 11232 3834
rect 11244 3782 11296 3834
rect 17680 3782 17732 3834
rect 17744 3782 17796 3834
rect 17808 3782 17860 3834
rect 17872 3782 17924 3834
rect 17936 3782 17988 3834
rect 24372 3782 24424 3834
rect 24436 3782 24488 3834
rect 24500 3782 24552 3834
rect 24564 3782 24616 3834
rect 24628 3782 24680 3834
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4620 3680 4672 3732
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 5448 3680 5500 3732
rect 5724 3680 5776 3732
rect 6828 3680 6880 3732
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 2596 3476 2648 3528
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 5172 3476 5224 3528
rect 2320 3451 2372 3460
rect 2320 3417 2354 3451
rect 2354 3417 2372 3451
rect 2320 3408 2372 3417
rect 7642 3238 7694 3290
rect 7706 3238 7758 3290
rect 7770 3238 7822 3290
rect 7834 3238 7886 3290
rect 7898 3238 7950 3290
rect 14334 3238 14386 3290
rect 14398 3238 14450 3290
rect 14462 3238 14514 3290
rect 14526 3238 14578 3290
rect 14590 3238 14642 3290
rect 21026 3238 21078 3290
rect 21090 3238 21142 3290
rect 21154 3238 21206 3290
rect 21218 3238 21270 3290
rect 21282 3238 21334 3290
rect 27718 3238 27770 3290
rect 27782 3238 27834 3290
rect 27846 3238 27898 3290
rect 27910 3238 27962 3290
rect 27974 3238 28026 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 3332 3111 3384 3120
rect 3332 3077 3341 3111
rect 3341 3077 3375 3111
rect 3375 3077 3384 3111
rect 3332 3068 3384 3077
rect 4160 3068 4212 3120
rect 2780 3000 2832 3052
rect 2596 2932 2648 2984
rect 4296 2694 4348 2746
rect 4360 2694 4412 2746
rect 4424 2694 4476 2746
rect 4488 2694 4540 2746
rect 4552 2694 4604 2746
rect 10988 2694 11040 2746
rect 11052 2694 11104 2746
rect 11116 2694 11168 2746
rect 11180 2694 11232 2746
rect 11244 2694 11296 2746
rect 17680 2694 17732 2746
rect 17744 2694 17796 2746
rect 17808 2694 17860 2746
rect 17872 2694 17924 2746
rect 17936 2694 17988 2746
rect 24372 2694 24424 2746
rect 24436 2694 24488 2746
rect 24500 2694 24552 2746
rect 24564 2694 24616 2746
rect 24628 2694 24680 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 3056 2592 3108 2644
rect 3608 2592 3660 2644
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 3792 2524 3844 2576
rect 8116 2524 8168 2576
rect 5724 2456 5776 2508
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 7642 2150 7694 2202
rect 7706 2150 7758 2202
rect 7770 2150 7822 2202
rect 7834 2150 7886 2202
rect 7898 2150 7950 2202
rect 14334 2150 14386 2202
rect 14398 2150 14450 2202
rect 14462 2150 14514 2202
rect 14526 2150 14578 2202
rect 14590 2150 14642 2202
rect 21026 2150 21078 2202
rect 21090 2150 21142 2202
rect 21154 2150 21206 2202
rect 21218 2150 21270 2202
rect 21282 2150 21334 2202
rect 27718 2150 27770 2202
rect 27782 2150 27834 2202
rect 27846 2150 27898 2202
rect 27910 2150 27962 2202
rect 27974 2150 28026 2202
<< metal2 >>
rect 1858 28200 1914 29000
rect 5446 28200 5502 29000
rect 9034 28200 9090 29000
rect 12622 28200 12678 29000
rect 16210 28200 16266 29000
rect 19798 28200 19854 29000
rect 23386 28200 23442 29000
rect 26974 28200 27030 29000
rect 1674 26888 1730 26897
rect 1674 26823 1730 26832
rect 1688 26382 1716 26823
rect 1872 26586 1900 28200
rect 4296 26684 4604 26693
rect 4296 26682 4302 26684
rect 4358 26682 4382 26684
rect 4438 26682 4462 26684
rect 4518 26682 4542 26684
rect 4598 26682 4604 26684
rect 4358 26630 4360 26682
rect 4540 26630 4542 26682
rect 4296 26628 4302 26630
rect 4358 26628 4382 26630
rect 4438 26628 4462 26630
rect 4518 26628 4542 26630
rect 4598 26628 4604 26630
rect 4296 26619 4604 26628
rect 5460 26586 5488 28200
rect 9048 26586 9076 28200
rect 10988 26684 11296 26693
rect 10988 26682 10994 26684
rect 11050 26682 11074 26684
rect 11130 26682 11154 26684
rect 11210 26682 11234 26684
rect 11290 26682 11296 26684
rect 11050 26630 11052 26682
rect 11232 26630 11234 26682
rect 10988 26628 10994 26630
rect 11050 26628 11074 26630
rect 11130 26628 11154 26630
rect 11210 26628 11234 26630
rect 11290 26628 11296 26630
rect 10988 26619 11296 26628
rect 1860 26580 1912 26586
rect 1860 26522 1912 26528
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 9036 26580 9088 26586
rect 9036 26522 9088 26528
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 4528 26376 4580 26382
rect 4528 26318 4580 26324
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 1688 26042 1716 26318
rect 4540 26042 4568 26318
rect 5000 26042 5028 26318
rect 5080 26308 5132 26314
rect 5080 26250 5132 26256
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 4528 26036 4580 26042
rect 4528 25978 4580 25984
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2228 25696 2280 25702
rect 2228 25638 2280 25644
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 1676 25220 1728 25226
rect 1676 25162 1728 25168
rect 1688 23866 1716 25162
rect 2056 24138 2084 25230
rect 2240 24206 2268 25638
rect 2516 24954 2544 25774
rect 2504 24948 2556 24954
rect 2504 24890 2556 24896
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2044 24132 2096 24138
rect 2044 24074 2096 24080
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 2976 23730 3004 25842
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4296 25596 4604 25605
rect 4296 25594 4302 25596
rect 4358 25594 4382 25596
rect 4438 25594 4462 25596
rect 4518 25594 4542 25596
rect 4598 25594 4604 25596
rect 4358 25542 4360 25594
rect 4540 25542 4542 25594
rect 4296 25540 4302 25542
rect 4358 25540 4382 25542
rect 4438 25540 4462 25542
rect 4518 25540 4542 25542
rect 4598 25540 4604 25542
rect 4296 25531 4604 25540
rect 4816 25498 4844 25774
rect 4804 25492 4856 25498
rect 4804 25434 4856 25440
rect 4160 25424 4212 25430
rect 4160 25366 4212 25372
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3620 24138 3648 24686
rect 3988 24410 4016 24754
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 4172 24274 4200 25366
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4356 24954 4384 25230
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4724 24886 4752 25230
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4816 24682 4844 25162
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4296 24508 4604 24517
rect 4296 24506 4302 24508
rect 4358 24506 4382 24508
rect 4438 24506 4462 24508
rect 4518 24506 4542 24508
rect 4598 24506 4604 24508
rect 4358 24454 4360 24506
rect 4540 24454 4542 24506
rect 4296 24452 4302 24454
rect 4358 24452 4382 24454
rect 4438 24452 4462 24454
rect 4518 24452 4542 24454
rect 4598 24452 4604 24454
rect 4296 24443 4604 24452
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 3056 24132 3108 24138
rect 3056 24074 3108 24080
rect 3608 24132 3660 24138
rect 3608 24074 3660 24080
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2044 22976 2096 22982
rect 2044 22918 2096 22924
rect 2056 22574 2084 22918
rect 2976 22642 3004 23666
rect 3068 23662 3096 24074
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 3252 23118 3280 24006
rect 4724 23730 4752 24142
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3344 23118 3372 23598
rect 3528 23361 3556 23666
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 3514 23352 3570 23361
rect 3514 23287 3570 23296
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3528 22778 3556 23287
rect 4172 23186 4200 23598
rect 4296 23420 4604 23429
rect 4296 23418 4302 23420
rect 4358 23418 4382 23420
rect 4438 23418 4462 23420
rect 4518 23418 4542 23420
rect 4598 23418 4604 23420
rect 4358 23366 4360 23418
rect 4540 23366 4542 23418
rect 4296 23364 4302 23366
rect 4358 23364 4382 23366
rect 4438 23364 4462 23366
rect 4518 23364 4542 23366
rect 4598 23364 4604 23366
rect 4296 23355 4604 23364
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 1860 22432 1912 22438
rect 1860 22374 1912 22380
rect 3516 22432 3568 22438
rect 3516 22374 3568 22380
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 1504 21010 1532 21422
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 1504 19922 1532 20946
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1596 17202 1624 21286
rect 1688 20466 1716 21830
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1688 19825 1716 20402
rect 1872 19854 1900 22374
rect 3528 21894 3556 22374
rect 3896 22030 3924 23054
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4296 22332 4604 22341
rect 4296 22330 4302 22332
rect 4358 22330 4382 22332
rect 4438 22330 4462 22332
rect 4518 22330 4542 22332
rect 4598 22330 4604 22332
rect 4358 22278 4360 22330
rect 4540 22278 4542 22330
rect 4296 22276 4302 22278
rect 4358 22276 4382 22278
rect 4438 22276 4462 22278
rect 4518 22276 4542 22278
rect 4598 22276 4604 22278
rect 4296 22267 4604 22276
rect 4632 22098 4660 22986
rect 4724 22642 4752 23666
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4724 22234 4752 22578
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3528 21690 3556 21830
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2700 21146 2728 21422
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2792 20602 2820 20742
rect 3436 20602 3464 21558
rect 3528 20874 3556 21626
rect 3896 21486 3924 21966
rect 4632 21690 4660 22034
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3896 21010 3924 21422
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3240 20528 3292 20534
rect 3528 20482 3556 20810
rect 3292 20476 3556 20482
rect 3240 20470 3556 20476
rect 3252 20466 3556 20470
rect 3896 20466 3924 20946
rect 3252 20460 3568 20466
rect 3252 20454 3516 20460
rect 3516 20402 3568 20408
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 1860 19848 1912 19854
rect 1674 19816 1730 19825
rect 1860 19790 1912 19796
rect 1674 19751 1730 19760
rect 3528 19718 3556 20402
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 2976 19446 3004 19654
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17746 1992 18022
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 2240 17338 2268 18566
rect 2608 18358 2636 18566
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2976 17882 3004 19246
rect 3344 18290 3372 19450
rect 3528 18630 3556 19654
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3068 17338 3096 17614
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2240 17218 2268 17274
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 2148 17190 2268 17218
rect 3528 17202 3556 18566
rect 3988 18222 4016 21490
rect 4296 21244 4604 21253
rect 4296 21242 4302 21244
rect 4358 21242 4382 21244
rect 4438 21242 4462 21244
rect 4518 21242 4542 21244
rect 4598 21242 4604 21244
rect 4358 21190 4360 21242
rect 4540 21190 4542 21242
rect 4296 21188 4302 21190
rect 4358 21188 4382 21190
rect 4438 21188 4462 21190
rect 4518 21188 4542 21190
rect 4598 21188 4604 21190
rect 4296 21179 4604 21188
rect 5000 20942 5028 21490
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 4816 20806 4844 20878
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4724 20534 4752 20742
rect 4816 20584 4844 20742
rect 4896 20596 4948 20602
rect 4816 20556 4896 20584
rect 4712 20528 4764 20534
rect 4712 20470 4764 20476
rect 4296 20156 4604 20165
rect 4296 20154 4302 20156
rect 4358 20154 4382 20156
rect 4438 20154 4462 20156
rect 4518 20154 4542 20156
rect 4598 20154 4604 20156
rect 4358 20102 4360 20154
rect 4540 20102 4542 20154
rect 4296 20100 4302 20102
rect 4358 20100 4382 20102
rect 4438 20100 4462 20102
rect 4518 20100 4542 20102
rect 4598 20100 4604 20102
rect 4296 20091 4604 20100
rect 4816 19514 4844 20556
rect 4896 20538 4948 20544
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4816 19258 4844 19450
rect 4724 19230 4844 19258
rect 4296 19068 4604 19077
rect 4296 19066 4302 19068
rect 4358 19066 4382 19068
rect 4438 19066 4462 19068
rect 4518 19066 4542 19068
rect 4598 19066 4604 19068
rect 4358 19014 4360 19066
rect 4540 19014 4542 19066
rect 4296 19012 4302 19014
rect 4358 19012 4382 19014
rect 4438 19012 4462 19014
rect 4518 19012 4542 19014
rect 4598 19012 4604 19014
rect 4296 19003 4604 19012
rect 4724 18766 4752 19230
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3988 17882 4016 18158
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3988 17678 4016 17818
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3516 17196 3568 17202
rect 1596 16289 1624 17138
rect 1768 17060 1820 17066
rect 1768 17002 1820 17008
rect 1582 16280 1638 16289
rect 1582 16215 1638 16224
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15094 1716 15438
rect 1676 15088 1728 15094
rect 1676 15030 1728 15036
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14482 1716 14758
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1582 12744 1638 12753
rect 1582 12679 1638 12688
rect 1596 12170 1624 12679
rect 1584 12164 1636 12170
rect 1584 12106 1636 12112
rect 1490 5672 1546 5681
rect 1490 5607 1546 5616
rect 1504 4146 1532 5607
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1596 2650 1624 12106
rect 1688 10266 1716 14418
rect 1780 14074 1808 17002
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2056 16182 2084 16390
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 2148 14362 2176 17190
rect 3516 17138 3568 17144
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2240 16250 2268 16526
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2240 15026 2268 16186
rect 2792 16046 2820 16390
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 15094 2912 15302
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 1860 14340 1912 14346
rect 2148 14334 2360 14362
rect 1860 14282 1912 14288
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1768 13796 1820 13802
rect 1768 13738 1820 13744
rect 1780 12850 1808 13738
rect 1872 12986 1900 14282
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2148 14006 2176 14214
rect 2240 14074 2268 14214
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1964 12986 1992 13262
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2240 12850 2268 13126
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 2056 9586 2084 12106
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2148 10810 2176 11018
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2056 9178 2084 9522
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 8090 2084 9114
rect 2148 8362 2176 9998
rect 2332 8566 2360 14334
rect 2504 14000 2556 14006
rect 2504 13942 2556 13948
rect 2516 13326 2544 13942
rect 2792 13938 2820 14962
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3068 14074 3096 14282
rect 3344 14074 3372 15370
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3436 15026 3464 15302
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12918 2820 13194
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2792 12238 2820 12854
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 11150 2912 11494
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2884 10470 2912 11086
rect 2872 10464 2924 10470
rect 2924 10412 3004 10418
rect 2872 10406 3004 10412
rect 2884 10390 3004 10406
rect 2976 10062 3004 10390
rect 2964 10056 3016 10062
rect 2792 10004 2964 10010
rect 2792 9998 3016 10004
rect 2792 9982 3004 9998
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2516 9654 2544 9862
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 8634 2728 8842
rect 2792 8634 2820 9982
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9217 3004 9862
rect 2962 9208 3018 9217
rect 2962 9143 3018 9152
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7410 2176 7822
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2056 6322 2084 6734
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5166 2084 6258
rect 2148 5710 2176 7346
rect 2332 5914 2360 8502
rect 2792 8430 2820 8570
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2884 5914 2912 6258
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2148 3942 2176 5646
rect 2332 5574 2360 5850
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5302 2360 5510
rect 2320 5296 2372 5302
rect 2240 5244 2320 5250
rect 2240 5238 2372 5244
rect 2240 5222 2360 5238
rect 2240 4146 2268 5222
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 3194 2084 3470
rect 2332 3466 2360 4422
rect 2608 4078 2636 5102
rect 2792 4690 2820 5782
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2792 4146 2820 4490
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2608 3534 2636 4014
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2608 2990 2636 3470
rect 2792 3058 2820 3946
rect 2884 3942 2912 5170
rect 2976 4570 3004 9143
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3160 8498 3188 8978
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3344 7546 3372 7754
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3068 4690 3096 5578
rect 3160 5370 3188 5646
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2976 4542 3096 4570
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2976 4214 3004 4422
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 3068 2650 3096 4542
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3252 2310 3280 7346
rect 3344 3126 3372 7482
rect 3528 7274 3556 17138
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3804 16250 3832 16526
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 3712 15162 3740 16118
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3896 9654 3924 16526
rect 3988 14414 4016 17614
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17338 4108 17478
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4172 17202 4200 18702
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4296 17980 4604 17989
rect 4296 17978 4302 17980
rect 4358 17978 4382 17980
rect 4438 17978 4462 17980
rect 4518 17978 4542 17980
rect 4598 17978 4604 17980
rect 4358 17926 4360 17978
rect 4540 17926 4542 17978
rect 4296 17924 4302 17926
rect 4358 17924 4382 17926
rect 4438 17924 4462 17926
rect 4518 17924 4542 17926
rect 4598 17924 4604 17926
rect 4296 17915 4604 17924
rect 4632 17338 4660 18226
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4724 17202 4752 18702
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4080 15434 4108 16730
rect 4172 15706 4200 17002
rect 4296 16892 4604 16901
rect 4296 16890 4302 16892
rect 4358 16890 4382 16892
rect 4438 16890 4462 16892
rect 4518 16890 4542 16892
rect 4598 16890 4604 16892
rect 4358 16838 4360 16890
rect 4540 16838 4542 16890
rect 4296 16836 4302 16838
rect 4358 16836 4382 16838
rect 4438 16836 4462 16838
rect 4518 16836 4542 16838
rect 4598 16836 4604 16838
rect 4296 16827 4604 16836
rect 4816 16590 4844 19110
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4908 16402 4936 20198
rect 5092 19718 5120 26250
rect 5368 24274 5396 26250
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5460 25362 5488 25842
rect 5540 25424 5592 25430
rect 5540 25366 5592 25372
rect 5448 25356 5500 25362
rect 5448 25298 5500 25304
rect 5460 24954 5488 25298
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5552 24070 5580 25366
rect 5736 25294 5764 26386
rect 6552 26376 6604 26382
rect 6552 26318 6604 26324
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 5908 26240 5960 26246
rect 5908 26182 5960 26188
rect 5920 25838 5948 26182
rect 5908 25832 5960 25838
rect 5908 25774 5960 25780
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5644 24818 5672 25094
rect 5736 24954 5764 25230
rect 5816 25220 5868 25226
rect 5816 25162 5868 25168
rect 5724 24948 5776 24954
rect 5724 24890 5776 24896
rect 5828 24818 5856 25162
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5644 23866 5672 24754
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 5736 24138 5764 24686
rect 5920 24614 5948 25230
rect 6380 25158 6408 26250
rect 6564 25294 6592 26318
rect 7642 26140 7950 26149
rect 7642 26138 7648 26140
rect 7704 26138 7728 26140
rect 7784 26138 7808 26140
rect 7864 26138 7888 26140
rect 7944 26138 7950 26140
rect 7704 26086 7706 26138
rect 7886 26086 7888 26138
rect 7642 26084 7648 26086
rect 7704 26084 7728 26086
rect 7784 26084 7808 26086
rect 7864 26084 7888 26086
rect 7944 26084 7950 26086
rect 7642 26075 7950 26084
rect 9140 26042 9168 26318
rect 9128 26036 9180 26042
rect 9128 25978 9180 25984
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 6276 24676 6328 24682
rect 6276 24618 6328 24624
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 6288 24154 6316 24618
rect 6380 24410 6408 25094
rect 6748 24886 6776 25842
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 6828 24948 6880 24954
rect 6828 24890 6880 24896
rect 6736 24880 6788 24886
rect 6736 24822 6788 24828
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 6748 24342 6776 24822
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6368 24200 6420 24206
rect 6288 24148 6368 24154
rect 6288 24142 6420 24148
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 6288 24126 6408 24142
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 5736 23322 5764 24074
rect 6288 23594 6316 24126
rect 6748 24070 6776 24278
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6276 23588 6328 23594
rect 6276 23530 6328 23536
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 5736 22094 5764 22986
rect 5644 22066 5764 22094
rect 6288 22094 6316 23530
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6380 22642 6408 23054
rect 6840 23050 6868 24890
rect 7024 24818 7052 25638
rect 7116 25362 7144 25638
rect 7392 25430 7420 25774
rect 9416 25430 9444 26318
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 7380 25424 7432 25430
rect 7380 25366 7432 25372
rect 9404 25424 9456 25430
rect 9404 25366 9456 25372
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 9508 25294 9536 26250
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 8116 25220 8168 25226
rect 8116 25162 8168 25168
rect 8300 25220 8352 25226
rect 8352 25180 8432 25208
rect 8300 25162 8352 25168
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7116 23866 7144 24754
rect 7392 24206 7420 25162
rect 7642 25052 7950 25061
rect 7642 25050 7648 25052
rect 7704 25050 7728 25052
rect 7784 25050 7808 25052
rect 7864 25050 7888 25052
rect 7944 25050 7950 25052
rect 7704 24998 7706 25050
rect 7886 24998 7888 25050
rect 7642 24996 7648 24998
rect 7704 24996 7728 24998
rect 7784 24996 7808 24998
rect 7864 24996 7888 24998
rect 7944 24996 7950 24998
rect 7642 24987 7950 24996
rect 8128 24818 8156 25162
rect 8404 24886 8432 25180
rect 8496 24954 8524 25230
rect 8852 25220 8904 25226
rect 8852 25162 8904 25168
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8392 24880 8444 24886
rect 8392 24822 8444 24828
rect 8116 24812 8168 24818
rect 8116 24754 8168 24760
rect 8300 24608 8352 24614
rect 8300 24550 8352 24556
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 7380 24200 7432 24206
rect 7432 24148 7512 24154
rect 7380 24142 7512 24148
rect 7392 24126 7512 24142
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 6828 23044 6880 23050
rect 6828 22986 6880 22992
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6288 22066 6408 22094
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 5368 21690 5396 21966
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5368 20806 5396 21490
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5368 20330 5396 20742
rect 5552 20602 5580 20878
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5644 20482 5672 22066
rect 5552 20454 5672 20482
rect 5552 20398 5580 20454
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 17270 5120 19654
rect 5276 19378 5304 19926
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5552 17882 5580 20334
rect 6380 19786 6408 22066
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21622 6592 21830
rect 6552 21616 6604 21622
rect 6552 21558 6604 21564
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 20602 6500 20810
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 5920 19514 5948 19722
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5736 18358 5764 19110
rect 6380 18426 6408 19722
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6564 18426 6592 18634
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 5724 18352 5776 18358
rect 5724 18294 5776 18300
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5092 16658 5120 17206
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 4816 16374 4936 16402
rect 4296 15804 4604 15813
rect 4296 15802 4302 15804
rect 4358 15802 4382 15804
rect 4438 15802 4462 15804
rect 4518 15802 4542 15804
rect 4598 15802 4604 15804
rect 4358 15750 4360 15802
rect 4540 15750 4542 15802
rect 4296 15748 4302 15750
rect 4358 15748 4382 15750
rect 4438 15748 4462 15750
rect 4518 15748 4542 15750
rect 4598 15748 4604 15750
rect 4296 15739 4604 15748
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4172 15502 4200 15642
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4172 15094 4200 15438
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 14618 4200 14894
rect 4296 14716 4604 14725
rect 4296 14714 4302 14716
rect 4358 14714 4382 14716
rect 4438 14714 4462 14716
rect 4518 14714 4542 14716
rect 4598 14714 4604 14716
rect 4358 14662 4360 14714
rect 4540 14662 4542 14714
rect 4296 14660 4302 14662
rect 4358 14660 4382 14662
rect 4438 14660 4462 14662
rect 4518 14660 4542 14662
rect 4598 14660 4604 14662
rect 4296 14651 4604 14660
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13512 4200 13806
rect 4296 13628 4604 13637
rect 4296 13626 4302 13628
rect 4358 13626 4382 13628
rect 4438 13626 4462 13628
rect 4518 13626 4542 13628
rect 4598 13626 4604 13628
rect 4358 13574 4360 13626
rect 4540 13574 4542 13626
rect 4296 13572 4302 13574
rect 4358 13572 4382 13574
rect 4438 13572 4462 13574
rect 4518 13572 4542 13574
rect 4598 13572 4604 13574
rect 4296 13563 4604 13572
rect 4172 13484 4292 13512
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12918 4200 13126
rect 4264 12986 4292 13484
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 12986 4752 13262
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4296 12540 4604 12549
rect 4296 12538 4302 12540
rect 4358 12538 4382 12540
rect 4438 12538 4462 12540
rect 4518 12538 4542 12540
rect 4598 12538 4604 12540
rect 4358 12486 4360 12538
rect 4540 12486 4542 12538
rect 4296 12484 4302 12486
rect 4358 12484 4382 12486
rect 4438 12484 4462 12486
rect 4518 12484 4542 12486
rect 4598 12484 4604 12486
rect 4296 12475 4604 12484
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 3988 11762 4016 12038
rect 4448 11898 4476 12038
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4632 11830 4660 12242
rect 4724 12238 4752 12786
rect 4816 12434 4844 16374
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4908 14414 4936 15438
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 5000 14618 5028 15030
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 13938 4936 14350
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4816 12406 4936 12434
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 10674 4200 11494
rect 4296 11452 4604 11461
rect 4296 11450 4302 11452
rect 4358 11450 4382 11452
rect 4438 11450 4462 11452
rect 4518 11450 4542 11452
rect 4598 11450 4604 11452
rect 4358 11398 4360 11450
rect 4540 11398 4542 11450
rect 4296 11396 4302 11398
rect 4358 11396 4382 11398
rect 4438 11396 4462 11398
rect 4518 11396 4542 11398
rect 4598 11396 4604 11398
rect 4296 11387 4604 11396
rect 4632 11218 4660 11766
rect 4724 11626 4752 12174
rect 4908 12102 4936 12406
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11762 4936 12038
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4264 10470 4292 11018
rect 4816 10742 4844 11222
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4908 10554 4936 11698
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5000 11354 5028 11630
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5000 10606 5028 11290
rect 5092 11150 5120 16594
rect 5736 16182 5764 16934
rect 6012 16794 6040 18158
rect 6656 17338 6684 22578
rect 6840 22234 6868 22986
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 7392 22094 7420 24126
rect 7484 24070 7512 24126
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 8024 24064 8076 24070
rect 8024 24006 8076 24012
rect 7642 23964 7950 23973
rect 7642 23962 7648 23964
rect 7704 23962 7728 23964
rect 7784 23962 7808 23964
rect 7864 23962 7888 23964
rect 7944 23962 7950 23964
rect 7704 23910 7706 23962
rect 7886 23910 7888 23962
rect 7642 23908 7648 23910
rect 7704 23908 7728 23910
rect 7784 23908 7808 23910
rect 7864 23908 7888 23910
rect 7944 23908 7950 23910
rect 7642 23899 7950 23908
rect 8036 23798 8064 24006
rect 8128 23866 8156 24210
rect 8208 24132 8260 24138
rect 8208 24074 8260 24080
rect 8220 23866 8248 24074
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8024 23792 8076 23798
rect 8024 23734 8076 23740
rect 8220 23322 8248 23802
rect 8312 23730 8340 24550
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 7642 22876 7950 22885
rect 7642 22874 7648 22876
rect 7704 22874 7728 22876
rect 7784 22874 7808 22876
rect 7864 22874 7888 22876
rect 7944 22874 7950 22876
rect 7704 22822 7706 22874
rect 7886 22822 7888 22874
rect 7642 22820 7648 22822
rect 7704 22820 7728 22822
rect 7784 22820 7808 22822
rect 7864 22820 7888 22822
rect 7944 22820 7950 22822
rect 7642 22811 7950 22820
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 7116 22066 7420 22094
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6840 21146 6868 21422
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6932 20466 6960 20878
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6932 19854 6960 20402
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6748 18290 6776 19110
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6932 17678 6960 19790
rect 7024 19378 7052 20742
rect 7116 19514 7144 22066
rect 7642 21788 7950 21797
rect 7642 21786 7648 21788
rect 7704 21786 7728 21788
rect 7784 21786 7808 21788
rect 7864 21786 7888 21788
rect 7944 21786 7950 21788
rect 7704 21734 7706 21786
rect 7886 21734 7888 21786
rect 7642 21732 7648 21734
rect 7704 21732 7728 21734
rect 7784 21732 7808 21734
rect 7864 21732 7888 21734
rect 7944 21732 7950 21734
rect 7642 21723 7950 21732
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6920 17536 6972 17542
rect 7024 17490 7052 19314
rect 7116 18970 7144 19450
rect 7300 19310 7328 19858
rect 7392 19310 7420 21422
rect 7484 21146 7512 21558
rect 8220 21350 8248 22578
rect 8312 22030 8340 22918
rect 8404 22778 8432 24822
rect 8496 24614 8524 24890
rect 8864 24682 8892 25162
rect 8852 24676 8904 24682
rect 8852 24618 8904 24624
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8864 24342 8892 24618
rect 9140 24410 9168 25230
rect 9220 25152 9272 25158
rect 9220 25094 9272 25100
rect 9232 24614 9260 25094
rect 9508 24886 9536 25230
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 9600 24818 9628 25298
rect 9784 24954 9812 25842
rect 9876 25838 9904 26182
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10704 25294 10732 25774
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10692 25152 10744 25158
rect 10796 25106 10824 25842
rect 11336 25696 11388 25702
rect 11336 25638 11388 25644
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 10988 25596 11296 25605
rect 10988 25594 10994 25596
rect 11050 25594 11074 25596
rect 11130 25594 11154 25596
rect 11210 25594 11234 25596
rect 11290 25594 11296 25596
rect 11050 25542 11052 25594
rect 11232 25542 11234 25594
rect 10988 25540 10994 25542
rect 11050 25540 11074 25542
rect 11130 25540 11154 25542
rect 11210 25540 11234 25542
rect 11290 25540 11296 25542
rect 10988 25531 11296 25540
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10744 25100 10824 25106
rect 10692 25094 10824 25100
rect 10704 25078 10824 25094
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 8852 24336 8904 24342
rect 8852 24278 8904 24284
rect 9232 23866 9260 24550
rect 9508 24410 9536 24618
rect 10704 24410 10732 25078
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10888 24206 10916 25230
rect 11348 24954 11376 25638
rect 11900 25362 11928 25638
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 12084 24818 12112 25842
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 11888 24608 11940 24614
rect 11888 24550 11940 24556
rect 10988 24508 11296 24517
rect 10988 24506 10994 24508
rect 11050 24506 11074 24508
rect 11130 24506 11154 24508
rect 11210 24506 11234 24508
rect 11290 24506 11296 24508
rect 11050 24454 11052 24506
rect 11232 24454 11234 24506
rect 10988 24452 10994 24454
rect 11050 24452 11074 24454
rect 11130 24452 11154 24454
rect 11210 24452 11234 24454
rect 11290 24452 11296 24454
rect 10988 24443 11296 24452
rect 11900 24274 11928 24550
rect 12084 24410 12112 24754
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 11888 24268 11940 24274
rect 11888 24210 11940 24216
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 9404 24132 9456 24138
rect 9404 24074 9456 24080
rect 9416 23866 9444 24074
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9600 23730 9628 24006
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 8220 21010 8248 21286
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7484 20534 7512 20878
rect 7642 20700 7950 20709
rect 7642 20698 7648 20700
rect 7704 20698 7728 20700
rect 7784 20698 7808 20700
rect 7864 20698 7888 20700
rect 7944 20698 7950 20700
rect 7704 20646 7706 20698
rect 7886 20646 7888 20698
rect 7642 20644 7648 20646
rect 7704 20644 7728 20646
rect 7784 20644 7808 20646
rect 7864 20644 7888 20646
rect 7944 20644 7950 20646
rect 7642 20635 7950 20644
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7484 19854 7512 20470
rect 8496 20330 8524 23462
rect 9508 23322 9536 23462
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 9508 23050 9536 23258
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 9232 21962 9260 22510
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 21350 9260 21898
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9232 20874 9260 21286
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7300 18834 7328 19246
rect 7392 18902 7420 19246
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18358 7420 18566
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7484 17678 7512 19790
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 19446 7604 19654
rect 7642 19612 7950 19621
rect 7642 19610 7648 19612
rect 7704 19610 7728 19612
rect 7784 19610 7808 19612
rect 7864 19610 7888 19612
rect 7944 19610 7950 19612
rect 7704 19558 7706 19610
rect 7886 19558 7888 19610
rect 7642 19556 7648 19558
rect 7704 19556 7728 19558
rect 7784 19556 7808 19558
rect 7864 19556 7888 19558
rect 7944 19556 7950 19558
rect 7642 19547 7950 19556
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7840 19304 7892 19310
rect 7892 19264 8064 19292
rect 7840 19246 7892 19252
rect 7642 18524 7950 18533
rect 7642 18522 7648 18524
rect 7704 18522 7728 18524
rect 7784 18522 7808 18524
rect 7864 18522 7888 18524
rect 7944 18522 7950 18524
rect 7704 18470 7706 18522
rect 7886 18470 7888 18522
rect 7642 18468 7648 18470
rect 7704 18468 7728 18470
rect 7784 18468 7808 18470
rect 7864 18468 7888 18470
rect 7944 18468 7950 18470
rect 7642 18459 7950 18468
rect 8036 18222 8064 19264
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 6972 17484 7052 17490
rect 6920 17478 7052 17484
rect 6932 17462 7052 17478
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 6656 16590 6684 17274
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6748 16794 6776 17138
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6932 16658 6960 17462
rect 7642 17436 7950 17445
rect 7642 17434 7648 17436
rect 7704 17434 7728 17436
rect 7784 17434 7808 17436
rect 7864 17434 7888 17436
rect 7944 17434 7950 17436
rect 7704 17382 7706 17434
rect 7886 17382 7888 17434
rect 7642 17380 7648 17382
rect 7704 17380 7728 17382
rect 7784 17380 7808 17382
rect 7864 17380 7888 17382
rect 7944 17380 7950 17382
rect 7642 17371 7950 17380
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7208 16794 7236 16934
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 6012 16114 6040 16390
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 14618 5580 15438
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5828 15162 5856 15370
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 6840 14958 6868 15574
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7116 14890 7144 15438
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5828 14414 5856 14826
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13938 6408 14214
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5368 13326 5396 13738
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5552 13326 5580 13466
rect 6288 13394 6316 13670
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5276 12918 5304 13262
rect 6748 13258 6776 13806
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5368 12434 5396 13126
rect 6564 12968 6592 13194
rect 6644 12980 6696 12986
rect 6564 12940 6644 12968
rect 6644 12922 6696 12928
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5368 12406 5488 12434
rect 5172 12368 5224 12374
rect 5224 12316 5304 12322
rect 5172 12310 5304 12316
rect 5184 12294 5304 12310
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 11354 5212 12174
rect 5276 11812 5304 12294
rect 5460 12170 5488 12406
rect 6012 12170 6040 12582
rect 6932 12442 6960 12650
rect 7116 12442 7144 12922
rect 7208 12832 7236 16730
rect 7944 16726 7972 17070
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8128 16522 8156 20198
rect 8312 18850 8340 20198
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19530 8616 19654
rect 8496 19514 8616 19530
rect 8484 19508 8616 19514
rect 8536 19502 8616 19508
rect 8484 19450 8536 19456
rect 8220 18822 8340 18850
rect 8220 18766 8248 18822
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7642 16348 7950 16357
rect 7642 16346 7648 16348
rect 7704 16346 7728 16348
rect 7784 16346 7808 16348
rect 7864 16346 7888 16348
rect 7944 16346 7950 16348
rect 7704 16294 7706 16346
rect 7886 16294 7888 16346
rect 7642 16292 7648 16294
rect 7704 16292 7728 16294
rect 7784 16292 7808 16294
rect 7864 16292 7888 16294
rect 7944 16292 7950 16294
rect 7642 16283 7950 16292
rect 8036 16114 8064 16390
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15026 7328 15302
rect 7642 15260 7950 15269
rect 7642 15258 7648 15260
rect 7704 15258 7728 15260
rect 7784 15258 7808 15260
rect 7864 15258 7888 15260
rect 7944 15258 7950 15260
rect 7704 15206 7706 15258
rect 7886 15206 7888 15258
rect 7642 15204 7648 15206
rect 7704 15204 7728 15206
rect 7784 15204 7808 15206
rect 7864 15204 7888 15206
rect 7944 15204 7950 15206
rect 7642 15195 7950 15204
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7300 13394 7328 14010
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7288 12844 7340 12850
rect 7208 12804 7288 12832
rect 7288 12786 7340 12792
rect 6920 12436 6972 12442
rect 7104 12436 7156 12442
rect 6972 12396 7052 12424
rect 6920 12378 6972 12384
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6932 12170 6960 12242
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 5448 11824 5500 11830
rect 5276 11784 5448 11812
rect 5448 11766 5500 11772
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4816 10526 4936 10554
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4296 10364 4604 10373
rect 4296 10362 4302 10364
rect 4358 10362 4382 10364
rect 4438 10362 4462 10364
rect 4518 10362 4542 10364
rect 4598 10362 4604 10364
rect 4358 10310 4360 10362
rect 4540 10310 4542 10362
rect 4296 10308 4302 10310
rect 4358 10308 4382 10310
rect 4438 10308 4462 10310
rect 4518 10308 4542 10310
rect 4598 10308 4604 10310
rect 4296 10299 4604 10308
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9654 4200 9862
rect 4540 9722 4568 9998
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3528 5710 3556 6190
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 4826 3556 5646
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3436 4486 3464 4694
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 3738 3464 4422
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3620 2650 3648 9318
rect 3896 8498 3924 9590
rect 4540 9450 4568 9658
rect 4632 9518 4660 10406
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4724 9330 4752 10066
rect 4632 9302 4752 9330
rect 4296 9276 4604 9285
rect 4296 9274 4302 9276
rect 4358 9274 4382 9276
rect 4438 9274 4462 9276
rect 4518 9274 4542 9276
rect 4598 9274 4604 9276
rect 4358 9222 4360 9274
rect 4540 9222 4542 9274
rect 4296 9220 4302 9222
rect 4358 9220 4382 9222
rect 4438 9220 4462 9222
rect 4518 9220 4542 9222
rect 4598 9220 4604 9222
rect 4296 9211 4604 9220
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3884 8492 3936 8498
rect 3804 8452 3884 8480
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3804 2582 3832 8452
rect 3884 8434 3936 8440
rect 4080 7886 4108 8570
rect 4172 8362 4200 8910
rect 4632 8838 4660 9302
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 8566 4660 8774
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4296 8188 4604 8197
rect 4296 8186 4302 8188
rect 4358 8186 4382 8188
rect 4438 8186 4462 8188
rect 4518 8186 4542 8188
rect 4598 8186 4604 8188
rect 4358 8134 4360 8186
rect 4540 8134 4542 8186
rect 4296 8132 4302 8134
rect 4358 8132 4382 8134
rect 4438 8132 4462 8134
rect 4518 8132 4542 8134
rect 4598 8132 4604 8134
rect 4296 8123 4604 8132
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4172 7002 4200 7278
rect 4296 7100 4604 7109
rect 4296 7098 4302 7100
rect 4358 7098 4382 7100
rect 4438 7098 4462 7100
rect 4518 7098 4542 7100
rect 4598 7098 4604 7100
rect 4358 7046 4360 7098
rect 4540 7046 4542 7098
rect 4296 7044 4302 7046
rect 4358 7044 4382 7046
rect 4438 7044 4462 7046
rect 4518 7044 4542 7046
rect 4598 7044 4604 7046
rect 4296 7035 4604 7044
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3988 6458 4016 6666
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3988 6322 4016 6394
rect 4080 6322 4108 6598
rect 3976 6316 4028 6322
rect 3896 6276 3976 6304
rect 3896 5778 3924 6276
rect 3976 6258 4028 6264
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4706 4016 4966
rect 4080 4758 4108 5510
rect 4172 5302 4200 6054
rect 4296 6012 4604 6021
rect 4296 6010 4302 6012
rect 4358 6010 4382 6012
rect 4438 6010 4462 6012
rect 4518 6010 4542 6012
rect 4598 6010 4604 6012
rect 4358 5958 4360 6010
rect 4540 5958 4542 6010
rect 4296 5956 4302 5958
rect 4358 5956 4382 5958
rect 4438 5956 4462 5958
rect 4518 5956 4542 5958
rect 4598 5956 4604 5958
rect 4296 5947 4604 5956
rect 4632 5710 4660 8502
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 5914 4752 8366
rect 4816 6662 4844 10526
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5184 9178 5212 9998
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4068 4752 4120 4758
rect 3988 4700 4068 4706
rect 3988 4694 4120 4700
rect 3988 4678 4108 4694
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3896 4282 3924 4558
rect 3988 4554 4016 4678
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 4080 4214 4108 4678
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4080 3534 4108 4150
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4172 3126 4200 4966
rect 4296 4924 4604 4933
rect 4296 4922 4302 4924
rect 4358 4922 4382 4924
rect 4438 4922 4462 4924
rect 4518 4922 4542 4924
rect 4598 4922 4604 4924
rect 4358 4870 4360 4922
rect 4540 4870 4542 4922
rect 4296 4868 4302 4870
rect 4358 4868 4382 4870
rect 4438 4868 4462 4870
rect 4518 4868 4542 4870
rect 4598 4868 4604 4870
rect 4296 4859 4604 4868
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 3942 4384 4422
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4296 3836 4604 3845
rect 4296 3834 4302 3836
rect 4358 3834 4382 3836
rect 4438 3834 4462 3836
rect 4518 3834 4542 3836
rect 4598 3834 4604 3836
rect 4358 3782 4360 3834
rect 4540 3782 4542 3834
rect 4296 3780 4302 3782
rect 4358 3780 4382 3782
rect 4438 3780 4462 3782
rect 4518 3780 4542 3782
rect 4598 3780 4604 3782
rect 4296 3771 4604 3780
rect 4632 3738 4660 5034
rect 4724 3942 4752 5578
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4816 3738 4844 6598
rect 4908 6118 4936 7142
rect 5000 6730 5028 9046
rect 5276 7886 5304 9522
rect 5264 7880 5316 7886
rect 5184 7828 5264 7834
rect 5184 7822 5316 7828
rect 5184 7806 5304 7822
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 5184 6662 5212 7806
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6798 5304 7142
rect 5368 7002 5396 7686
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 5302 4936 5510
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 5368 5234 5396 6598
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5000 4690 5028 5170
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5000 4282 5028 4626
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5184 4214 5212 4558
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 5184 3534 5212 4150
rect 5460 3738 5488 11766
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6380 11286 6408 11698
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 10266 5580 10406
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5644 10146 5672 10950
rect 5552 10130 5672 10146
rect 5540 10124 5672 10130
rect 5592 10118 5672 10124
rect 5540 10066 5592 10072
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8634 5580 8910
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 7410 5672 8298
rect 5736 7410 5764 8502
rect 5828 8090 5856 8842
rect 6472 8566 6500 11698
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6564 11082 6592 11630
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6656 10606 6684 12106
rect 7024 11830 7052 12396
rect 7104 12378 7156 12384
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 7392 11286 7420 13942
rect 7484 13938 7512 14758
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 14074 7604 14214
rect 7642 14172 7950 14181
rect 7642 14170 7648 14172
rect 7704 14170 7728 14172
rect 7784 14170 7808 14172
rect 7864 14170 7888 14172
rect 7944 14170 7950 14172
rect 7704 14118 7706 14170
rect 7886 14118 7888 14170
rect 7642 14116 7648 14118
rect 7704 14116 7728 14118
rect 7784 14116 7808 14118
rect 7864 14116 7888 14118
rect 7944 14116 7950 14118
rect 7642 14107 7950 14116
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 8036 13190 8064 14282
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11830 7512 12038
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7576 11694 7604 13126
rect 7642 13084 7950 13093
rect 7642 13082 7648 13084
rect 7704 13082 7728 13084
rect 7784 13082 7808 13084
rect 7864 13082 7888 13084
rect 7944 13082 7950 13084
rect 7704 13030 7706 13082
rect 7886 13030 7888 13082
rect 7642 13028 7648 13030
rect 7704 13028 7728 13030
rect 7784 13028 7808 13030
rect 7864 13028 7888 13030
rect 7944 13028 7950 13030
rect 7642 13019 7950 13028
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7668 12306 7696 12718
rect 8128 12434 8156 16458
rect 8220 15162 8248 18702
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8312 17882 8340 18294
rect 8588 17882 8616 19502
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16046 8340 17002
rect 8680 16046 8708 18158
rect 8772 16794 8800 20266
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8864 17678 8892 20198
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9140 19310 9168 19654
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9232 19174 9260 20810
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 18358 9260 18566
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 16998 8892 17478
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8864 16794 8892 16934
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8864 16130 8892 16730
rect 8956 16658 8984 17138
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8772 16114 8892 16130
rect 8760 16108 8892 16114
rect 8812 16102 8892 16108
rect 8760 16050 8812 16056
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8312 15366 8340 15642
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8220 12442 8248 15098
rect 8312 14482 8340 15302
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8312 13326 8340 13466
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8036 12406 8156 12434
rect 8208 12436 8260 12442
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7642 11996 7950 12005
rect 7642 11994 7648 11996
rect 7704 11994 7728 11996
rect 7784 11994 7808 11996
rect 7864 11994 7888 11996
rect 7944 11994 7950 11996
rect 7704 11942 7706 11994
rect 7886 11942 7888 11994
rect 7642 11940 7648 11942
rect 7704 11940 7728 11942
rect 7784 11940 7808 11942
rect 7864 11940 7888 11942
rect 7944 11940 7950 11942
rect 7642 11931 7950 11940
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7944 11778 7972 11834
rect 8036 11778 8064 12406
rect 8208 12378 8260 12384
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7852 11370 7880 11766
rect 7944 11750 8064 11778
rect 8128 11744 8156 12242
rect 8312 12170 8340 13262
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8128 11716 8248 11744
rect 8220 11676 8248 11716
rect 8300 11688 8352 11694
rect 8220 11648 8300 11676
rect 8300 11630 8352 11636
rect 7760 11354 7880 11370
rect 7748 11348 7880 11354
rect 7800 11342 7880 11348
rect 7748 11290 7800 11296
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 8404 11218 8432 12378
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9654 6592 9998
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6552 8900 6604 8906
rect 6552 8842 6604 8848
rect 6564 8634 6592 8842
rect 6840 8838 6868 11086
rect 7012 11008 7064 11014
rect 6932 10968 7012 10996
rect 6932 10742 6960 10968
rect 7012 10950 7064 10956
rect 8404 10962 8432 11154
rect 8496 11082 8524 14962
rect 8680 14958 8708 15982
rect 8864 15706 8892 16102
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8588 12170 8616 13466
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8588 11150 8616 12106
rect 8864 11830 8892 15642
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8404 10934 8616 10962
rect 7642 10908 7950 10917
rect 7642 10906 7648 10908
rect 7704 10906 7728 10908
rect 7784 10906 7808 10908
rect 7864 10906 7888 10908
rect 7944 10906 7950 10908
rect 7704 10854 7706 10906
rect 7886 10854 7888 10906
rect 7642 10852 7648 10854
rect 7704 10852 7728 10854
rect 7784 10852 7808 10854
rect 7864 10852 7888 10854
rect 7944 10852 7950 10854
rect 7642 10843 7950 10852
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6932 9926 6960 10678
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6840 8650 6868 8774
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6748 8622 6868 8650
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5552 5166 5580 6190
rect 5920 5778 5948 8366
rect 6748 7954 6776 8622
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5370 5672 5646
rect 6012 5642 6040 6190
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 6196 5234 6224 7822
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6288 5914 6316 7346
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6564 6730 6592 7278
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6840 5574 6868 8502
rect 6932 8498 6960 9862
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7024 8498 7052 9522
rect 7208 8498 7236 9522
rect 7392 9178 7420 9930
rect 7484 9450 7512 10066
rect 7668 10062 7696 10406
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7642 9820 7950 9829
rect 7642 9818 7648 9820
rect 7704 9818 7728 9820
rect 7784 9818 7808 9820
rect 7864 9818 7888 9820
rect 7944 9818 7950 9820
rect 7704 9766 7706 9818
rect 7886 9766 7888 9818
rect 7642 9764 7648 9766
rect 7704 9764 7728 9766
rect 7784 9764 7808 9766
rect 7864 9764 7888 9766
rect 7944 9764 7950 9766
rect 7642 9755 7950 9764
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7300 8498 7328 9114
rect 7642 8732 7950 8741
rect 7642 8730 7648 8732
rect 7704 8730 7728 8732
rect 7784 8730 7808 8732
rect 7864 8730 7888 8732
rect 7944 8730 7950 8732
rect 7704 8678 7706 8730
rect 7886 8678 7888 8730
rect 7642 8676 7648 8678
rect 7704 8676 7728 8678
rect 7784 8676 7808 8678
rect 7864 8676 7888 8678
rect 7944 8676 7950 8678
rect 7642 8667 7950 8676
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7024 7410 7052 8434
rect 7208 8090 7236 8434
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6932 6322 6960 7210
rect 7024 6914 7052 7346
rect 7024 6886 7144 6914
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4826 5580 5102
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6840 3738 6868 5510
rect 7116 5166 7144 6886
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 5370 7236 6734
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7392 4146 7420 8026
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7484 6458 7512 7346
rect 7576 6798 7604 7754
rect 7642 7644 7950 7653
rect 7642 7642 7648 7644
rect 7704 7642 7728 7644
rect 7784 7642 7808 7644
rect 7864 7642 7888 7644
rect 7944 7642 7950 7644
rect 7704 7590 7706 7642
rect 7886 7590 7888 7642
rect 7642 7588 7648 7590
rect 7704 7588 7728 7590
rect 7784 7588 7808 7590
rect 7864 7588 7888 7590
rect 7944 7588 7950 7590
rect 7642 7579 7950 7588
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7484 5234 7512 6394
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7576 4622 7604 6734
rect 7642 6556 7950 6565
rect 7642 6554 7648 6556
rect 7704 6554 7728 6556
rect 7784 6554 7808 6556
rect 7864 6554 7888 6556
rect 7944 6554 7950 6556
rect 7704 6502 7706 6554
rect 7886 6502 7888 6554
rect 7642 6500 7648 6502
rect 7704 6500 7728 6502
rect 7784 6500 7808 6502
rect 7864 6500 7888 6502
rect 7944 6500 7950 6502
rect 7642 6491 7950 6500
rect 8128 6458 8156 10610
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8220 6866 8248 10474
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8404 9654 8432 9930
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8496 9450 8524 9930
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5914 8064 6190
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8128 5710 8156 6394
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8220 5574 8248 6802
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7642 5468 7950 5477
rect 7642 5466 7648 5468
rect 7704 5466 7728 5468
rect 7784 5466 7808 5468
rect 7864 5466 7888 5468
rect 7944 5466 7950 5468
rect 7704 5414 7706 5466
rect 7886 5414 7888 5466
rect 7642 5412 7648 5414
rect 7704 5412 7728 5414
rect 7784 5412 7808 5414
rect 7864 5412 7888 5414
rect 7944 5412 7950 5414
rect 7642 5403 7950 5412
rect 8312 5370 8340 6326
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 4690 7696 5170
rect 8588 4826 8616 10934
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 8974 8800 9522
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8362 8800 8910
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8772 7886 8800 8298
rect 8956 8090 8984 16594
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 15026 9076 15846
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9048 14006 9076 14758
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 9140 13818 9168 14010
rect 9048 13790 9168 13818
rect 9048 12170 9076 13790
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13530 9168 13670
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 13410 9260 15438
rect 9140 13382 9260 13410
rect 9140 12374 9168 13382
rect 9324 13297 9352 21966
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9600 19718 9628 20402
rect 9692 20398 9720 20742
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 18698 9628 19654
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18426 9628 18634
rect 9692 18426 9720 18702
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9416 17202 9444 17750
rect 9508 17746 9536 18022
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16590 9536 16934
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 14414 9536 16526
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9508 14074 9536 14350
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9310 13288 9366 13297
rect 9310 13223 9366 13232
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11286 9260 11494
rect 9324 11354 9352 12718
rect 9416 12170 9444 13194
rect 9600 12764 9628 18158
rect 9784 18086 9812 23462
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10060 22710 10088 22918
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 10060 21146 10088 21490
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9968 19514 9996 19790
rect 10152 19786 10180 20402
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10336 19854 10364 20266
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10152 19446 10180 19722
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10336 18970 10364 19790
rect 10428 19718 10456 20402
rect 10612 20058 10640 24142
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 10988 23420 11296 23429
rect 10988 23418 10994 23420
rect 11050 23418 11074 23420
rect 11130 23418 11154 23420
rect 11210 23418 11234 23420
rect 11290 23418 11296 23420
rect 11050 23366 11052 23418
rect 11232 23366 11234 23418
rect 10988 23364 10994 23366
rect 11050 23364 11074 23366
rect 11130 23364 11154 23366
rect 11210 23364 11234 23366
rect 11290 23364 11296 23366
rect 10988 23355 11296 23364
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11164 22778 11192 23054
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 10988 22332 11296 22341
rect 10988 22330 10994 22332
rect 11050 22330 11074 22332
rect 11130 22330 11154 22332
rect 11210 22330 11234 22332
rect 11290 22330 11296 22332
rect 11050 22278 11052 22330
rect 11232 22278 11234 22330
rect 10988 22276 10994 22278
rect 11050 22276 11074 22278
rect 11130 22276 11154 22278
rect 11210 22276 11234 22278
rect 11290 22276 11296 22278
rect 10988 22267 11296 22276
rect 11440 22250 11468 23122
rect 11348 22234 11468 22250
rect 11336 22228 11468 22234
rect 11388 22222 11468 22228
rect 11336 22170 11388 22176
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 10988 21244 11296 21253
rect 10988 21242 10994 21244
rect 11050 21242 11074 21244
rect 11130 21242 11154 21244
rect 11210 21242 11234 21244
rect 11290 21242 11296 21244
rect 11050 21190 11052 21242
rect 11232 21190 11234 21242
rect 10988 21188 10994 21190
rect 11050 21188 11074 21190
rect 11130 21188 11154 21190
rect 11210 21188 11234 21190
rect 11290 21188 11296 21190
rect 10988 21179 11296 21188
rect 11348 21146 11376 21422
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11440 21010 11468 22222
rect 11532 22094 11560 24074
rect 11624 22778 11652 24142
rect 12084 23730 12112 24346
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11992 23118 12020 23598
rect 12176 23594 12204 24754
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 12176 23118 12204 23530
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 11532 22066 11652 22094
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20602 11100 20810
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10988 20156 11296 20165
rect 10988 20154 10994 20156
rect 11050 20154 11074 20156
rect 11130 20154 11154 20156
rect 11210 20154 11234 20156
rect 11290 20154 11296 20156
rect 11050 20102 11052 20154
rect 11232 20102 11234 20154
rect 10988 20100 10994 20102
rect 11050 20100 11074 20102
rect 11130 20100 11154 20102
rect 11210 20100 11234 20102
rect 11290 20100 11296 20102
rect 10988 20091 11296 20100
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 11440 19922 11468 20946
rect 11624 20534 11652 22066
rect 12176 21554 12204 22578
rect 12268 21894 12296 23462
rect 12452 22710 12480 25162
rect 12544 24818 12572 26250
rect 12636 26246 12664 28200
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12728 25498 12756 25842
rect 12716 25492 12768 25498
rect 12716 25434 12768 25440
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12452 21962 12480 22510
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12176 21078 12204 21490
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11532 20262 11560 20402
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10428 18426 10456 19654
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9680 17672 9732 17678
rect 9732 17632 9812 17660
rect 9680 17614 9732 17620
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9692 15366 9720 16594
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 15094 9720 15302
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9680 12776 9732 12782
rect 9600 12736 9680 12764
rect 9680 12718 9732 12724
rect 9784 12646 9812 17632
rect 9968 17134 9996 17682
rect 10520 17678 10548 19654
rect 10988 19068 11296 19077
rect 10988 19066 10994 19068
rect 11050 19066 11074 19068
rect 11130 19066 11154 19068
rect 11210 19066 11234 19068
rect 11290 19066 11296 19068
rect 11050 19014 11052 19066
rect 11232 19014 11234 19066
rect 10988 19012 10994 19014
rect 11050 19012 11074 19014
rect 11130 19012 11154 19014
rect 11210 19012 11234 19014
rect 11290 19012 11296 19014
rect 10988 19003 11296 19012
rect 11348 18698 11376 19722
rect 11440 19514 11468 19858
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11532 19378 11560 20198
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 11440 18834 11468 19246
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 10988 17980 11296 17989
rect 10988 17978 10994 17980
rect 11050 17978 11074 17980
rect 11130 17978 11154 17980
rect 11210 17978 11234 17980
rect 11290 17978 11296 17980
rect 11050 17926 11052 17978
rect 11232 17926 11234 17978
rect 10988 17924 10994 17926
rect 11050 17924 11074 17926
rect 11130 17924 11154 17926
rect 11210 17924 11234 17926
rect 11290 17924 11296 17926
rect 10988 17915 11296 17924
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9968 16658 9996 17070
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10060 16590 10088 17274
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10508 17060 10560 17066
rect 10508 17002 10560 17008
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 15978 10088 16526
rect 10520 16046 10548 17002
rect 10612 16794 10640 17138
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10704 16658 10732 17206
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 10060 14362 10088 15914
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10428 14414 10456 14758
rect 10416 14408 10468 14414
rect 9876 13530 9904 14350
rect 10060 14334 10180 14362
rect 10416 14350 10468 14356
rect 10520 14346 10548 15846
rect 10612 15502 10640 16186
rect 10704 16182 10732 16594
rect 10796 16454 10824 17274
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10704 15570 10732 16118
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10704 15162 10732 15506
rect 10796 15502 10824 15914
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10796 15026 10824 15098
rect 10888 15026 10916 17478
rect 11440 17270 11468 18770
rect 11532 17678 11560 19314
rect 11716 18834 11744 20538
rect 11808 20534 11836 20742
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 12176 19786 12204 20266
rect 12268 19990 12296 21830
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 20942 12388 21354
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12636 20602 12664 22986
rect 12728 22642 12756 25434
rect 13280 25294 13308 26250
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13648 24954 13676 26318
rect 13832 25974 13860 26318
rect 14334 26140 14642 26149
rect 14334 26138 14340 26140
rect 14396 26138 14420 26140
rect 14476 26138 14500 26140
rect 14556 26138 14580 26140
rect 14636 26138 14642 26140
rect 14396 26086 14398 26138
rect 14578 26086 14580 26138
rect 14334 26084 14340 26086
rect 14396 26084 14420 26086
rect 14476 26084 14500 26086
rect 14556 26084 14580 26086
rect 14636 26084 14642 26086
rect 14334 26075 14642 26084
rect 13820 25968 13872 25974
rect 13820 25910 13872 25916
rect 14096 25968 14148 25974
rect 14096 25910 14148 25916
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13188 23186 13216 24074
rect 13648 23866 13676 24890
rect 14016 24682 14044 25094
rect 14108 24818 14136 25910
rect 15304 25838 15332 26386
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 14188 25832 14240 25838
rect 14188 25774 14240 25780
rect 15016 25832 15068 25838
rect 15016 25774 15068 25780
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14004 24676 14056 24682
rect 14004 24618 14056 24624
rect 14200 24410 14228 25774
rect 14924 25220 14976 25226
rect 14924 25162 14976 25168
rect 14334 25052 14642 25061
rect 14334 25050 14340 25052
rect 14396 25050 14420 25052
rect 14476 25050 14500 25052
rect 14556 25050 14580 25052
rect 14636 25050 14642 25052
rect 14396 24998 14398 25050
rect 14578 24998 14580 25050
rect 14334 24996 14340 24998
rect 14396 24996 14420 24998
rect 14476 24996 14500 24998
rect 14556 24996 14580 24998
rect 14636 24996 14642 24998
rect 14334 24987 14642 24996
rect 14936 24886 14964 25162
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 15028 24206 15056 25774
rect 15304 25158 15332 25774
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15120 24410 15148 25094
rect 15488 24750 15516 25638
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15580 24750 15608 25230
rect 15764 24954 15792 26318
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15120 24206 15148 24346
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 14334 23964 14642 23973
rect 14334 23962 14340 23964
rect 14396 23962 14420 23964
rect 14476 23962 14500 23964
rect 14556 23962 14580 23964
rect 14636 23962 14642 23964
rect 14396 23910 14398 23962
rect 14578 23910 14580 23962
rect 14334 23908 14340 23910
rect 14396 23908 14420 23910
rect 14476 23908 14500 23910
rect 14556 23908 14580 23910
rect 14636 23908 14642 23910
rect 14334 23899 14642 23908
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13176 23180 13228 23186
rect 13176 23122 13228 23128
rect 13648 23118 13676 23802
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 15028 23050 15056 24142
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15016 23044 15068 23050
rect 15016 22986 15068 22992
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22710 13768 22918
rect 14334 22876 14642 22885
rect 14334 22874 14340 22876
rect 14396 22874 14420 22876
rect 14476 22874 14500 22876
rect 14556 22874 14580 22876
rect 14636 22874 14642 22876
rect 14396 22822 14398 22874
rect 14578 22822 14580 22874
rect 14334 22820 14340 22822
rect 14396 22820 14420 22822
rect 14476 22820 14500 22822
rect 14556 22820 14580 22822
rect 14636 22820 14642 22822
rect 14334 22811 14642 22820
rect 15212 22778 15240 23054
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 13728 22704 13780 22710
rect 13464 22664 13728 22692
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13096 21146 13124 21490
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 13096 19854 13124 20334
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11808 17882 11836 18634
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11716 16998 11744 17546
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 10988 16892 11296 16901
rect 10988 16890 10994 16892
rect 11050 16890 11074 16892
rect 11130 16890 11154 16892
rect 11210 16890 11234 16892
rect 11290 16890 11296 16892
rect 11050 16838 11052 16890
rect 11232 16838 11234 16890
rect 10988 16836 10994 16838
rect 11050 16836 11074 16838
rect 11130 16836 11154 16838
rect 11210 16836 11234 16838
rect 11290 16836 11296 16838
rect 10988 16827 11296 16836
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16250 11008 16390
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10980 16114 11008 16186
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10988 15804 11296 15813
rect 10988 15802 10994 15804
rect 11050 15802 11074 15804
rect 11130 15802 11154 15804
rect 11210 15802 11234 15804
rect 11290 15802 11296 15804
rect 11050 15750 11052 15802
rect 11232 15750 11234 15802
rect 10988 15748 10994 15750
rect 11050 15748 11074 15750
rect 11130 15748 11154 15750
rect 11210 15748 11234 15750
rect 11290 15748 11296 15750
rect 10988 15739 11296 15748
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10988 14716 11296 14725
rect 10988 14714 10994 14716
rect 11050 14714 11074 14716
rect 11130 14714 11154 14716
rect 11210 14714 11234 14716
rect 11290 14714 11296 14716
rect 11050 14662 11052 14714
rect 11232 14662 11234 14714
rect 10988 14660 10994 14662
rect 11050 14660 11074 14662
rect 11130 14660 11154 14662
rect 11210 14660 11234 14662
rect 11290 14660 11296 14662
rect 10988 14651 11296 14660
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13938 10088 14214
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9508 11150 9536 11222
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9140 10266 9168 11086
rect 9692 10810 9720 11630
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9784 10674 9812 12582
rect 9968 12442 9996 13806
rect 9956 12436 10008 12442
rect 10152 12434 10180 14334
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10612 13938 10640 14282
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10244 12850 10272 13126
rect 10520 12986 10548 13330
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9956 12378 10008 12384
rect 10060 12406 10180 12434
rect 9968 11830 9996 12378
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10060 10674 10088 12406
rect 10244 11762 10272 12582
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10152 10606 10180 11154
rect 10336 11150 10364 12922
rect 10888 12646 10916 13806
rect 10988 13628 11296 13637
rect 10988 13626 10994 13628
rect 11050 13626 11074 13628
rect 11130 13626 11154 13628
rect 11210 13626 11234 13628
rect 11290 13626 11296 13628
rect 11050 13574 11052 13626
rect 11232 13574 11234 13626
rect 10988 13572 10994 13574
rect 11050 13572 11074 13574
rect 11130 13572 11154 13574
rect 11210 13572 11234 13574
rect 11290 13572 11296 13574
rect 10988 13563 11296 13572
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 11898 10456 12106
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10612 11762 10640 12310
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11830 10732 12174
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10796 11642 10824 12038
rect 10888 11762 10916 12582
rect 10988 12540 11296 12549
rect 10988 12538 10994 12540
rect 11050 12538 11074 12540
rect 11130 12538 11154 12540
rect 11210 12538 11234 12540
rect 11290 12538 11296 12540
rect 11050 12486 11052 12538
rect 11232 12486 11234 12538
rect 10988 12484 10994 12486
rect 11050 12484 11074 12486
rect 11130 12484 11154 12486
rect 11210 12484 11234 12486
rect 11290 12484 11296 12486
rect 10988 12475 11296 12484
rect 11348 12306 11376 16458
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 15434 11836 16390
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11428 15428 11480 15434
rect 11796 15428 11848 15434
rect 11480 15388 11560 15416
rect 11428 15370 11480 15376
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10796 11614 10916 11642
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5234 8892 5646
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 9048 4622 9076 7142
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 5302 9168 6734
rect 9232 6458 9260 8502
rect 9692 6914 9720 10542
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9784 9178 9812 10474
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9692 6886 9812 6914
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9784 5114 9812 6886
rect 9876 6254 9904 9998
rect 10060 9722 10088 10406
rect 10152 9722 10180 10542
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10244 9586 10272 9862
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 8906 10180 9318
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10244 8090 10272 8366
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10336 7886 10364 10678
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9518 10732 9930
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10796 9382 10824 9998
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10520 6390 10548 8366
rect 10888 7410 10916 11614
rect 10988 11452 11296 11461
rect 10988 11450 10994 11452
rect 11050 11450 11074 11452
rect 11130 11450 11154 11452
rect 11210 11450 11234 11452
rect 11290 11450 11296 11452
rect 11050 11398 11052 11450
rect 11232 11398 11234 11450
rect 10988 11396 10994 11398
rect 11050 11396 11074 11398
rect 11130 11396 11154 11398
rect 11210 11396 11234 11398
rect 11290 11396 11296 11398
rect 10988 11387 11296 11396
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 10742 11376 10950
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 10988 10364 11296 10373
rect 10988 10362 10994 10364
rect 11050 10362 11074 10364
rect 11130 10362 11154 10364
rect 11210 10362 11234 10364
rect 11290 10362 11296 10364
rect 11050 10310 11052 10362
rect 11232 10310 11234 10362
rect 10988 10308 10994 10310
rect 11050 10308 11074 10310
rect 11130 10308 11154 10310
rect 11210 10308 11234 10310
rect 11290 10308 11296 10310
rect 10988 10299 11296 10308
rect 10988 9276 11296 9285
rect 10988 9274 10994 9276
rect 11050 9274 11074 9276
rect 11130 9274 11154 9276
rect 11210 9274 11234 9276
rect 11290 9274 11296 9276
rect 11050 9222 11052 9274
rect 11232 9222 11234 9274
rect 10988 9220 10994 9222
rect 11050 9220 11074 9222
rect 11130 9220 11154 9222
rect 11210 9220 11234 9222
rect 11290 9220 11296 9222
rect 10988 9211 11296 9220
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8634 11008 8842
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11348 8498 11376 10406
rect 11440 9722 11468 13874
rect 11532 13802 11560 15388
rect 11796 15370 11848 15376
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11624 14482 11652 14758
rect 11716 14618 11744 14758
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11808 14498 11836 15370
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11716 14470 11836 14498
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11716 13190 11744 14470
rect 11900 13920 11928 15438
rect 12084 14346 12112 19314
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18630 12204 19110
rect 12636 18698 12664 19382
rect 13096 18970 13124 19790
rect 13188 19446 13216 20402
rect 13464 19786 13492 22664
rect 13728 22646 13780 22652
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13832 22030 13860 22374
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13740 21350 13768 21898
rect 14334 21788 14642 21797
rect 14334 21786 14340 21788
rect 14396 21786 14420 21788
rect 14476 21786 14500 21788
rect 14556 21786 14580 21788
rect 14636 21786 14642 21788
rect 14396 21734 14398 21786
rect 14578 21734 14580 21786
rect 14334 21732 14340 21734
rect 14396 21732 14420 21734
rect 14476 21732 14500 21734
rect 14556 21732 14580 21734
rect 14636 21732 14642 21734
rect 14334 21723 14642 21732
rect 14936 21418 14964 22442
rect 15212 22234 15240 22714
rect 15304 22642 15332 23054
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 14924 21412 14976 21418
rect 14924 21354 14976 21360
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13556 19854 13584 20402
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 20058 13676 20198
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13740 19854 13768 21286
rect 14936 21010 14964 21354
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 18290 12204 18566
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12636 18222 12664 18634
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12176 14278 12204 14894
rect 12360 14618 12388 17478
rect 12544 15706 12572 18158
rect 12636 17796 12664 18158
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12716 17808 12768 17814
rect 12636 17768 12716 17796
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12176 14074 12204 14214
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12360 13938 12388 14554
rect 12072 13932 12124 13938
rect 11900 13892 12072 13920
rect 12072 13874 12124 13880
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11992 13190 12020 13738
rect 12084 13394 12112 13874
rect 12164 13728 12216 13734
rect 12440 13728 12492 13734
rect 12164 13670 12216 13676
rect 12438 13696 12440 13705
rect 12492 13696 12494 13705
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11704 13184 11756 13190
rect 11888 13184 11940 13190
rect 11704 13126 11756 13132
rect 11886 13152 11888 13161
rect 11980 13184 12032 13190
rect 11940 13152 11942 13161
rect 11980 13126 12032 13132
rect 11886 13087 11942 13096
rect 12084 13025 12112 13330
rect 12176 13326 12204 13670
rect 12438 13631 12494 13640
rect 12438 13560 12494 13569
rect 12438 13495 12440 13504
rect 12492 13495 12494 13504
rect 12440 13466 12492 13472
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12070 13016 12126 13025
rect 11520 12980 11572 12986
rect 12070 12951 12126 12960
rect 11520 12922 11572 12928
rect 11532 11694 11560 12922
rect 12544 12850 12572 15642
rect 12636 15638 12664 17768
rect 12716 17750 12768 17756
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12728 17105 12756 17546
rect 12714 17096 12770 17105
rect 12714 17031 12770 17040
rect 12820 16250 12848 17614
rect 13096 17270 13124 17818
rect 13280 17746 13308 19654
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13648 18290 13676 18566
rect 13740 18426 13768 19790
rect 14108 19786 14136 20742
rect 14200 20602 14228 20878
rect 14334 20700 14642 20709
rect 14334 20698 14340 20700
rect 14396 20698 14420 20700
rect 14476 20698 14500 20700
rect 14556 20698 14580 20700
rect 14636 20698 14642 20700
rect 14396 20646 14398 20698
rect 14578 20646 14580 20698
rect 14334 20644 14340 20646
rect 14396 20644 14420 20646
rect 14476 20644 14500 20646
rect 14556 20644 14580 20646
rect 14636 20644 14642 20646
rect 14334 20635 14642 20644
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14936 20398 14964 20946
rect 15212 20942 15240 21626
rect 15396 21350 15424 23462
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15488 21486 15516 23122
rect 15580 22642 15608 24686
rect 15764 24206 15792 24890
rect 16132 24886 16160 26250
rect 16224 26246 16252 28200
rect 17680 26684 17988 26693
rect 17680 26682 17686 26684
rect 17742 26682 17766 26684
rect 17822 26682 17846 26684
rect 17902 26682 17926 26684
rect 17982 26682 17988 26684
rect 17742 26630 17744 26682
rect 17924 26630 17926 26682
rect 17680 26628 17686 26630
rect 17742 26628 17766 26630
rect 17822 26628 17846 26630
rect 17902 26628 17926 26630
rect 17982 26628 17988 26630
rect 17680 26619 17988 26628
rect 19812 26586 19840 28200
rect 23400 26602 23428 28200
rect 24372 26684 24680 26693
rect 24372 26682 24378 26684
rect 24434 26682 24458 26684
rect 24514 26682 24538 26684
rect 24594 26682 24618 26684
rect 24674 26682 24680 26684
rect 24434 26630 24436 26682
rect 24616 26630 24618 26682
rect 24372 26628 24378 26630
rect 24434 26628 24458 26630
rect 24514 26628 24538 26630
rect 24594 26628 24618 26630
rect 24674 26628 24680 26630
rect 24372 26619 24680 26628
rect 23400 26586 23520 26602
rect 26988 26586 27016 28200
rect 19800 26580 19852 26586
rect 23400 26580 23532 26586
rect 23400 26574 23480 26580
rect 19800 26522 19852 26528
rect 23480 26522 23532 26528
rect 26976 26580 27028 26586
rect 26976 26522 27028 26528
rect 16856 26376 16908 26382
rect 16856 26318 16908 26324
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16868 25770 16896 26318
rect 19352 25906 19380 26318
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 17316 25900 17368 25906
rect 17316 25842 17368 25848
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 16856 25764 16908 25770
rect 16856 25706 16908 25712
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16592 24274 16620 25162
rect 17144 24274 17172 25638
rect 17328 25158 17356 25842
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 17680 25596 17988 25605
rect 17680 25594 17686 25596
rect 17742 25594 17766 25596
rect 17822 25594 17846 25596
rect 17902 25594 17926 25596
rect 17982 25594 17988 25596
rect 17742 25542 17744 25594
rect 17924 25542 17926 25594
rect 17680 25540 17686 25542
rect 17742 25540 17766 25542
rect 17822 25540 17846 25542
rect 17902 25540 17926 25542
rect 17982 25540 17988 25542
rect 17680 25531 17988 25540
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17316 25152 17368 25158
rect 17316 25094 17368 25100
rect 17328 24818 17356 25094
rect 17420 24886 17448 25230
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 18328 25220 18380 25226
rect 18328 25162 18380 25168
rect 17604 24886 17632 25162
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 17408 24880 17460 24886
rect 17408 24822 17460 24828
rect 17592 24880 17644 24886
rect 17592 24822 17644 24828
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 16316 22574 16344 22986
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 15856 21690 15884 22510
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16224 21690 16252 21966
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16316 21622 16344 21830
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15856 21010 15884 21286
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 20602 16068 20878
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14334 19612 14642 19621
rect 14334 19610 14340 19612
rect 14396 19610 14420 19612
rect 14476 19610 14500 19612
rect 14556 19610 14580 19612
rect 14636 19610 14642 19612
rect 14396 19558 14398 19610
rect 14578 19558 14580 19610
rect 14334 19556 14340 19558
rect 14396 19556 14420 19558
rect 14476 19556 14500 19558
rect 14556 19556 14580 19558
rect 14636 19556 14642 19558
rect 14334 19547 14642 19556
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12912 14090 12940 17206
rect 13280 16794 13308 17682
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13464 17270 13492 17546
rect 13740 17338 13768 17546
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13832 17134 13860 18090
rect 14016 17678 14044 18702
rect 14200 18426 14228 19314
rect 14936 18834 14964 20334
rect 15580 20058 15608 20402
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15108 18896 15160 18902
rect 15108 18838 15160 18844
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14334 18524 14642 18533
rect 14334 18522 14340 18524
rect 14396 18522 14420 18524
rect 14476 18522 14500 18524
rect 14556 18522 14580 18524
rect 14636 18522 14642 18524
rect 14396 18470 14398 18522
rect 14578 18470 14580 18522
rect 14334 18468 14340 18470
rect 14396 18468 14420 18470
rect 14476 18468 14500 18470
rect 14556 18468 14580 18470
rect 14636 18468 14642 18470
rect 14334 18459 14642 18468
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13910 17096 13966 17105
rect 13910 17031 13912 17040
rect 13964 17031 13966 17040
rect 13912 17002 13964 17008
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13004 14346 13216 14362
rect 12992 14340 13216 14346
rect 13044 14334 13216 14340
rect 12992 14282 13044 14288
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12820 14062 12940 14090
rect 12820 13938 12848 14062
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13530 12664 13670
rect 12714 13560 12770 13569
rect 12624 13524 12676 13530
rect 12714 13495 12716 13504
rect 12624 13466 12676 13472
rect 12768 13495 12770 13504
rect 12716 13466 12768 13472
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12452 12730 12480 12786
rect 12716 12776 12768 12782
rect 12452 12702 12664 12730
rect 12820 12764 12848 13874
rect 12768 12736 12848 12764
rect 12716 12718 12768 12724
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 10198 11560 11630
rect 11624 11626 11652 12242
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11716 10674 11744 12038
rect 11808 11898 11836 12106
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 10988 8188 11296 8197
rect 10988 8186 10994 8188
rect 11050 8186 11074 8188
rect 11130 8186 11154 8188
rect 11210 8186 11234 8188
rect 11290 8186 11296 8188
rect 11050 8134 11052 8186
rect 11232 8134 11234 8186
rect 10988 8132 10994 8134
rect 11050 8132 11074 8134
rect 11130 8132 11154 8134
rect 11210 8132 11234 8134
rect 11290 8132 11296 8134
rect 10988 8123 11296 8132
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 10988 7100 11296 7109
rect 10988 7098 10994 7100
rect 11050 7098 11074 7100
rect 11130 7098 11154 7100
rect 11210 7098 11234 7100
rect 11290 7098 11296 7100
rect 11050 7046 11052 7098
rect 11232 7046 11234 7098
rect 10988 7044 10994 7046
rect 11050 7044 11074 7046
rect 11130 7044 11154 7046
rect 11210 7044 11234 7046
rect 11290 7044 11296 7046
rect 10988 7035 11296 7044
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9968 5710 9996 6258
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10244 5710 10272 6190
rect 10612 5778 10640 6666
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10796 5710 10824 6802
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10980 6322 11008 6666
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10988 6012 11296 6021
rect 10988 6010 10994 6012
rect 11050 6010 11074 6012
rect 11130 6010 11154 6012
rect 11210 6010 11234 6012
rect 11290 6010 11296 6012
rect 11050 5958 11052 6010
rect 11232 5958 11234 6010
rect 10988 5956 10994 5958
rect 11050 5956 11074 5958
rect 11130 5956 11154 5958
rect 11210 5956 11234 5958
rect 11290 5956 11296 5958
rect 10988 5947 11296 5956
rect 11348 5778 11376 7142
rect 11440 6662 11468 8910
rect 11532 8906 11560 10134
rect 11808 9042 11836 11834
rect 12360 11762 12388 12582
rect 12452 11830 12480 12582
rect 12636 12170 12664 12702
rect 12912 12617 12940 13874
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 12646 13032 13670
rect 13096 13258 13124 14214
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13188 12850 13216 14334
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 12992 12640 13044 12646
rect 12898 12608 12954 12617
rect 12992 12582 13044 12588
rect 12898 12543 12954 12552
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 11992 10810 12020 11698
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10810 12480 10950
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12544 10674 12572 12038
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9042 11928 9318
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11624 6322 11652 8366
rect 12084 7410 12112 8910
rect 12176 7954 12204 10542
rect 12728 10266 12756 11018
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12728 9450 12756 9658
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12728 7954 12756 9386
rect 12820 9178 12848 10202
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12912 8566 12940 12543
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7546 12940 7686
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13004 7478 13032 10406
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 9968 5234 9996 5646
rect 10796 5234 10824 5646
rect 11716 5234 11744 6394
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 5370 11836 5578
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11900 5234 11928 6598
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11992 5302 12020 6190
rect 12544 5370 12572 6870
rect 13096 6866 13124 9998
rect 13188 8634 13216 12038
rect 13280 9926 13308 16730
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13464 15434 13492 16390
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13556 15026 13584 15914
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 14074 13492 14418
rect 13648 14414 13676 16390
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13464 13258 13492 14010
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13464 12782 13492 13194
rect 13556 12986 13584 13194
rect 13648 13002 13676 14350
rect 13740 13462 13768 16526
rect 14016 14618 14044 17614
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14108 15434 14136 17478
rect 14200 16182 14228 18362
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14334 17436 14642 17445
rect 14334 17434 14340 17436
rect 14396 17434 14420 17436
rect 14476 17434 14500 17436
rect 14556 17434 14580 17436
rect 14636 17434 14642 17436
rect 14396 17382 14398 17434
rect 14578 17382 14580 17434
rect 14334 17380 14340 17382
rect 14396 17380 14420 17382
rect 14476 17380 14500 17382
rect 14556 17380 14580 17382
rect 14636 17380 14642 17382
rect 14334 17371 14642 17380
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14568 16794 14596 17138
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16794 14688 16934
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14334 16348 14642 16357
rect 14334 16346 14340 16348
rect 14396 16346 14420 16348
rect 14476 16346 14500 16348
rect 14556 16346 14580 16348
rect 14636 16346 14642 16348
rect 14396 16294 14398 16346
rect 14578 16294 14580 16346
rect 14334 16292 14340 16294
rect 14396 16292 14420 16294
rect 14476 16292 14500 16294
rect 14556 16292 14580 16294
rect 14636 16292 14642 16294
rect 14334 16283 14642 16292
rect 14752 16182 14780 18022
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14188 16176 14240 16182
rect 14188 16118 14240 16124
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14738 16008 14794 16017
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14016 13870 14044 14554
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13726 13016 13782 13025
rect 13544 12980 13596 12986
rect 13648 12974 13726 13002
rect 13726 12951 13782 12960
rect 13544 12922 13596 12928
rect 13542 12880 13598 12889
rect 13740 12850 13768 12951
rect 13542 12815 13544 12824
rect 13596 12815 13598 12824
rect 13728 12844 13780 12850
rect 13544 12786 13596 12792
rect 13728 12786 13780 12792
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11014 13676 12038
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10198 13676 10950
rect 13740 10266 13768 12786
rect 13832 12374 13860 13806
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14108 13705 14136 13738
rect 14094 13696 14150 13705
rect 14094 13631 14150 13640
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12434 13952 13330
rect 14002 13152 14058 13161
rect 14002 13087 14058 13096
rect 14016 12986 14044 13087
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13924 12406 14044 12434
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 11762 13860 12310
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13924 10810 13952 12174
rect 14016 11694 14044 12406
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14108 11014 14136 13398
rect 14200 13326 14228 15982
rect 14738 15943 14794 15952
rect 14334 15260 14642 15269
rect 14334 15258 14340 15260
rect 14396 15258 14420 15260
rect 14476 15258 14500 15260
rect 14556 15258 14580 15260
rect 14636 15258 14642 15260
rect 14396 15206 14398 15258
rect 14578 15206 14580 15258
rect 14334 15204 14340 15206
rect 14396 15204 14420 15206
rect 14476 15204 14500 15206
rect 14556 15204 14580 15206
rect 14636 15204 14642 15206
rect 14334 15195 14642 15204
rect 14334 14172 14642 14181
rect 14334 14170 14340 14172
rect 14396 14170 14420 14172
rect 14476 14170 14500 14172
rect 14556 14170 14580 14172
rect 14636 14170 14642 14172
rect 14396 14118 14398 14170
rect 14578 14118 14580 14170
rect 14334 14116 14340 14118
rect 14396 14116 14420 14118
rect 14476 14116 14500 14118
rect 14556 14116 14580 14118
rect 14636 14116 14642 14118
rect 14334 14107 14642 14116
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14292 13258 14320 14010
rect 14752 13954 14780 15943
rect 14844 15502 14872 16662
rect 14936 16561 14964 17546
rect 15016 16584 15068 16590
rect 14922 16552 14978 16561
rect 15016 16526 15068 16532
rect 14922 16487 14978 16496
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14660 13926 14780 13954
rect 14660 13802 14688 13926
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14660 13190 14688 13738
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14200 12918 14228 13126
rect 14334 13084 14642 13093
rect 14334 13082 14340 13084
rect 14396 13082 14420 13084
rect 14476 13082 14500 13084
rect 14556 13082 14580 13084
rect 14636 13082 14642 13084
rect 14396 13030 14398 13082
rect 14578 13030 14580 13082
rect 14334 13028 14340 13030
rect 14396 13028 14420 13030
rect 14476 13028 14500 13030
rect 14556 13028 14580 13030
rect 14636 13028 14642 13030
rect 14334 13019 14642 13028
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12617 14596 12718
rect 14554 12608 14610 12617
rect 14554 12543 14610 12552
rect 14752 12306 14780 13806
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14334 11996 14642 12005
rect 14334 11994 14340 11996
rect 14396 11994 14420 11996
rect 14476 11994 14500 11996
rect 14556 11994 14580 11996
rect 14636 11994 14642 11996
rect 14396 11942 14398 11994
rect 14578 11942 14580 11994
rect 14334 11940 14340 11942
rect 14396 11940 14420 11942
rect 14476 11940 14500 11942
rect 14556 11940 14580 11942
rect 14636 11940 14642 11942
rect 14334 11931 14642 11940
rect 14936 11830 14964 16390
rect 15028 14414 15056 16526
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15028 12918 15056 14350
rect 15120 14090 15148 18838
rect 15212 18222 15240 19654
rect 15856 19446 15884 19654
rect 15948 19446 15976 20198
rect 16040 20058 16068 20402
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15936 19440 15988 19446
rect 15936 19382 15988 19388
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15212 17338 15240 18158
rect 15396 17882 15424 19246
rect 15856 18970 15884 19382
rect 16132 19174 16160 20742
rect 16868 19514 16896 23666
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 20942 17080 22918
rect 17236 22574 17264 23054
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 17328 21026 17356 24754
rect 17680 24508 17988 24517
rect 17680 24506 17686 24508
rect 17742 24506 17766 24508
rect 17822 24506 17846 24508
rect 17902 24506 17926 24508
rect 17982 24506 17988 24508
rect 17742 24454 17744 24506
rect 17924 24454 17926 24506
rect 17680 24452 17686 24454
rect 17742 24452 17766 24454
rect 17822 24452 17846 24454
rect 17902 24452 17926 24454
rect 17982 24452 17988 24454
rect 17680 24443 17988 24452
rect 18064 24274 18092 25094
rect 18340 24818 18368 25162
rect 18616 24886 18644 25638
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 17680 23420 17988 23429
rect 17680 23418 17686 23420
rect 17742 23418 17766 23420
rect 17822 23418 17846 23420
rect 17902 23418 17926 23420
rect 17982 23418 17988 23420
rect 17742 23366 17744 23418
rect 17924 23366 17926 23418
rect 17680 23364 17686 23366
rect 17742 23364 17766 23366
rect 17822 23364 17846 23366
rect 17902 23364 17926 23366
rect 17982 23364 17988 23366
rect 17680 23355 17988 23364
rect 18524 23186 18552 24142
rect 18892 24070 18920 25230
rect 19352 24614 19380 25842
rect 19444 25362 19472 26250
rect 19892 25900 19944 25906
rect 19892 25842 19944 25848
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18696 23248 18748 23254
rect 18696 23190 18748 23196
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17500 22568 17552 22574
rect 17500 22510 17552 22516
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17420 21486 17448 21966
rect 17512 21894 17540 22510
rect 17680 22332 17988 22341
rect 17680 22330 17686 22332
rect 17742 22330 17766 22332
rect 17822 22330 17846 22332
rect 17902 22330 17926 22332
rect 17982 22330 17988 22332
rect 17742 22278 17744 22330
rect 17924 22278 17926 22330
rect 17680 22276 17686 22278
rect 17742 22276 17766 22278
rect 17822 22276 17846 22278
rect 17902 22276 17926 22278
rect 17982 22276 17988 22278
rect 17680 22267 17988 22276
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17512 21690 17540 21830
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17680 21244 17988 21253
rect 17680 21242 17686 21244
rect 17742 21242 17766 21244
rect 17822 21242 17846 21244
rect 17902 21242 17926 21244
rect 17982 21242 17988 21244
rect 17742 21190 17744 21242
rect 17924 21190 17926 21242
rect 17680 21188 17686 21190
rect 17742 21188 17766 21190
rect 17822 21188 17846 21190
rect 17902 21188 17926 21190
rect 17982 21188 17988 21190
rect 17680 21179 17988 21188
rect 18156 21146 18184 21490
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 17328 20998 17448 21026
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 17316 20868 17368 20874
rect 17316 20810 17368 20816
rect 17328 20534 17356 20810
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 17316 20528 17368 20534
rect 17316 20470 17368 20476
rect 16960 20058 16988 20470
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17144 19786 17172 19926
rect 17420 19854 17448 20998
rect 18248 20466 18276 23054
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18340 21010 18368 21286
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18432 20466 18460 22918
rect 18708 22574 18736 23190
rect 18892 22642 18920 24006
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 22710 19288 22918
rect 18972 22704 19024 22710
rect 19248 22704 19300 22710
rect 19024 22664 19196 22692
rect 18972 22646 19024 22652
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18696 22568 18748 22574
rect 19168 22556 19196 22664
rect 19248 22646 19300 22652
rect 19248 22568 19300 22574
rect 19168 22528 19248 22556
rect 18696 22510 18748 22516
rect 19248 22510 19300 22516
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18708 21622 18736 21830
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 21010 19104 21286
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 17604 20058 17632 20402
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17680 20156 17988 20165
rect 17680 20154 17686 20156
rect 17742 20154 17766 20156
rect 17822 20154 17846 20156
rect 17902 20154 17926 20156
rect 17982 20154 17988 20156
rect 17742 20102 17744 20154
rect 17924 20102 17926 20154
rect 17680 20100 17686 20102
rect 17742 20100 17766 20102
rect 17822 20100 17846 20102
rect 17902 20100 17926 20102
rect 17982 20100 17988 20102
rect 17680 20091 17988 20100
rect 18064 20058 18092 20334
rect 18616 20330 18644 20878
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18144 20256 18196 20262
rect 18512 20256 18564 20262
rect 18196 20204 18512 20210
rect 18144 20198 18564 20204
rect 18156 20182 18552 20198
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 18696 19780 18748 19786
rect 18696 19722 18748 19728
rect 18708 19514 18736 19722
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 16868 18766 16896 19110
rect 17420 18902 17448 19110
rect 17680 19068 17988 19077
rect 17680 19066 17686 19068
rect 17742 19066 17766 19068
rect 17822 19066 17846 19068
rect 17902 19066 17926 19068
rect 17982 19066 17988 19068
rect 17742 19014 17744 19066
rect 17924 19014 17926 19066
rect 17680 19012 17686 19014
rect 17742 19012 17766 19014
rect 17822 19012 17846 19014
rect 17902 19012 17926 19014
rect 17982 19012 17988 19014
rect 17680 19003 17988 19012
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16408 18358 16436 18634
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15212 15162 15240 17138
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15396 15706 15424 16458
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15672 15502 15700 16390
rect 15764 16182 15792 17070
rect 15948 16250 15976 18226
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15672 15094 15700 15438
rect 16408 15366 16436 18294
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16960 17746 16988 18022
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 17052 17542 17080 18022
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16868 15706 16896 17138
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17328 16250 17356 17070
rect 17420 16998 17448 18838
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18290 17540 18702
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17512 17542 17540 18226
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17604 17796 17632 18158
rect 17680 17980 17988 17989
rect 17680 17978 17686 17980
rect 17742 17978 17766 17980
rect 17822 17978 17846 17980
rect 17902 17978 17926 17980
rect 17982 17978 17988 17980
rect 17742 17926 17744 17978
rect 17924 17926 17926 17978
rect 17680 17924 17686 17926
rect 17742 17924 17766 17926
rect 17822 17924 17846 17926
rect 17902 17924 17926 17926
rect 17982 17924 17988 17926
rect 17680 17915 17988 17924
rect 17684 17808 17736 17814
rect 17604 17768 17684 17796
rect 17684 17750 17736 17756
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16250 17448 16934
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 16408 14958 16436 15302
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 15672 14278 15700 14894
rect 16408 14498 16436 14894
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16316 14470 16436 14498
rect 16316 14414 16344 14470
rect 16868 14414 16896 14758
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15120 14062 15332 14090
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15120 12434 15148 13738
rect 15212 13530 15240 13874
rect 15304 13734 15332 14062
rect 15764 13938 15792 14282
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 15304 13530 15332 13670
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15028 12406 15148 12434
rect 15028 11898 15056 12406
rect 15212 11898 15240 13330
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15304 12306 15332 13194
rect 15856 12918 15884 13670
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14108 10742 14136 10950
rect 14334 10908 14642 10917
rect 14334 10906 14340 10908
rect 14396 10906 14420 10908
rect 14476 10906 14500 10908
rect 14556 10906 14580 10908
rect 14636 10906 14642 10908
rect 14396 10854 14398 10906
rect 14578 10854 14580 10906
rect 14334 10852 14340 10854
rect 14396 10852 14420 10854
rect 14476 10852 14500 10854
rect 14556 10852 14580 10854
rect 14636 10852 14642 10854
rect 14334 10843 14642 10852
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14108 10538 14136 10678
rect 14844 10674 14872 10950
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9178 13308 9862
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13372 6866 13400 7482
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13464 6798 13492 8434
rect 13556 7410 13584 9318
rect 13740 8090 13768 9522
rect 13832 8838 13860 9590
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13832 7954 13860 8774
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6390 12664 6598
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 13464 6322 13492 6734
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13464 5846 13492 6258
rect 13740 5846 13768 6734
rect 13924 6458 13952 7822
rect 14108 7546 14136 10474
rect 14844 10130 14872 10610
rect 15304 10606 15332 11630
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14200 8090 14228 9930
rect 14334 9820 14642 9829
rect 14334 9818 14340 9820
rect 14396 9818 14420 9820
rect 14476 9818 14500 9820
rect 14556 9818 14580 9820
rect 14636 9818 14642 9820
rect 14396 9766 14398 9818
rect 14578 9766 14580 9818
rect 14334 9764 14340 9766
rect 14396 9764 14420 9766
rect 14476 9764 14500 9766
rect 14556 9764 14580 9766
rect 14636 9764 14642 9766
rect 14334 9755 14642 9764
rect 14844 9518 14872 9930
rect 15212 9602 15240 10474
rect 15304 10130 15332 10542
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15396 10062 15424 11698
rect 15948 11082 15976 12174
rect 16040 11762 16068 13126
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16132 11898 16160 12106
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16684 11762 16712 12582
rect 16776 12442 16804 13262
rect 16960 12986 16988 13670
rect 17144 12986 17172 15098
rect 17236 14822 17264 15982
rect 17328 15162 17356 16186
rect 17420 15978 17448 16186
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17512 15502 17540 17478
rect 17604 16658 17632 17546
rect 17696 17202 17724 17750
rect 18248 17746 18276 19246
rect 18432 18970 18460 19314
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18708 18766 18736 19110
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 18290 18460 18566
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18156 17270 18184 17478
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 18800 17134 18828 20402
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19076 19378 19104 20198
rect 19260 19922 19288 20334
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 17680 16892 17988 16901
rect 17680 16890 17686 16892
rect 17742 16890 17766 16892
rect 17822 16890 17846 16892
rect 17902 16890 17926 16892
rect 17982 16890 17988 16892
rect 17742 16838 17744 16890
rect 17924 16838 17926 16890
rect 17680 16836 17686 16838
rect 17742 16836 17766 16838
rect 17822 16836 17846 16838
rect 17902 16836 17926 16838
rect 17982 16836 17988 16838
rect 17680 16827 17988 16836
rect 18800 16794 18828 17070
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18708 16250 18736 16526
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 17680 15804 17988 15813
rect 17680 15802 17686 15804
rect 17742 15802 17766 15804
rect 17822 15802 17846 15804
rect 17902 15802 17926 15804
rect 17982 15802 17988 15804
rect 17742 15750 17744 15802
rect 17924 15750 17926 15802
rect 17680 15748 17686 15750
rect 17742 15748 17766 15750
rect 17822 15748 17846 15750
rect 17902 15748 17926 15750
rect 17982 15748 17988 15750
rect 17680 15739 17988 15748
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17604 15094 17632 15506
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 13530 17264 14758
rect 17604 14618 17632 15030
rect 17680 14716 17988 14725
rect 17680 14714 17686 14716
rect 17742 14714 17766 14716
rect 17822 14714 17846 14716
rect 17902 14714 17926 14716
rect 17982 14714 17988 14716
rect 17742 14662 17744 14714
rect 17924 14662 17926 14714
rect 17680 14660 17686 14662
rect 17742 14660 17766 14662
rect 17822 14660 17846 14662
rect 17902 14660 17926 14662
rect 17982 14660 17988 14662
rect 17680 14651 17988 14660
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17328 13394 17356 13806
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17328 12986 17356 13330
rect 17420 13326 17448 13738
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17498 13288 17554 13297
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 17144 12170 17172 12922
rect 17420 12918 17448 13262
rect 17498 13223 17500 13232
rect 17552 13223 17554 13232
rect 17500 13194 17552 13200
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 12442 17356 12582
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15028 9586 15240 9602
rect 15016 9580 15240 9586
rect 15068 9574 15240 9580
rect 15016 9522 15068 9528
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8974 14596 9318
rect 15212 9042 15240 9574
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14334 8732 14642 8741
rect 14334 8730 14340 8732
rect 14396 8730 14420 8732
rect 14476 8730 14500 8732
rect 14556 8730 14580 8732
rect 14636 8730 14642 8732
rect 14396 8678 14398 8730
rect 14578 8678 14580 8730
rect 14334 8676 14340 8678
rect 14396 8676 14420 8678
rect 14476 8676 14500 8678
rect 14556 8676 14580 8678
rect 14636 8676 14642 8678
rect 14334 8667 14642 8676
rect 15396 8498 15424 9998
rect 15488 9654 15516 10610
rect 15948 10538 15976 11018
rect 16684 10810 16712 11086
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16776 10062 16804 10474
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15856 9722 15884 9862
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 8634 15976 9522
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16132 8498 16160 9862
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16316 9042 16344 9658
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16592 8634 16620 9930
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16868 8566 16896 11698
rect 17144 11354 17172 12106
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17328 11082 17356 11698
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17328 10674 17356 11018
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 10010 17356 10066
rect 17420 10010 17448 12718
rect 17604 12434 17632 13874
rect 17680 13628 17988 13637
rect 17680 13626 17686 13628
rect 17742 13626 17766 13628
rect 17822 13626 17846 13628
rect 17902 13626 17926 13628
rect 17982 13626 17988 13628
rect 17742 13574 17744 13626
rect 17924 13574 17926 13626
rect 17680 13572 17686 13574
rect 17742 13572 17766 13574
rect 17822 13572 17846 13574
rect 17902 13572 17926 13574
rect 17982 13572 17988 13574
rect 17680 13563 17988 13572
rect 18340 13530 18368 14418
rect 18984 14006 19012 14486
rect 19076 14278 19104 19314
rect 19260 19242 19288 19858
rect 19352 19854 19380 24550
rect 19720 24138 19748 24754
rect 19904 24206 19932 25842
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20088 24274 20116 25774
rect 20180 25498 20208 26318
rect 21026 26140 21334 26149
rect 21026 26138 21032 26140
rect 21088 26138 21112 26140
rect 21168 26138 21192 26140
rect 21248 26138 21272 26140
rect 21328 26138 21334 26140
rect 21088 26086 21090 26138
rect 21270 26086 21272 26138
rect 21026 26084 21032 26086
rect 21088 26084 21112 26086
rect 21168 26084 21192 26086
rect 21248 26084 21272 26086
rect 21328 26084 21334 26086
rect 21026 26075 21334 26084
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 20720 25356 20772 25362
rect 20720 25298 20772 25304
rect 20732 24954 20760 25298
rect 20824 25294 20852 25774
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20916 24818 20944 25298
rect 21026 25052 21334 25061
rect 21026 25050 21032 25052
rect 21088 25050 21112 25052
rect 21168 25050 21192 25052
rect 21248 25050 21272 25052
rect 21328 25050 21334 25052
rect 21088 24998 21090 25050
rect 21270 24998 21272 25050
rect 21026 24996 21032 24998
rect 21088 24996 21112 24998
rect 21168 24996 21192 24998
rect 21248 24996 21272 24998
rect 21328 24996 21334 24998
rect 21026 24987 21334 24996
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19904 23866 19932 24142
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 20088 23576 20116 24210
rect 20916 24206 20944 24754
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 19812 23548 20116 23576
rect 19812 22642 19840 23548
rect 20180 23186 20208 23802
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20180 22642 20208 23122
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 19432 22500 19484 22506
rect 19432 22442 19484 22448
rect 19444 22234 19472 22442
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 19524 21888 19576 21894
rect 19524 21830 19576 21836
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19536 19718 19564 21830
rect 20364 21690 20392 22034
rect 20456 22030 20484 22918
rect 20732 22710 20760 22986
rect 20916 22778 20944 24142
rect 21456 24132 21508 24138
rect 21456 24074 21508 24080
rect 21026 23964 21334 23973
rect 21026 23962 21032 23964
rect 21088 23962 21112 23964
rect 21168 23962 21192 23964
rect 21248 23962 21272 23964
rect 21328 23962 21334 23964
rect 21088 23910 21090 23962
rect 21270 23910 21272 23962
rect 21026 23908 21032 23910
rect 21088 23908 21112 23910
rect 21168 23908 21192 23910
rect 21248 23908 21272 23910
rect 21328 23908 21334 23910
rect 21026 23899 21334 23908
rect 21468 23186 21496 24074
rect 21456 23180 21508 23186
rect 21456 23122 21508 23128
rect 21026 22876 21334 22885
rect 21026 22874 21032 22876
rect 21088 22874 21112 22876
rect 21168 22874 21192 22876
rect 21248 22874 21272 22876
rect 21328 22874 21334 22876
rect 21088 22822 21090 22874
rect 21270 22822 21272 22874
rect 21026 22820 21032 22822
rect 21088 22820 21112 22822
rect 21168 22820 21192 22822
rect 21248 22820 21272 22822
rect 21328 22820 21334 22822
rect 21026 22811 21334 22820
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20720 22704 20772 22710
rect 20720 22646 20772 22652
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 19812 20058 19840 21490
rect 20364 20602 20392 21626
rect 20824 21146 20852 22170
rect 22020 22030 22048 22374
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19352 19446 19380 19654
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19616 19236 19668 19242
rect 19616 19178 19668 19184
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19352 17270 19380 18294
rect 19628 17882 19656 19178
rect 20180 18970 20208 20402
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20548 19378 20576 19654
rect 20640 19514 20668 20402
rect 20824 19854 20852 21082
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20916 19786 20944 21966
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21026 21788 21334 21797
rect 21026 21786 21032 21788
rect 21088 21786 21112 21788
rect 21168 21786 21192 21788
rect 21248 21786 21272 21788
rect 21328 21786 21334 21788
rect 21088 21734 21090 21786
rect 21270 21734 21272 21786
rect 21026 21732 21032 21734
rect 21088 21732 21112 21734
rect 21168 21732 21192 21734
rect 21248 21732 21272 21734
rect 21328 21732 21334 21734
rect 21026 21723 21334 21732
rect 21376 21554 21404 21830
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21284 21146 21312 21490
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21026 20700 21334 20709
rect 21026 20698 21032 20700
rect 21088 20698 21112 20700
rect 21168 20698 21192 20700
rect 21248 20698 21272 20700
rect 21328 20698 21334 20700
rect 21088 20646 21090 20698
rect 21270 20646 21272 20698
rect 21026 20644 21032 20646
rect 21088 20644 21112 20646
rect 21168 20644 21192 20646
rect 21248 20644 21272 20646
rect 21328 20644 21334 20646
rect 21026 20635 21334 20644
rect 21376 20262 21404 21286
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21560 20602 21588 20878
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21744 20330 21772 21966
rect 22020 21690 22048 21966
rect 23492 21894 23520 26318
rect 24372 25596 24680 25605
rect 24372 25594 24378 25596
rect 24434 25594 24458 25596
rect 24514 25594 24538 25596
rect 24594 25594 24618 25596
rect 24674 25594 24680 25596
rect 24434 25542 24436 25594
rect 24616 25542 24618 25594
rect 24372 25540 24378 25542
rect 24434 25540 24458 25542
rect 24514 25540 24538 25542
rect 24594 25540 24618 25542
rect 24674 25540 24680 25542
rect 24372 25531 24680 25540
rect 24372 24508 24680 24517
rect 24372 24506 24378 24508
rect 24434 24506 24458 24508
rect 24514 24506 24538 24508
rect 24594 24506 24618 24508
rect 24674 24506 24680 24508
rect 24434 24454 24436 24506
rect 24616 24454 24618 24506
rect 24372 24452 24378 24454
rect 24434 24452 24458 24454
rect 24514 24452 24538 24454
rect 24594 24452 24618 24454
rect 24674 24452 24680 24454
rect 24372 24443 24680 24452
rect 24372 23420 24680 23429
rect 24372 23418 24378 23420
rect 24434 23418 24458 23420
rect 24514 23418 24538 23420
rect 24594 23418 24618 23420
rect 24674 23418 24680 23420
rect 24434 23366 24436 23418
rect 24616 23366 24618 23418
rect 24372 23364 24378 23366
rect 24434 23364 24458 23366
rect 24514 23364 24538 23366
rect 24594 23364 24618 23366
rect 24674 23364 24680 23366
rect 24372 23355 24680 23364
rect 24372 22332 24680 22341
rect 24372 22330 24378 22332
rect 24434 22330 24458 22332
rect 24514 22330 24538 22332
rect 24594 22330 24618 22332
rect 24674 22330 24680 22332
rect 24434 22278 24436 22330
rect 24616 22278 24618 22330
rect 24372 22276 24378 22278
rect 24434 22276 24458 22278
rect 24514 22276 24538 22278
rect 24594 22276 24618 22278
rect 24674 22276 24680 22278
rect 24372 22267 24680 22276
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 26344 21690 26372 26318
rect 27718 26140 28026 26149
rect 27718 26138 27724 26140
rect 27780 26138 27804 26140
rect 27860 26138 27884 26140
rect 27940 26138 27964 26140
rect 28020 26138 28026 26140
rect 27780 26086 27782 26138
rect 27962 26086 27964 26138
rect 27718 26084 27724 26086
rect 27780 26084 27804 26086
rect 27860 26084 27884 26086
rect 27940 26084 27964 26086
rect 28020 26084 28026 26086
rect 27718 26075 28026 26084
rect 27718 25052 28026 25061
rect 27718 25050 27724 25052
rect 27780 25050 27804 25052
rect 27860 25050 27884 25052
rect 27940 25050 27964 25052
rect 28020 25050 28026 25052
rect 27780 24998 27782 25050
rect 27962 24998 27964 25050
rect 27718 24996 27724 24998
rect 27780 24996 27804 24998
rect 27860 24996 27884 24998
rect 27940 24996 27964 24998
rect 28020 24996 28026 24998
rect 27718 24987 28026 24996
rect 27718 23964 28026 23973
rect 27718 23962 27724 23964
rect 27780 23962 27804 23964
rect 27860 23962 27884 23964
rect 27940 23962 27964 23964
rect 28020 23962 28026 23964
rect 27780 23910 27782 23962
rect 27962 23910 27964 23962
rect 27718 23908 27724 23910
rect 27780 23908 27804 23910
rect 27860 23908 27884 23910
rect 27940 23908 27964 23910
rect 28020 23908 28026 23910
rect 27718 23899 28026 23908
rect 27718 22876 28026 22885
rect 27718 22874 27724 22876
rect 27780 22874 27804 22876
rect 27860 22874 27884 22876
rect 27940 22874 27964 22876
rect 28020 22874 28026 22876
rect 27780 22822 27782 22874
rect 27962 22822 27964 22874
rect 27718 22820 27724 22822
rect 27780 22820 27804 22822
rect 27860 22820 27884 22822
rect 27940 22820 27964 22822
rect 28020 22820 28026 22822
rect 27718 22811 28026 22820
rect 27718 21788 28026 21797
rect 27718 21786 27724 21788
rect 27780 21786 27804 21788
rect 27860 21786 27884 21788
rect 27940 21786 27964 21788
rect 28020 21786 28026 21788
rect 27780 21734 27782 21786
rect 27962 21734 27964 21786
rect 27718 21732 27724 21734
rect 27780 21732 27804 21734
rect 27860 21732 27884 21734
rect 27940 21732 27964 21734
rect 28020 21732 28026 21734
rect 27718 21723 28026 21732
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 26332 21684 26384 21690
rect 26332 21626 26384 21632
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21928 20942 21956 21422
rect 24372 21244 24680 21253
rect 24372 21242 24378 21244
rect 24434 21242 24458 21244
rect 24514 21242 24538 21244
rect 24594 21242 24618 21244
rect 24674 21242 24680 21244
rect 24434 21190 24436 21242
rect 24616 21190 24618 21242
rect 24372 21188 24378 21190
rect 24434 21188 24458 21190
rect 24514 21188 24538 21190
rect 24594 21188 24618 21190
rect 24674 21188 24680 21190
rect 24372 21179 24680 21188
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21928 19854 21956 20878
rect 23480 20868 23532 20874
rect 23480 20810 23532 20816
rect 23492 20602 23520 20810
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20602 23704 20742
rect 27718 20700 28026 20709
rect 27718 20698 27724 20700
rect 27780 20698 27804 20700
rect 27860 20698 27884 20700
rect 27940 20698 27964 20700
rect 28020 20698 28026 20700
rect 27780 20646 27782 20698
rect 27962 20646 27964 20698
rect 27718 20644 27724 20646
rect 27780 20644 27804 20646
rect 27860 20644 27884 20646
rect 27940 20644 27964 20646
rect 28020 20644 28026 20646
rect 27718 20635 28026 20644
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19708 17536 19760 17542
rect 19984 17536 20036 17542
rect 19760 17496 19840 17524
rect 19708 17478 19760 17484
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16590 19196 17070
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19628 16590 19656 16730
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19524 16176 19576 16182
rect 19524 16118 19576 16124
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15094 19472 15302
rect 19536 15094 19564 16118
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15502 19656 15846
rect 19720 15706 19748 16458
rect 19708 15700 19760 15706
rect 19708 15642 19760 15648
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19352 14414 19380 14962
rect 19536 14414 19564 15030
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 19352 14074 19380 14350
rect 19812 14346 19840 17496
rect 19984 17478 20036 17484
rect 19996 17270 20024 17478
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20180 15162 20208 17138
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12918 18552 13126
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 17680 12540 17988 12549
rect 17680 12538 17686 12540
rect 17742 12538 17766 12540
rect 17822 12538 17846 12540
rect 17902 12538 17926 12540
rect 17982 12538 17988 12540
rect 17742 12486 17744 12538
rect 17924 12486 17926 12538
rect 17680 12484 17686 12486
rect 17742 12484 17766 12486
rect 17822 12484 17846 12486
rect 17902 12484 17926 12486
rect 17982 12484 17988 12486
rect 17680 12475 17988 12484
rect 17604 12406 17724 12434
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17500 11688 17552 11694
rect 17500 11630 17552 11636
rect 17512 10606 17540 11630
rect 17604 11354 17632 11766
rect 17696 11762 17724 12406
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17680 11452 17988 11461
rect 17680 11450 17686 11452
rect 17742 11450 17766 11452
rect 17822 11450 17846 11452
rect 17902 11450 17926 11452
rect 17982 11450 17988 11452
rect 17742 11398 17744 11450
rect 17924 11398 17926 11450
rect 17680 11396 17686 11398
rect 17742 11396 17766 11398
rect 17822 11396 17846 11398
rect 17902 11396 17926 11398
rect 17982 11396 17988 11398
rect 17680 11387 17988 11396
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 18064 11150 18092 12038
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17512 10062 17540 10542
rect 17680 10364 17988 10373
rect 17680 10362 17686 10364
rect 17742 10362 17766 10364
rect 17822 10362 17846 10364
rect 17902 10362 17926 10364
rect 17982 10362 17988 10364
rect 17742 10310 17744 10362
rect 17924 10310 17926 10362
rect 17680 10308 17686 10310
rect 17742 10308 17766 10310
rect 17822 10308 17846 10310
rect 17902 10308 17926 10310
rect 17982 10308 17988 10310
rect 17680 10299 17988 10308
rect 17328 9982 17448 10010
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17420 9518 17448 9982
rect 17512 9654 17540 9998
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17592 9580 17644 9586
rect 17592 9522 17644 9528
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17328 9178 17356 9454
rect 17604 9178 17632 9522
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17680 9276 17988 9285
rect 17680 9274 17686 9276
rect 17742 9274 17766 9276
rect 17822 9274 17846 9276
rect 17902 9274 17926 9276
rect 17982 9274 17988 9276
rect 17742 9222 17744 9274
rect 17924 9222 17926 9274
rect 17680 9220 17686 9222
rect 17742 9220 17766 9222
rect 17822 9220 17846 9222
rect 17902 9220 17926 9222
rect 17982 9220 17988 9222
rect 17680 9211 17988 9220
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14334 7644 14642 7653
rect 14334 7642 14340 7644
rect 14396 7642 14420 7644
rect 14476 7642 14500 7644
rect 14556 7642 14580 7644
rect 14636 7642 14642 7644
rect 14396 7590 14398 7642
rect 14578 7590 14580 7642
rect 14334 7588 14340 7590
rect 14396 7588 14420 7590
rect 14476 7588 14500 7590
rect 14556 7588 14580 7590
rect 14636 7588 14642 7590
rect 14334 7579 14642 7588
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14844 7478 14872 7686
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 15028 7206 15056 7822
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14334 6556 14642 6565
rect 14334 6554 14340 6556
rect 14396 6554 14420 6556
rect 14476 6554 14500 6556
rect 14556 6554 14580 6556
rect 14636 6554 14642 6556
rect 14396 6502 14398 6554
rect 14578 6502 14580 6554
rect 14334 6500 14340 6502
rect 14396 6500 14420 6502
rect 14476 6500 14500 6502
rect 14556 6500 14580 6502
rect 14636 6500 14642 6502
rect 14334 6491 14642 6500
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5914 14044 6054
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 15028 5710 15056 7142
rect 15212 7002 15240 7754
rect 15304 7342 15332 8230
rect 16960 7886 16988 9114
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15948 6458 15976 7346
rect 16500 7002 16528 7686
rect 16960 7410 16988 7822
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 17236 6798 17264 8910
rect 17680 8188 17988 8197
rect 17680 8186 17686 8188
rect 17742 8186 17766 8188
rect 17822 8186 17846 8188
rect 17902 8186 17926 8188
rect 17982 8186 17988 8188
rect 17742 8134 17744 8186
rect 17924 8134 17926 8186
rect 17680 8132 17686 8134
rect 17742 8132 17766 8134
rect 17822 8132 17846 8134
rect 17902 8132 17926 8134
rect 17982 8132 17988 8134
rect 17680 8123 17988 8132
rect 18064 7970 18092 9386
rect 18156 9178 18184 12854
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18524 10606 18552 12242
rect 18708 11354 18736 12786
rect 18892 12646 18920 13262
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12850 19380 13126
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18892 12238 18920 12582
rect 18984 12306 19012 12582
rect 19076 12442 19104 12650
rect 19064 12436 19116 12442
rect 19444 12434 19472 13262
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19064 12378 19116 12384
rect 19352 12406 19472 12434
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 19352 12170 19380 12406
rect 19536 12238 19564 13194
rect 19628 12986 19656 13874
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11898 19012 12038
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18800 11150 18828 11698
rect 18984 11218 19012 11834
rect 19352 11354 19380 12106
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 19536 10792 19564 12174
rect 19720 11898 19748 12854
rect 19812 12850 19840 14282
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 19996 12986 20024 13330
rect 20088 13190 20116 13330
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 20180 11898 20208 14894
rect 20364 14618 20392 17138
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20456 12889 20484 19314
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20640 17678 20668 18362
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20548 17202 20576 17478
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20732 16590 20760 19654
rect 21026 19612 21334 19621
rect 21026 19610 21032 19612
rect 21088 19610 21112 19612
rect 21168 19610 21192 19612
rect 21248 19610 21272 19612
rect 21328 19610 21334 19612
rect 21088 19558 21090 19610
rect 21270 19558 21272 19610
rect 21026 19556 21032 19558
rect 21088 19556 21112 19558
rect 21168 19556 21192 19558
rect 21248 19556 21272 19558
rect 21328 19556 21334 19558
rect 21026 19547 21334 19556
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20824 18970 20852 19382
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20824 17746 20852 18906
rect 20916 18426 20944 19314
rect 21026 18524 21334 18533
rect 21026 18522 21032 18524
rect 21088 18522 21112 18524
rect 21168 18522 21192 18524
rect 21248 18522 21272 18524
rect 21328 18522 21334 18524
rect 21088 18470 21090 18522
rect 21270 18470 21272 18522
rect 21026 18468 21032 18470
rect 21088 18468 21112 18470
rect 21168 18468 21192 18470
rect 21248 18468 21272 18470
rect 21328 18468 21334 18470
rect 21026 18459 21334 18468
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20916 18290 20944 18362
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20442 12880 20498 12889
rect 20442 12815 20444 12824
rect 20496 12815 20498 12824
rect 20444 12786 20496 12792
rect 20456 12755 20484 12786
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11898 20484 12038
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 19708 11620 19760 11626
rect 19708 11562 19760 11568
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19352 10764 19564 10792
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 9518 18368 10202
rect 18432 9926 18460 10542
rect 18524 10130 18552 10542
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18432 9330 18460 9862
rect 18340 9302 18460 9330
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18340 8430 18368 9302
rect 18524 9194 18552 10066
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19260 9586 19288 9930
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18432 9166 18552 9194
rect 18432 8430 18460 9166
rect 18892 8974 18920 9318
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 17972 7942 18092 7970
rect 17972 7750 18000 7942
rect 18248 7886 18276 8230
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18144 7812 18196 7818
rect 18144 7754 18196 7760
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7342 18000 7686
rect 18156 7546 18184 7754
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18340 7478 18368 8366
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 7546 18460 7822
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18524 7392 18552 8434
rect 18616 8090 18644 8910
rect 18708 8362 18736 8910
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18604 7404 18656 7410
rect 18524 7364 18604 7392
rect 18604 7346 18656 7352
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17680 7100 17988 7109
rect 17680 7098 17686 7100
rect 17742 7098 17766 7100
rect 17822 7098 17846 7100
rect 17902 7098 17926 7100
rect 17982 7098 17988 7100
rect 17742 7046 17744 7098
rect 17924 7046 17926 7098
rect 17680 7044 17686 7046
rect 17742 7044 17766 7046
rect 17822 7044 17846 7046
rect 17902 7044 17926 7046
rect 17982 7044 17988 7046
rect 17680 7035 17988 7044
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 17224 6792 17276 6798
rect 17144 6752 17224 6780
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5710 15148 6190
rect 15580 5710 15608 6258
rect 16132 5778 16160 6666
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6458 16528 6598
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16500 5710 16528 6394
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 14334 5468 14642 5477
rect 14334 5466 14340 5468
rect 14396 5466 14420 5468
rect 14476 5466 14500 5468
rect 14556 5466 14580 5468
rect 14636 5466 14642 5468
rect 14396 5414 14398 5466
rect 14578 5414 14580 5466
rect 14334 5412 14340 5414
rect 14396 5412 14420 5414
rect 14476 5412 14500 5414
rect 14556 5412 14580 5414
rect 14636 5412 14642 5414
rect 14334 5403 14642 5412
rect 15120 5370 15148 5646
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 16868 5302 16896 6190
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 17144 5234 17172 6752
rect 17224 6734 17276 6740
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6390 17264 6598
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17604 5778 17632 6326
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 17680 6012 17988 6021
rect 17680 6010 17686 6012
rect 17742 6010 17766 6012
rect 17822 6010 17846 6012
rect 17902 6010 17926 6012
rect 17982 6010 17988 6012
rect 17742 5958 17744 6010
rect 17924 5958 17926 6010
rect 17680 5956 17686 5958
rect 17742 5956 17766 5958
rect 17822 5956 17846 5958
rect 17902 5956 17926 5958
rect 17982 5956 17988 5958
rect 17680 5947 17988 5956
rect 18432 5914 18460 6190
rect 18524 6118 18552 6802
rect 18616 6798 18644 7346
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 18524 5710 18552 6054
rect 18800 5778 18828 6598
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18892 5642 18920 7346
rect 18984 7342 19012 8434
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19352 6866 19380 10764
rect 19628 10742 19656 11018
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19444 9586 19472 10406
rect 19536 10266 19564 10610
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19444 8430 19472 8774
rect 19536 8566 19564 9998
rect 19720 8566 19748 11562
rect 20180 11150 20208 11834
rect 20456 11626 20484 11834
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20456 11082 20484 11562
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19812 10062 19840 10950
rect 20548 10810 20576 16526
rect 20824 16250 20852 17546
rect 20916 16726 20944 18022
rect 21026 17436 21334 17445
rect 21026 17434 21032 17436
rect 21088 17434 21112 17436
rect 21168 17434 21192 17436
rect 21248 17434 21272 17436
rect 21328 17434 21334 17436
rect 21088 17382 21090 17434
rect 21270 17382 21272 17434
rect 21026 17380 21032 17382
rect 21088 17380 21112 17382
rect 21168 17380 21192 17382
rect 21248 17380 21272 17382
rect 21328 17380 21334 17382
rect 21026 17371 21334 17380
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 21100 16590 21128 17002
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21026 16348 21334 16357
rect 21026 16346 21032 16348
rect 21088 16346 21112 16348
rect 21168 16346 21192 16348
rect 21248 16346 21272 16348
rect 21328 16346 21334 16348
rect 21088 16294 21090 16346
rect 21270 16294 21272 16346
rect 21026 16292 21032 16294
rect 21088 16292 21112 16294
rect 21168 16292 21192 16294
rect 21248 16292 21272 16294
rect 21328 16292 21334 16294
rect 21026 16283 21334 16292
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20824 15706 20852 15982
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20916 14958 20944 15914
rect 21376 15502 21404 16934
rect 21468 15502 21496 19790
rect 21640 19440 21692 19446
rect 21640 19382 21692 19388
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21560 18834 21588 19110
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21652 16114 21680 19382
rect 22112 19310 22140 20334
rect 23676 19922 23704 20538
rect 24372 20156 24680 20165
rect 24372 20154 24378 20156
rect 24434 20154 24458 20156
rect 24514 20154 24538 20156
rect 24594 20154 24618 20156
rect 24674 20154 24680 20156
rect 24434 20102 24436 20154
rect 24616 20102 24618 20154
rect 24372 20100 24378 20102
rect 24434 20100 24458 20102
rect 24514 20100 24538 20102
rect 24594 20100 24618 20102
rect 24674 20100 24680 20102
rect 24372 20091 24680 20100
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 23664 19916 23716 19922
rect 23664 19858 23716 19864
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22296 19514 22324 19654
rect 23584 19514 23612 19790
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21836 17882 21864 19246
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21928 17066 21956 18226
rect 22112 17678 22140 18566
rect 22296 17814 22324 19450
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23492 18766 23520 19314
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22848 18358 22876 18634
rect 23584 18426 23612 19314
rect 24372 19068 24680 19077
rect 24372 19066 24378 19068
rect 24434 19066 24458 19068
rect 24514 19066 24538 19068
rect 24594 19066 24618 19068
rect 24674 19066 24680 19068
rect 24434 19014 24436 19066
rect 24616 19014 24618 19066
rect 24372 19012 24378 19014
rect 24434 19012 24458 19014
rect 24514 19012 24538 19014
rect 24594 19012 24618 19014
rect 24674 19012 24680 19014
rect 24372 19003 24680 19012
rect 24676 18760 24728 18766
rect 24728 18720 24808 18748
rect 24676 18702 24728 18708
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21928 16794 21956 17002
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 22020 16114 22048 17478
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 22020 15450 22048 15914
rect 22112 15638 22140 17070
rect 22204 16522 22232 17206
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22296 16250 22324 17614
rect 22388 17202 22416 18226
rect 24372 17980 24680 17989
rect 24372 17978 24378 17980
rect 24434 17978 24458 17980
rect 24514 17978 24538 17980
rect 24594 17978 24618 17980
rect 24674 17978 24680 17980
rect 24434 17926 24436 17978
rect 24616 17926 24618 17978
rect 24372 17924 24378 17926
rect 24434 17924 24458 17926
rect 24514 17924 24538 17926
rect 24594 17924 24618 17926
rect 24674 17924 24680 17926
rect 24372 17915 24680 17924
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22480 16794 22508 17682
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22388 16182 22416 16390
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 21026 15260 21334 15269
rect 21026 15258 21032 15260
rect 21088 15258 21112 15260
rect 21168 15258 21192 15260
rect 21248 15258 21272 15260
rect 21328 15258 21334 15260
rect 21088 15206 21090 15258
rect 21270 15206 21272 15258
rect 21026 15204 21032 15206
rect 21088 15204 21112 15206
rect 21168 15204 21192 15206
rect 21248 15204 21272 15206
rect 21328 15204 21334 15206
rect 21026 15195 21334 15204
rect 21468 15026 21496 15438
rect 22020 15422 22140 15450
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 14074 20944 14350
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21026 14172 21334 14181
rect 21026 14170 21032 14172
rect 21088 14170 21112 14172
rect 21168 14170 21192 14172
rect 21248 14170 21272 14172
rect 21328 14170 21334 14172
rect 21088 14118 21090 14170
rect 21270 14118 21272 14170
rect 21026 14116 21032 14118
rect 21088 14116 21112 14118
rect 21168 14116 21192 14118
rect 21248 14116 21272 14118
rect 21328 14116 21334 14118
rect 21026 14107 21334 14116
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20916 13870 20944 14010
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20732 13394 20760 13670
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 21026 13084 21334 13093
rect 21026 13082 21032 13084
rect 21088 13082 21112 13084
rect 21168 13082 21192 13084
rect 21248 13082 21272 13084
rect 21328 13082 21334 13084
rect 21088 13030 21090 13082
rect 21270 13030 21272 13082
rect 21026 13028 21032 13030
rect 21088 13028 21112 13030
rect 21168 13028 21192 13030
rect 21248 13028 21272 13030
rect 21328 13028 21334 13030
rect 21026 13019 21334 13028
rect 21376 12986 21404 14282
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21468 12850 21496 14758
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21928 12986 21956 13874
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22020 13394 22048 13806
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20640 11354 20668 11494
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 11218 20760 12582
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21026 11996 21334 12005
rect 21026 11994 21032 11996
rect 21088 11994 21112 11996
rect 21168 11994 21192 11996
rect 21248 11994 21272 11996
rect 21328 11994 21334 11996
rect 21088 11942 21090 11994
rect 21270 11942 21272 11994
rect 21026 11940 21032 11942
rect 21088 11940 21112 11942
rect 21168 11940 21192 11942
rect 21248 11940 21272 11942
rect 21328 11940 21334 11942
rect 21026 11931 21334 11940
rect 21744 11354 21772 12174
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11830 21956 12038
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21026 10908 21334 10917
rect 21026 10906 21032 10908
rect 21088 10906 21112 10908
rect 21168 10906 21192 10908
rect 21248 10906 21272 10908
rect 21328 10906 21334 10908
rect 21088 10854 21090 10906
rect 21270 10854 21272 10906
rect 21026 10852 21032 10854
rect 21088 10852 21112 10854
rect 21168 10852 21192 10854
rect 21248 10852 21272 10854
rect 21328 10852 21334 10854
rect 21026 10843 21334 10852
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 21376 10674 21404 10950
rect 22020 10674 22048 13330
rect 22112 12850 22140 15422
rect 22940 15366 22968 17478
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23308 16182 23336 17070
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22480 14618 22508 15030
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22664 14634 22692 14962
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 22664 14618 22784 14634
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22652 14612 22784 14618
rect 22704 14606 22784 14612
rect 22652 14554 22704 14560
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22664 13190 22692 14418
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22664 12782 22692 13126
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22480 12442 22508 12718
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22756 11898 22784 14606
rect 23216 14278 23244 14894
rect 23308 14414 23336 15846
rect 23400 15706 23428 16458
rect 23492 16266 23520 16594
rect 23584 16522 23612 17614
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23492 16238 23704 16266
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23216 13530 23244 14214
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23308 12918 23336 14350
rect 23400 13734 23428 15506
rect 23492 15502 23520 15914
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23492 13938 23520 14962
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 12986 23428 13670
rect 23676 13462 23704 16238
rect 23768 15026 23796 17614
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 23952 17202 23980 17478
rect 24228 17270 24256 17478
rect 24596 17338 24624 17614
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 24372 16892 24680 16901
rect 24372 16890 24378 16892
rect 24434 16890 24458 16892
rect 24514 16890 24538 16892
rect 24594 16890 24618 16892
rect 24674 16890 24680 16892
rect 24434 16838 24436 16890
rect 24616 16838 24618 16890
rect 24372 16836 24378 16838
rect 24434 16836 24458 16838
rect 24514 16836 24538 16838
rect 24594 16836 24618 16838
rect 24674 16836 24680 16838
rect 24372 16827 24680 16836
rect 24676 16652 24728 16658
rect 24780 16640 24808 18720
rect 24728 16612 24808 16640
rect 24676 16594 24728 16600
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23952 15978 23980 16458
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 24372 15804 24680 15813
rect 24372 15802 24378 15804
rect 24434 15802 24458 15804
rect 24514 15802 24538 15804
rect 24594 15802 24618 15804
rect 24674 15802 24680 15804
rect 24434 15750 24436 15802
rect 24616 15750 24618 15802
rect 24372 15748 24378 15750
rect 24434 15748 24458 15750
rect 24514 15748 24538 15750
rect 24594 15748 24618 15750
rect 24674 15748 24680 15750
rect 24372 15739 24680 15748
rect 24872 15706 24900 19994
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19310 25452 19654
rect 25884 19514 25912 19790
rect 27718 19612 28026 19621
rect 27718 19610 27724 19612
rect 27780 19610 27804 19612
rect 27860 19610 27884 19612
rect 27940 19610 27964 19612
rect 28020 19610 28026 19612
rect 27780 19558 27782 19610
rect 27962 19558 27964 19610
rect 27718 19556 27724 19558
rect 27780 19556 27804 19558
rect 27860 19556 27884 19558
rect 27940 19556 27964 19558
rect 28020 19556 28026 19558
rect 27718 19547 28026 19556
rect 25872 19508 25924 19514
rect 25872 19450 25924 19456
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25516 18834 25544 19314
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25320 18760 25372 18766
rect 25320 18702 25372 18708
rect 25332 18290 25360 18702
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25332 16590 25360 18226
rect 25412 17128 25464 17134
rect 25412 17070 25464 17076
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25424 16538 25452 17070
rect 25596 16584 25648 16590
rect 25424 16522 25544 16538
rect 25596 16526 25648 16532
rect 25424 16516 25556 16522
rect 25424 16510 25504 16516
rect 25504 16458 25556 16464
rect 25608 15910 25636 16526
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 24872 14958 24900 15438
rect 25044 15428 25096 15434
rect 25044 15370 25096 15376
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 25056 14890 25084 15370
rect 25608 15026 25636 15846
rect 25792 15570 25820 18634
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26252 16658 26280 18090
rect 26344 17542 26372 19314
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26528 17610 26556 18158
rect 26516 17604 26568 17610
rect 26516 17546 26568 17552
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26344 15706 26372 16934
rect 26332 15700 26384 15706
rect 26332 15642 26384 15648
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 26436 15162 26464 17138
rect 26620 15366 26648 18702
rect 27080 17746 27108 19110
rect 27344 18692 27396 18698
rect 27344 18634 27396 18640
rect 27356 17746 27384 18634
rect 27718 18524 28026 18533
rect 27718 18522 27724 18524
rect 27780 18522 27804 18524
rect 27860 18522 27884 18524
rect 27940 18522 27964 18524
rect 28020 18522 28026 18524
rect 27780 18470 27782 18522
rect 27962 18470 27964 18522
rect 27718 18468 27724 18470
rect 27780 18468 27804 18470
rect 27860 18468 27884 18470
rect 27940 18468 27964 18470
rect 28020 18468 28026 18470
rect 27718 18459 28026 18468
rect 27068 17740 27120 17746
rect 27068 17682 27120 17688
rect 27344 17740 27396 17746
rect 27344 17682 27396 17688
rect 27718 17436 28026 17445
rect 27718 17434 27724 17436
rect 27780 17434 27804 17436
rect 27860 17434 27884 17436
rect 27940 17434 27964 17436
rect 28020 17434 28026 17436
rect 27780 17382 27782 17434
rect 27962 17382 27964 17434
rect 27718 17380 27724 17382
rect 27780 17380 27804 17382
rect 27860 17380 27884 17382
rect 27940 17380 27964 17382
rect 28020 17380 28026 17382
rect 27718 17371 28026 17380
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 26988 15570 27016 16458
rect 27172 16250 27200 16594
rect 27718 16348 28026 16357
rect 27718 16346 27724 16348
rect 27780 16346 27804 16348
rect 27860 16346 27884 16348
rect 27940 16346 27964 16348
rect 28020 16346 28026 16348
rect 27780 16294 27782 16346
rect 27962 16294 27964 16346
rect 27718 16292 27724 16294
rect 27780 16292 27804 16294
rect 27860 16292 27884 16294
rect 27940 16292 27964 16294
rect 28020 16292 28026 16294
rect 27718 16283 28026 16292
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 26976 15564 27028 15570
rect 26976 15506 27028 15512
rect 26608 15360 26660 15366
rect 26608 15302 26660 15308
rect 27172 15162 27200 16186
rect 27718 15260 28026 15269
rect 27718 15258 27724 15260
rect 27780 15258 27804 15260
rect 27860 15258 27884 15260
rect 27940 15258 27964 15260
rect 28020 15258 28026 15260
rect 27780 15206 27782 15258
rect 27962 15206 27964 15258
rect 27718 15204 27724 15206
rect 27780 15204 27804 15206
rect 27860 15204 27884 15206
rect 27940 15204 27964 15206
rect 28020 15204 28026 15206
rect 27718 15195 28026 15204
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24372 14716 24680 14725
rect 24372 14714 24378 14716
rect 24434 14714 24458 14716
rect 24514 14714 24538 14716
rect 24594 14714 24618 14716
rect 24674 14714 24680 14716
rect 24434 14662 24436 14714
rect 24616 14662 24618 14714
rect 24372 14660 24378 14662
rect 24434 14660 24458 14662
rect 24514 14660 24538 14662
rect 24594 14660 24618 14662
rect 24674 14660 24680 14662
rect 24372 14651 24680 14660
rect 25332 14414 25360 14962
rect 25608 14414 25636 14962
rect 26436 14414 26464 15098
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 24044 13326 24072 14214
rect 25056 14074 25084 14350
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 24768 13728 24820 13734
rect 24768 13670 24820 13676
rect 24372 13628 24680 13637
rect 24372 13626 24378 13628
rect 24434 13626 24458 13628
rect 24514 13626 24538 13628
rect 24594 13626 24618 13628
rect 24674 13626 24680 13628
rect 24434 13574 24436 13626
rect 24616 13574 24618 13626
rect 24372 13572 24378 13574
rect 24434 13572 24458 13574
rect 24514 13572 24538 13574
rect 24594 13572 24618 13574
rect 24674 13572 24680 13574
rect 24372 13563 24680 13572
rect 24780 13530 24808 13670
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22204 11218 22232 11494
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 20272 10266 20300 10610
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 21008 10062 21036 10406
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 22020 9994 22048 10610
rect 22112 10198 22140 11086
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 22008 9988 22060 9994
rect 22008 9930 22060 9936
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9722 20576 9862
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19812 8634 19840 9522
rect 20548 9518 20576 9658
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20732 8974 20760 9318
rect 20824 9042 20852 9930
rect 21026 9820 21334 9829
rect 21026 9818 21032 9820
rect 21088 9818 21112 9820
rect 21168 9818 21192 9820
rect 21248 9818 21272 9820
rect 21328 9818 21334 9820
rect 21088 9766 21090 9818
rect 21270 9766 21272 9818
rect 21026 9764 21032 9766
rect 21088 9764 21112 9766
rect 21168 9764 21192 9766
rect 21248 9764 21272 9766
rect 21328 9764 21334 9766
rect 21026 9755 21334 9764
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21100 9178 21128 9318
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 22112 9042 22140 10134
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21026 8732 21334 8741
rect 21026 8730 21032 8732
rect 21088 8730 21112 8732
rect 21168 8730 21192 8732
rect 21248 8730 21272 8732
rect 21328 8730 21334 8732
rect 21088 8678 21090 8730
rect 21270 8678 21272 8730
rect 21026 8676 21032 8678
rect 21088 8676 21112 8678
rect 21168 8676 21192 8678
rect 21248 8676 21272 8678
rect 21328 8676 21334 8678
rect 21026 8667 21334 8676
rect 19800 8628 19852 8634
rect 19800 8570 19852 8576
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19708 8560 19760 8566
rect 19708 8502 19760 8508
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19536 8090 19564 8502
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 20824 7818 20852 8230
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18892 5370 18920 5578
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 9784 5086 9904 5114
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9876 4486 9904 5086
rect 9968 4690 9996 5170
rect 10796 4826 10824 5170
rect 10988 4924 11296 4933
rect 10988 4922 10994 4924
rect 11050 4922 11074 4924
rect 11130 4922 11154 4924
rect 11210 4922 11234 4924
rect 11290 4922 11296 4924
rect 11050 4870 11052 4922
rect 11232 4870 11234 4922
rect 10988 4868 10994 4870
rect 11050 4868 11074 4870
rect 11130 4868 11154 4870
rect 11210 4868 11234 4870
rect 11290 4868 11296 4870
rect 10988 4859 11296 4868
rect 17680 4924 17988 4933
rect 17680 4922 17686 4924
rect 17742 4922 17766 4924
rect 17822 4922 17846 4924
rect 17902 4922 17926 4924
rect 17982 4922 17988 4924
rect 17742 4870 17744 4922
rect 17924 4870 17926 4922
rect 17680 4868 17686 4870
rect 17742 4868 17766 4870
rect 17822 4868 17846 4870
rect 17902 4868 17926 4870
rect 17982 4868 17988 4870
rect 17680 4859 17988 4868
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 7642 4380 7950 4389
rect 7642 4378 7648 4380
rect 7704 4378 7728 4380
rect 7784 4378 7808 4380
rect 7864 4378 7888 4380
rect 7944 4378 7950 4380
rect 7704 4326 7706 4378
rect 7886 4326 7888 4378
rect 7642 4324 7648 4326
rect 7704 4324 7728 4326
rect 7784 4324 7808 4326
rect 7864 4324 7888 4326
rect 7944 4324 7950 4326
rect 7642 4315 7950 4324
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 9876 4010 9904 4422
rect 14334 4380 14642 4389
rect 14334 4378 14340 4380
rect 14396 4378 14420 4380
rect 14476 4378 14500 4380
rect 14556 4378 14580 4380
rect 14636 4378 14642 4380
rect 14396 4326 14398 4378
rect 14578 4326 14580 4378
rect 14334 4324 14340 4326
rect 14396 4324 14420 4326
rect 14476 4324 14500 4326
rect 14556 4324 14580 4326
rect 14636 4324 14642 4326
rect 14334 4315 14642 4324
rect 18892 4078 18920 5306
rect 18984 4146 19012 6394
rect 19352 6390 19380 6598
rect 19536 6458 19564 7346
rect 20180 7002 20208 7686
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19616 6384 19668 6390
rect 19616 6326 19668 6332
rect 19628 4146 19656 6326
rect 19720 5778 19748 6598
rect 19996 6458 20024 6734
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 20732 5642 20760 7278
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20824 5302 20852 7754
rect 21026 7644 21334 7653
rect 21026 7642 21032 7644
rect 21088 7642 21112 7644
rect 21168 7642 21192 7644
rect 21248 7642 21272 7644
rect 21328 7642 21334 7644
rect 21088 7590 21090 7642
rect 21270 7590 21272 7642
rect 21026 7588 21032 7590
rect 21088 7588 21112 7590
rect 21168 7588 21192 7590
rect 21248 7588 21272 7590
rect 21328 7588 21334 7590
rect 21026 7579 21334 7588
rect 21376 7410 21404 8434
rect 22020 8090 22048 8910
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6866 20944 7142
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21192 6730 21220 7346
rect 22296 6798 22324 8774
rect 22572 7546 22600 11698
rect 22756 11354 22784 11834
rect 23124 11558 23152 12242
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23216 11762 23244 12174
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23308 11354 23336 12854
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23400 12646 23428 12786
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23124 10130 23152 11154
rect 23308 11082 23336 11290
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23308 9926 23336 10406
rect 23400 9994 23428 12582
rect 24372 12540 24680 12549
rect 24372 12538 24378 12540
rect 24434 12538 24458 12540
rect 24514 12538 24538 12540
rect 24594 12538 24618 12540
rect 24674 12538 24680 12540
rect 24434 12486 24436 12538
rect 24616 12486 24618 12538
rect 24372 12484 24378 12486
rect 24434 12484 24458 12486
rect 24514 12484 24538 12486
rect 24594 12484 24618 12486
rect 24674 12484 24680 12486
rect 24372 12475 24680 12484
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24372 11452 24680 11461
rect 24372 11450 24378 11452
rect 24434 11450 24458 11452
rect 24514 11450 24538 11452
rect 24594 11450 24618 11452
rect 24674 11450 24680 11452
rect 24434 11398 24436 11450
rect 24616 11398 24618 11450
rect 24372 11396 24378 11398
rect 24434 11396 24458 11398
rect 24514 11396 24538 11398
rect 24594 11396 24618 11398
rect 24674 11396 24680 11398
rect 24372 11387 24680 11396
rect 24872 11218 24900 11494
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24372 10364 24680 10373
rect 24372 10362 24378 10364
rect 24434 10362 24458 10364
rect 24514 10362 24538 10364
rect 24594 10362 24618 10364
rect 24674 10362 24680 10364
rect 24434 10310 24436 10362
rect 24616 10310 24618 10362
rect 24372 10308 24378 10310
rect 24434 10308 24458 10310
rect 24514 10308 24538 10310
rect 24594 10308 24618 10310
rect 24674 10308 24680 10310
rect 24372 10299 24680 10308
rect 24780 10266 24808 11018
rect 24964 10810 24992 11018
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 25056 10690 25084 14010
rect 26344 14006 26372 14282
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25148 13326 25176 13806
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25148 12850 25176 13262
rect 25332 12986 25360 13262
rect 26620 13258 26648 14894
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26792 14340 26844 14346
rect 26792 14282 26844 14288
rect 26804 13394 26832 14282
rect 27080 13530 27108 14350
rect 27172 14074 27200 15098
rect 27718 14172 28026 14181
rect 27718 14170 27724 14172
rect 27780 14170 27804 14172
rect 27860 14170 27884 14172
rect 27940 14170 27964 14172
rect 28020 14170 28026 14172
rect 27780 14118 27782 14170
rect 27962 14118 27964 14170
rect 27718 14116 27724 14118
rect 27780 14116 27804 14118
rect 27860 14116 27884 14118
rect 27940 14116 27964 14118
rect 28020 14116 28026 14118
rect 27718 14107 28026 14116
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27068 13524 27120 13530
rect 27068 13466 27120 13472
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 26608 13252 26660 13258
rect 26608 13194 26660 13200
rect 27718 13084 28026 13093
rect 27718 13082 27724 13084
rect 27780 13082 27804 13084
rect 27860 13082 27884 13084
rect 27940 13082 27964 13084
rect 28020 13082 28026 13084
rect 27780 13030 27782 13082
rect 27962 13030 27964 13082
rect 27718 13028 27724 13030
rect 27780 13028 27804 13030
rect 27860 13028 27884 13030
rect 27940 13028 27964 13030
rect 28020 13028 28026 13030
rect 27718 13019 28026 13028
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 27718 11996 28026 12005
rect 27718 11994 27724 11996
rect 27780 11994 27804 11996
rect 27860 11994 27884 11996
rect 27940 11994 27964 11996
rect 28020 11994 28026 11996
rect 27780 11942 27782 11994
rect 27962 11942 27964 11994
rect 27718 11940 27724 11942
rect 27780 11940 27804 11942
rect 27860 11940 27884 11942
rect 27940 11940 27964 11942
rect 28020 11940 28026 11942
rect 27718 11931 28026 11940
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26344 11354 26372 11698
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 27718 10908 28026 10917
rect 27718 10906 27724 10908
rect 27780 10906 27804 10908
rect 27860 10906 27884 10908
rect 27940 10906 27964 10908
rect 28020 10906 28026 10908
rect 27780 10854 27782 10906
rect 27962 10854 27964 10906
rect 27718 10852 27724 10854
rect 27780 10852 27804 10854
rect 27860 10852 27884 10854
rect 27940 10852 27964 10854
rect 28020 10852 28026 10854
rect 27718 10843 28026 10852
rect 24964 10662 25084 10690
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25136 10668 25188 10674
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 23756 10056 23808 10062
rect 23756 9998 23808 10004
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22664 7818 22692 9522
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22848 9178 22876 9386
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22940 8566 22968 9862
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22928 8560 22980 8566
rect 22928 8502 22980 8508
rect 23032 8090 23060 9590
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23216 8974 23244 9522
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23216 8634 23244 8910
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23308 7954 23336 9862
rect 23768 9382 23796 9998
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23584 8566 23612 9318
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23768 7886 23796 9318
rect 24372 9276 24680 9285
rect 24372 9274 24378 9276
rect 24434 9274 24458 9276
rect 24514 9274 24538 9276
rect 24594 9274 24618 9276
rect 24674 9274 24680 9276
rect 24434 9222 24436 9274
rect 24616 9222 24618 9274
rect 24372 9220 24378 9222
rect 24434 9220 24458 9222
rect 24514 9220 24538 9222
rect 24594 9220 24618 9222
rect 24674 9220 24680 9222
rect 24372 9211 24680 9220
rect 24780 9042 24808 9590
rect 24964 9110 24992 10662
rect 25136 10610 25188 10616
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 25148 8974 25176 10610
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25240 9654 25268 9930
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25332 8974 25360 10678
rect 27718 9820 28026 9829
rect 27718 9818 27724 9820
rect 27780 9818 27804 9820
rect 27860 9818 27884 9820
rect 27940 9818 27964 9820
rect 28020 9818 28026 9820
rect 27780 9766 27782 9818
rect 27962 9766 27964 9818
rect 27718 9764 27724 9766
rect 27780 9764 27804 9766
rect 27860 9764 27884 9766
rect 27940 9764 27964 9766
rect 28020 9764 28026 9766
rect 27718 9755 28026 9764
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22664 6866 22692 7754
rect 23952 7546 23980 8366
rect 24372 8188 24680 8197
rect 24372 8186 24378 8188
rect 24434 8186 24458 8188
rect 24514 8186 24538 8188
rect 24594 8186 24618 8188
rect 24674 8186 24680 8188
rect 24434 8134 24436 8186
rect 24616 8134 24618 8186
rect 24372 8132 24378 8134
rect 24434 8132 24458 8134
rect 24514 8132 24538 8134
rect 24594 8132 24618 8134
rect 24674 8132 24680 8134
rect 24372 8123 24680 8132
rect 24780 7954 24808 8366
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 25148 7886 25176 8910
rect 25516 8634 25544 9454
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 26160 8090 26188 8910
rect 27718 8732 28026 8741
rect 27718 8730 27724 8732
rect 27780 8730 27804 8732
rect 27860 8730 27884 8732
rect 27940 8730 27964 8732
rect 28020 8730 28026 8732
rect 27780 8678 27782 8730
rect 27962 8678 27964 8730
rect 27718 8676 27724 8678
rect 27780 8676 27804 8678
rect 27860 8676 27884 8678
rect 27940 8676 27964 8678
rect 28020 8676 28026 8678
rect 27718 8667 28026 8676
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26160 7886 26188 8026
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 21180 6724 21232 6730
rect 21180 6666 21232 6672
rect 20916 5914 20944 6666
rect 21026 6556 21334 6565
rect 21026 6554 21032 6556
rect 21088 6554 21112 6556
rect 21168 6554 21192 6556
rect 21248 6554 21272 6556
rect 21328 6554 21334 6556
rect 21088 6502 21090 6554
rect 21270 6502 21272 6554
rect 21026 6500 21032 6502
rect 21088 6500 21112 6502
rect 21168 6500 21192 6502
rect 21248 6500 21272 6502
rect 21328 6500 21334 6502
rect 21026 6491 21334 6500
rect 22848 6458 22876 7414
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24412 7206 24440 7278
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 23492 6866 23520 7142
rect 24372 7100 24680 7109
rect 24372 7098 24378 7100
rect 24434 7098 24458 7100
rect 24514 7098 24538 7100
rect 24594 7098 24618 7100
rect 24674 7098 24680 7100
rect 24434 7046 24436 7098
rect 24616 7046 24618 7098
rect 24372 7044 24378 7046
rect 24434 7044 24458 7046
rect 24514 7044 24538 7046
rect 24594 7044 24618 7046
rect 24674 7044 24680 7046
rect 24372 7035 24680 7044
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 25148 6322 25176 7822
rect 25240 6390 25268 7822
rect 27718 7644 28026 7653
rect 27718 7642 27724 7644
rect 27780 7642 27804 7644
rect 27860 7642 27884 7644
rect 27940 7642 27964 7644
rect 28020 7642 28026 7644
rect 27780 7590 27782 7642
rect 27962 7590 27964 7642
rect 27718 7588 27724 7590
rect 27780 7588 27804 7590
rect 27860 7588 27884 7590
rect 27940 7588 27964 7590
rect 28020 7588 28026 7590
rect 27718 7579 28026 7588
rect 27718 6556 28026 6565
rect 27718 6554 27724 6556
rect 27780 6554 27804 6556
rect 27860 6554 27884 6556
rect 27940 6554 27964 6556
rect 28020 6554 28026 6556
rect 27780 6502 27782 6554
rect 27962 6502 27964 6554
rect 27718 6500 27724 6502
rect 27780 6500 27804 6502
rect 27860 6500 27884 6502
rect 27940 6500 27964 6502
rect 28020 6500 28026 6502
rect 27718 6491 28026 6500
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 24372 6012 24680 6021
rect 24372 6010 24378 6012
rect 24434 6010 24458 6012
rect 24514 6010 24538 6012
rect 24594 6010 24618 6012
rect 24674 6010 24680 6012
rect 24434 5958 24436 6010
rect 24616 5958 24618 6010
rect 24372 5956 24378 5958
rect 24434 5956 24458 5958
rect 24514 5956 24538 5958
rect 24594 5956 24618 5958
rect 24674 5956 24680 5958
rect 24372 5947 24680 5956
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21026 5468 21334 5477
rect 21026 5466 21032 5468
rect 21088 5466 21112 5468
rect 21168 5466 21192 5468
rect 21248 5466 21272 5468
rect 21328 5466 21334 5468
rect 21088 5414 21090 5466
rect 21270 5414 21272 5466
rect 21026 5412 21032 5414
rect 21088 5412 21112 5414
rect 21168 5412 21192 5414
rect 21248 5412 21272 5414
rect 21328 5412 21334 5414
rect 21026 5403 21334 5412
rect 27718 5468 28026 5477
rect 27718 5466 27724 5468
rect 27780 5466 27804 5468
rect 27860 5466 27884 5468
rect 27940 5466 27964 5468
rect 28020 5466 28026 5468
rect 27780 5414 27782 5466
rect 27962 5414 27964 5466
rect 27718 5412 27724 5414
rect 27780 5412 27804 5414
rect 27860 5412 27884 5414
rect 27940 5412 27964 5414
rect 28020 5412 28026 5414
rect 27718 5403 28026 5412
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 24372 4924 24680 4933
rect 24372 4922 24378 4924
rect 24434 4922 24458 4924
rect 24514 4922 24538 4924
rect 24594 4922 24618 4924
rect 24674 4922 24680 4924
rect 24434 4870 24436 4922
rect 24616 4870 24618 4922
rect 24372 4868 24378 4870
rect 24434 4868 24458 4870
rect 24514 4868 24538 4870
rect 24594 4868 24618 4870
rect 24674 4868 24680 4870
rect 24372 4859 24680 4868
rect 21026 4380 21334 4389
rect 21026 4378 21032 4380
rect 21088 4378 21112 4380
rect 21168 4378 21192 4380
rect 21248 4378 21272 4380
rect 21328 4378 21334 4380
rect 21088 4326 21090 4378
rect 21270 4326 21272 4378
rect 21026 4324 21032 4326
rect 21088 4324 21112 4326
rect 21168 4324 21192 4326
rect 21248 4324 21272 4326
rect 21328 4324 21334 4326
rect 21026 4315 21334 4324
rect 27718 4380 28026 4389
rect 27718 4378 27724 4380
rect 27780 4378 27804 4380
rect 27860 4378 27884 4380
rect 27940 4378 27964 4380
rect 28020 4378 28026 4380
rect 27780 4326 27782 4378
rect 27962 4326 27964 4378
rect 27718 4324 27724 4326
rect 27780 4324 27804 4326
rect 27860 4324 27884 4326
rect 27940 4324 27964 4326
rect 28020 4324 28026 4326
rect 27718 4315 28026 4324
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5184 3194 5212 3470
rect 5736 3194 5764 3674
rect 7642 3292 7950 3301
rect 7642 3290 7648 3292
rect 7704 3290 7728 3292
rect 7784 3290 7808 3292
rect 7864 3290 7888 3292
rect 7944 3290 7950 3292
rect 7704 3238 7706 3290
rect 7886 3238 7888 3290
rect 7642 3236 7648 3238
rect 7704 3236 7728 3238
rect 7784 3236 7808 3238
rect 7864 3236 7888 3238
rect 7944 3236 7950 3238
rect 7642 3227 7950 3236
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4296 2748 4604 2757
rect 4296 2746 4302 2748
rect 4358 2746 4382 2748
rect 4438 2746 4462 2748
rect 4518 2746 4542 2748
rect 4598 2746 4604 2748
rect 4358 2694 4360 2746
rect 4540 2694 4542 2746
rect 4296 2692 4302 2694
rect 4358 2692 4382 2694
rect 4438 2692 4462 2694
rect 4518 2692 4542 2694
rect 4598 2692 4604 2694
rect 4296 2683 4604 2692
rect 5736 2650 5764 3130
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 3792 2576 3844 2582
rect 3792 2518 3844 2524
rect 5736 2514 5764 2586
rect 8128 2582 8156 3878
rect 10988 3836 11296 3845
rect 10988 3834 10994 3836
rect 11050 3834 11074 3836
rect 11130 3834 11154 3836
rect 11210 3834 11234 3836
rect 11290 3834 11296 3836
rect 11050 3782 11052 3834
rect 11232 3782 11234 3834
rect 10988 3780 10994 3782
rect 11050 3780 11074 3782
rect 11130 3780 11154 3782
rect 11210 3780 11234 3782
rect 11290 3780 11296 3782
rect 10988 3771 11296 3780
rect 17680 3836 17988 3845
rect 17680 3834 17686 3836
rect 17742 3834 17766 3836
rect 17822 3834 17846 3836
rect 17902 3834 17926 3836
rect 17982 3834 17988 3836
rect 17742 3782 17744 3834
rect 17924 3782 17926 3834
rect 17680 3780 17686 3782
rect 17742 3780 17766 3782
rect 17822 3780 17846 3782
rect 17902 3780 17926 3782
rect 17982 3780 17988 3782
rect 17680 3771 17988 3780
rect 24372 3836 24680 3845
rect 24372 3834 24378 3836
rect 24434 3834 24458 3836
rect 24514 3834 24538 3836
rect 24594 3834 24618 3836
rect 24674 3834 24680 3836
rect 24434 3782 24436 3834
rect 24616 3782 24618 3834
rect 24372 3780 24378 3782
rect 24434 3780 24458 3782
rect 24514 3780 24538 3782
rect 24594 3780 24618 3782
rect 24674 3780 24680 3782
rect 24372 3771 24680 3780
rect 14334 3292 14642 3301
rect 14334 3290 14340 3292
rect 14396 3290 14420 3292
rect 14476 3290 14500 3292
rect 14556 3290 14580 3292
rect 14636 3290 14642 3292
rect 14396 3238 14398 3290
rect 14578 3238 14580 3290
rect 14334 3236 14340 3238
rect 14396 3236 14420 3238
rect 14476 3236 14500 3238
rect 14556 3236 14580 3238
rect 14636 3236 14642 3238
rect 14334 3227 14642 3236
rect 21026 3292 21334 3301
rect 21026 3290 21032 3292
rect 21088 3290 21112 3292
rect 21168 3290 21192 3292
rect 21248 3290 21272 3292
rect 21328 3290 21334 3292
rect 21088 3238 21090 3290
rect 21270 3238 21272 3290
rect 21026 3236 21032 3238
rect 21088 3236 21112 3238
rect 21168 3236 21192 3238
rect 21248 3236 21272 3238
rect 21328 3236 21334 3238
rect 21026 3227 21334 3236
rect 27718 3292 28026 3301
rect 27718 3290 27724 3292
rect 27780 3290 27804 3292
rect 27860 3290 27884 3292
rect 27940 3290 27964 3292
rect 28020 3290 28026 3292
rect 27780 3238 27782 3290
rect 27962 3238 27964 3290
rect 27718 3236 27724 3238
rect 27780 3236 27804 3238
rect 27860 3236 27884 3238
rect 27940 3236 27964 3238
rect 28020 3236 28026 3238
rect 27718 3227 28026 3236
rect 10988 2748 11296 2757
rect 10988 2746 10994 2748
rect 11050 2746 11074 2748
rect 11130 2746 11154 2748
rect 11210 2746 11234 2748
rect 11290 2746 11296 2748
rect 11050 2694 11052 2746
rect 11232 2694 11234 2746
rect 10988 2692 10994 2694
rect 11050 2692 11074 2694
rect 11130 2692 11154 2694
rect 11210 2692 11234 2694
rect 11290 2692 11296 2694
rect 10988 2683 11296 2692
rect 17680 2748 17988 2757
rect 17680 2746 17686 2748
rect 17742 2746 17766 2748
rect 17822 2746 17846 2748
rect 17902 2746 17926 2748
rect 17982 2746 17988 2748
rect 17742 2694 17744 2746
rect 17924 2694 17926 2746
rect 17680 2692 17686 2694
rect 17742 2692 17766 2694
rect 17822 2692 17846 2694
rect 17902 2692 17926 2694
rect 17982 2692 17988 2694
rect 17680 2683 17988 2692
rect 24372 2748 24680 2757
rect 24372 2746 24378 2748
rect 24434 2746 24458 2748
rect 24514 2746 24538 2748
rect 24594 2746 24618 2748
rect 24674 2746 24680 2748
rect 24434 2694 24436 2746
rect 24616 2694 24618 2746
rect 24372 2692 24378 2694
rect 24434 2692 24458 2694
rect 24514 2692 24538 2694
rect 24594 2692 24618 2694
rect 24674 2692 24680 2694
rect 24372 2683 24680 2692
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 2145 3280 2246
rect 7642 2204 7950 2213
rect 7642 2202 7648 2204
rect 7704 2202 7728 2204
rect 7784 2202 7808 2204
rect 7864 2202 7888 2204
rect 7944 2202 7950 2204
rect 7704 2150 7706 2202
rect 7886 2150 7888 2202
rect 7642 2148 7648 2150
rect 7704 2148 7728 2150
rect 7784 2148 7808 2150
rect 7864 2148 7888 2150
rect 7944 2148 7950 2150
rect 3238 2136 3294 2145
rect 7642 2139 7950 2148
rect 14334 2204 14642 2213
rect 14334 2202 14340 2204
rect 14396 2202 14420 2204
rect 14476 2202 14500 2204
rect 14556 2202 14580 2204
rect 14636 2202 14642 2204
rect 14396 2150 14398 2202
rect 14578 2150 14580 2202
rect 14334 2148 14340 2150
rect 14396 2148 14420 2150
rect 14476 2148 14500 2150
rect 14556 2148 14580 2150
rect 14636 2148 14642 2150
rect 14334 2139 14642 2148
rect 21026 2204 21334 2213
rect 21026 2202 21032 2204
rect 21088 2202 21112 2204
rect 21168 2202 21192 2204
rect 21248 2202 21272 2204
rect 21328 2202 21334 2204
rect 21088 2150 21090 2202
rect 21270 2150 21272 2202
rect 21026 2148 21032 2150
rect 21088 2148 21112 2150
rect 21168 2148 21192 2150
rect 21248 2148 21272 2150
rect 21328 2148 21334 2150
rect 21026 2139 21334 2148
rect 27718 2204 28026 2213
rect 27718 2202 27724 2204
rect 27780 2202 27804 2204
rect 27860 2202 27884 2204
rect 27940 2202 27964 2204
rect 28020 2202 28026 2204
rect 27780 2150 27782 2202
rect 27962 2150 27964 2202
rect 27718 2148 27724 2150
rect 27780 2148 27804 2150
rect 27860 2148 27884 2150
rect 27940 2148 27964 2150
rect 28020 2148 28026 2150
rect 27718 2139 28026 2148
rect 3238 2071 3294 2080
<< via2 >>
rect 1674 26832 1730 26888
rect 4302 26682 4358 26684
rect 4382 26682 4438 26684
rect 4462 26682 4518 26684
rect 4542 26682 4598 26684
rect 4302 26630 4348 26682
rect 4348 26630 4358 26682
rect 4382 26630 4412 26682
rect 4412 26630 4424 26682
rect 4424 26630 4438 26682
rect 4462 26630 4476 26682
rect 4476 26630 4488 26682
rect 4488 26630 4518 26682
rect 4542 26630 4552 26682
rect 4552 26630 4598 26682
rect 4302 26628 4358 26630
rect 4382 26628 4438 26630
rect 4462 26628 4518 26630
rect 4542 26628 4598 26630
rect 10994 26682 11050 26684
rect 11074 26682 11130 26684
rect 11154 26682 11210 26684
rect 11234 26682 11290 26684
rect 10994 26630 11040 26682
rect 11040 26630 11050 26682
rect 11074 26630 11104 26682
rect 11104 26630 11116 26682
rect 11116 26630 11130 26682
rect 11154 26630 11168 26682
rect 11168 26630 11180 26682
rect 11180 26630 11210 26682
rect 11234 26630 11244 26682
rect 11244 26630 11290 26682
rect 10994 26628 11050 26630
rect 11074 26628 11130 26630
rect 11154 26628 11210 26630
rect 11234 26628 11290 26630
rect 4302 25594 4358 25596
rect 4382 25594 4438 25596
rect 4462 25594 4518 25596
rect 4542 25594 4598 25596
rect 4302 25542 4348 25594
rect 4348 25542 4358 25594
rect 4382 25542 4412 25594
rect 4412 25542 4424 25594
rect 4424 25542 4438 25594
rect 4462 25542 4476 25594
rect 4476 25542 4488 25594
rect 4488 25542 4518 25594
rect 4542 25542 4552 25594
rect 4552 25542 4598 25594
rect 4302 25540 4358 25542
rect 4382 25540 4438 25542
rect 4462 25540 4518 25542
rect 4542 25540 4598 25542
rect 4302 24506 4358 24508
rect 4382 24506 4438 24508
rect 4462 24506 4518 24508
rect 4542 24506 4598 24508
rect 4302 24454 4348 24506
rect 4348 24454 4358 24506
rect 4382 24454 4412 24506
rect 4412 24454 4424 24506
rect 4424 24454 4438 24506
rect 4462 24454 4476 24506
rect 4476 24454 4488 24506
rect 4488 24454 4518 24506
rect 4542 24454 4552 24506
rect 4552 24454 4598 24506
rect 4302 24452 4358 24454
rect 4382 24452 4438 24454
rect 4462 24452 4518 24454
rect 4542 24452 4598 24454
rect 3514 23296 3570 23352
rect 4302 23418 4358 23420
rect 4382 23418 4438 23420
rect 4462 23418 4518 23420
rect 4542 23418 4598 23420
rect 4302 23366 4348 23418
rect 4348 23366 4358 23418
rect 4382 23366 4412 23418
rect 4412 23366 4424 23418
rect 4424 23366 4438 23418
rect 4462 23366 4476 23418
rect 4476 23366 4488 23418
rect 4488 23366 4518 23418
rect 4542 23366 4552 23418
rect 4552 23366 4598 23418
rect 4302 23364 4358 23366
rect 4382 23364 4438 23366
rect 4462 23364 4518 23366
rect 4542 23364 4598 23366
rect 4302 22330 4358 22332
rect 4382 22330 4438 22332
rect 4462 22330 4518 22332
rect 4542 22330 4598 22332
rect 4302 22278 4348 22330
rect 4348 22278 4358 22330
rect 4382 22278 4412 22330
rect 4412 22278 4424 22330
rect 4424 22278 4438 22330
rect 4462 22278 4476 22330
rect 4476 22278 4488 22330
rect 4488 22278 4518 22330
rect 4542 22278 4552 22330
rect 4552 22278 4598 22330
rect 4302 22276 4358 22278
rect 4382 22276 4438 22278
rect 4462 22276 4518 22278
rect 4542 22276 4598 22278
rect 1674 19760 1730 19816
rect 4302 21242 4358 21244
rect 4382 21242 4438 21244
rect 4462 21242 4518 21244
rect 4542 21242 4598 21244
rect 4302 21190 4348 21242
rect 4348 21190 4358 21242
rect 4382 21190 4412 21242
rect 4412 21190 4424 21242
rect 4424 21190 4438 21242
rect 4462 21190 4476 21242
rect 4476 21190 4488 21242
rect 4488 21190 4518 21242
rect 4542 21190 4552 21242
rect 4552 21190 4598 21242
rect 4302 21188 4358 21190
rect 4382 21188 4438 21190
rect 4462 21188 4518 21190
rect 4542 21188 4598 21190
rect 4302 20154 4358 20156
rect 4382 20154 4438 20156
rect 4462 20154 4518 20156
rect 4542 20154 4598 20156
rect 4302 20102 4348 20154
rect 4348 20102 4358 20154
rect 4382 20102 4412 20154
rect 4412 20102 4424 20154
rect 4424 20102 4438 20154
rect 4462 20102 4476 20154
rect 4476 20102 4488 20154
rect 4488 20102 4518 20154
rect 4542 20102 4552 20154
rect 4552 20102 4598 20154
rect 4302 20100 4358 20102
rect 4382 20100 4438 20102
rect 4462 20100 4518 20102
rect 4542 20100 4598 20102
rect 4302 19066 4358 19068
rect 4382 19066 4438 19068
rect 4462 19066 4518 19068
rect 4542 19066 4598 19068
rect 4302 19014 4348 19066
rect 4348 19014 4358 19066
rect 4382 19014 4412 19066
rect 4412 19014 4424 19066
rect 4424 19014 4438 19066
rect 4462 19014 4476 19066
rect 4476 19014 4488 19066
rect 4488 19014 4518 19066
rect 4542 19014 4552 19066
rect 4552 19014 4598 19066
rect 4302 19012 4358 19014
rect 4382 19012 4438 19014
rect 4462 19012 4518 19014
rect 4542 19012 4598 19014
rect 1582 16224 1638 16280
rect 1582 12688 1638 12744
rect 1490 5616 1546 5672
rect 2962 9152 3018 9208
rect 4302 17978 4358 17980
rect 4382 17978 4438 17980
rect 4462 17978 4518 17980
rect 4542 17978 4598 17980
rect 4302 17926 4348 17978
rect 4348 17926 4358 17978
rect 4382 17926 4412 17978
rect 4412 17926 4424 17978
rect 4424 17926 4438 17978
rect 4462 17926 4476 17978
rect 4476 17926 4488 17978
rect 4488 17926 4518 17978
rect 4542 17926 4552 17978
rect 4552 17926 4598 17978
rect 4302 17924 4358 17926
rect 4382 17924 4438 17926
rect 4462 17924 4518 17926
rect 4542 17924 4598 17926
rect 4302 16890 4358 16892
rect 4382 16890 4438 16892
rect 4462 16890 4518 16892
rect 4542 16890 4598 16892
rect 4302 16838 4348 16890
rect 4348 16838 4358 16890
rect 4382 16838 4412 16890
rect 4412 16838 4424 16890
rect 4424 16838 4438 16890
rect 4462 16838 4476 16890
rect 4476 16838 4488 16890
rect 4488 16838 4518 16890
rect 4542 16838 4552 16890
rect 4552 16838 4598 16890
rect 4302 16836 4358 16838
rect 4382 16836 4438 16838
rect 4462 16836 4518 16838
rect 4542 16836 4598 16838
rect 7648 26138 7704 26140
rect 7728 26138 7784 26140
rect 7808 26138 7864 26140
rect 7888 26138 7944 26140
rect 7648 26086 7694 26138
rect 7694 26086 7704 26138
rect 7728 26086 7758 26138
rect 7758 26086 7770 26138
rect 7770 26086 7784 26138
rect 7808 26086 7822 26138
rect 7822 26086 7834 26138
rect 7834 26086 7864 26138
rect 7888 26086 7898 26138
rect 7898 26086 7944 26138
rect 7648 26084 7704 26086
rect 7728 26084 7784 26086
rect 7808 26084 7864 26086
rect 7888 26084 7944 26086
rect 7648 25050 7704 25052
rect 7728 25050 7784 25052
rect 7808 25050 7864 25052
rect 7888 25050 7944 25052
rect 7648 24998 7694 25050
rect 7694 24998 7704 25050
rect 7728 24998 7758 25050
rect 7758 24998 7770 25050
rect 7770 24998 7784 25050
rect 7808 24998 7822 25050
rect 7822 24998 7834 25050
rect 7834 24998 7864 25050
rect 7888 24998 7898 25050
rect 7898 24998 7944 25050
rect 7648 24996 7704 24998
rect 7728 24996 7784 24998
rect 7808 24996 7864 24998
rect 7888 24996 7944 24998
rect 4302 15802 4358 15804
rect 4382 15802 4438 15804
rect 4462 15802 4518 15804
rect 4542 15802 4598 15804
rect 4302 15750 4348 15802
rect 4348 15750 4358 15802
rect 4382 15750 4412 15802
rect 4412 15750 4424 15802
rect 4424 15750 4438 15802
rect 4462 15750 4476 15802
rect 4476 15750 4488 15802
rect 4488 15750 4518 15802
rect 4542 15750 4552 15802
rect 4552 15750 4598 15802
rect 4302 15748 4358 15750
rect 4382 15748 4438 15750
rect 4462 15748 4518 15750
rect 4542 15748 4598 15750
rect 4302 14714 4358 14716
rect 4382 14714 4438 14716
rect 4462 14714 4518 14716
rect 4542 14714 4598 14716
rect 4302 14662 4348 14714
rect 4348 14662 4358 14714
rect 4382 14662 4412 14714
rect 4412 14662 4424 14714
rect 4424 14662 4438 14714
rect 4462 14662 4476 14714
rect 4476 14662 4488 14714
rect 4488 14662 4518 14714
rect 4542 14662 4552 14714
rect 4552 14662 4598 14714
rect 4302 14660 4358 14662
rect 4382 14660 4438 14662
rect 4462 14660 4518 14662
rect 4542 14660 4598 14662
rect 4302 13626 4358 13628
rect 4382 13626 4438 13628
rect 4462 13626 4518 13628
rect 4542 13626 4598 13628
rect 4302 13574 4348 13626
rect 4348 13574 4358 13626
rect 4382 13574 4412 13626
rect 4412 13574 4424 13626
rect 4424 13574 4438 13626
rect 4462 13574 4476 13626
rect 4476 13574 4488 13626
rect 4488 13574 4518 13626
rect 4542 13574 4552 13626
rect 4552 13574 4598 13626
rect 4302 13572 4358 13574
rect 4382 13572 4438 13574
rect 4462 13572 4518 13574
rect 4542 13572 4598 13574
rect 4302 12538 4358 12540
rect 4382 12538 4438 12540
rect 4462 12538 4518 12540
rect 4542 12538 4598 12540
rect 4302 12486 4348 12538
rect 4348 12486 4358 12538
rect 4382 12486 4412 12538
rect 4412 12486 4424 12538
rect 4424 12486 4438 12538
rect 4462 12486 4476 12538
rect 4476 12486 4488 12538
rect 4488 12486 4518 12538
rect 4542 12486 4552 12538
rect 4552 12486 4598 12538
rect 4302 12484 4358 12486
rect 4382 12484 4438 12486
rect 4462 12484 4518 12486
rect 4542 12484 4598 12486
rect 4302 11450 4358 11452
rect 4382 11450 4438 11452
rect 4462 11450 4518 11452
rect 4542 11450 4598 11452
rect 4302 11398 4348 11450
rect 4348 11398 4358 11450
rect 4382 11398 4412 11450
rect 4412 11398 4424 11450
rect 4424 11398 4438 11450
rect 4462 11398 4476 11450
rect 4476 11398 4488 11450
rect 4488 11398 4518 11450
rect 4542 11398 4552 11450
rect 4552 11398 4598 11450
rect 4302 11396 4358 11398
rect 4382 11396 4438 11398
rect 4462 11396 4518 11398
rect 4542 11396 4598 11398
rect 7648 23962 7704 23964
rect 7728 23962 7784 23964
rect 7808 23962 7864 23964
rect 7888 23962 7944 23964
rect 7648 23910 7694 23962
rect 7694 23910 7704 23962
rect 7728 23910 7758 23962
rect 7758 23910 7770 23962
rect 7770 23910 7784 23962
rect 7808 23910 7822 23962
rect 7822 23910 7834 23962
rect 7834 23910 7864 23962
rect 7888 23910 7898 23962
rect 7898 23910 7944 23962
rect 7648 23908 7704 23910
rect 7728 23908 7784 23910
rect 7808 23908 7864 23910
rect 7888 23908 7944 23910
rect 7648 22874 7704 22876
rect 7728 22874 7784 22876
rect 7808 22874 7864 22876
rect 7888 22874 7944 22876
rect 7648 22822 7694 22874
rect 7694 22822 7704 22874
rect 7728 22822 7758 22874
rect 7758 22822 7770 22874
rect 7770 22822 7784 22874
rect 7808 22822 7822 22874
rect 7822 22822 7834 22874
rect 7834 22822 7864 22874
rect 7888 22822 7898 22874
rect 7898 22822 7944 22874
rect 7648 22820 7704 22822
rect 7728 22820 7784 22822
rect 7808 22820 7864 22822
rect 7888 22820 7944 22822
rect 7648 21786 7704 21788
rect 7728 21786 7784 21788
rect 7808 21786 7864 21788
rect 7888 21786 7944 21788
rect 7648 21734 7694 21786
rect 7694 21734 7704 21786
rect 7728 21734 7758 21786
rect 7758 21734 7770 21786
rect 7770 21734 7784 21786
rect 7808 21734 7822 21786
rect 7822 21734 7834 21786
rect 7834 21734 7864 21786
rect 7888 21734 7898 21786
rect 7898 21734 7944 21786
rect 7648 21732 7704 21734
rect 7728 21732 7784 21734
rect 7808 21732 7864 21734
rect 7888 21732 7944 21734
rect 10994 25594 11050 25596
rect 11074 25594 11130 25596
rect 11154 25594 11210 25596
rect 11234 25594 11290 25596
rect 10994 25542 11040 25594
rect 11040 25542 11050 25594
rect 11074 25542 11104 25594
rect 11104 25542 11116 25594
rect 11116 25542 11130 25594
rect 11154 25542 11168 25594
rect 11168 25542 11180 25594
rect 11180 25542 11210 25594
rect 11234 25542 11244 25594
rect 11244 25542 11290 25594
rect 10994 25540 11050 25542
rect 11074 25540 11130 25542
rect 11154 25540 11210 25542
rect 11234 25540 11290 25542
rect 10994 24506 11050 24508
rect 11074 24506 11130 24508
rect 11154 24506 11210 24508
rect 11234 24506 11290 24508
rect 10994 24454 11040 24506
rect 11040 24454 11050 24506
rect 11074 24454 11104 24506
rect 11104 24454 11116 24506
rect 11116 24454 11130 24506
rect 11154 24454 11168 24506
rect 11168 24454 11180 24506
rect 11180 24454 11210 24506
rect 11234 24454 11244 24506
rect 11244 24454 11290 24506
rect 10994 24452 11050 24454
rect 11074 24452 11130 24454
rect 11154 24452 11210 24454
rect 11234 24452 11290 24454
rect 7648 20698 7704 20700
rect 7728 20698 7784 20700
rect 7808 20698 7864 20700
rect 7888 20698 7944 20700
rect 7648 20646 7694 20698
rect 7694 20646 7704 20698
rect 7728 20646 7758 20698
rect 7758 20646 7770 20698
rect 7770 20646 7784 20698
rect 7808 20646 7822 20698
rect 7822 20646 7834 20698
rect 7834 20646 7864 20698
rect 7888 20646 7898 20698
rect 7898 20646 7944 20698
rect 7648 20644 7704 20646
rect 7728 20644 7784 20646
rect 7808 20644 7864 20646
rect 7888 20644 7944 20646
rect 7648 19610 7704 19612
rect 7728 19610 7784 19612
rect 7808 19610 7864 19612
rect 7888 19610 7944 19612
rect 7648 19558 7694 19610
rect 7694 19558 7704 19610
rect 7728 19558 7758 19610
rect 7758 19558 7770 19610
rect 7770 19558 7784 19610
rect 7808 19558 7822 19610
rect 7822 19558 7834 19610
rect 7834 19558 7864 19610
rect 7888 19558 7898 19610
rect 7898 19558 7944 19610
rect 7648 19556 7704 19558
rect 7728 19556 7784 19558
rect 7808 19556 7864 19558
rect 7888 19556 7944 19558
rect 7648 18522 7704 18524
rect 7728 18522 7784 18524
rect 7808 18522 7864 18524
rect 7888 18522 7944 18524
rect 7648 18470 7694 18522
rect 7694 18470 7704 18522
rect 7728 18470 7758 18522
rect 7758 18470 7770 18522
rect 7770 18470 7784 18522
rect 7808 18470 7822 18522
rect 7822 18470 7834 18522
rect 7834 18470 7864 18522
rect 7888 18470 7898 18522
rect 7898 18470 7944 18522
rect 7648 18468 7704 18470
rect 7728 18468 7784 18470
rect 7808 18468 7864 18470
rect 7888 18468 7944 18470
rect 7648 17434 7704 17436
rect 7728 17434 7784 17436
rect 7808 17434 7864 17436
rect 7888 17434 7944 17436
rect 7648 17382 7694 17434
rect 7694 17382 7704 17434
rect 7728 17382 7758 17434
rect 7758 17382 7770 17434
rect 7770 17382 7784 17434
rect 7808 17382 7822 17434
rect 7822 17382 7834 17434
rect 7834 17382 7864 17434
rect 7888 17382 7898 17434
rect 7898 17382 7944 17434
rect 7648 17380 7704 17382
rect 7728 17380 7784 17382
rect 7808 17380 7864 17382
rect 7888 17380 7944 17382
rect 7648 16346 7704 16348
rect 7728 16346 7784 16348
rect 7808 16346 7864 16348
rect 7888 16346 7944 16348
rect 7648 16294 7694 16346
rect 7694 16294 7704 16346
rect 7728 16294 7758 16346
rect 7758 16294 7770 16346
rect 7770 16294 7784 16346
rect 7808 16294 7822 16346
rect 7822 16294 7834 16346
rect 7834 16294 7864 16346
rect 7888 16294 7898 16346
rect 7898 16294 7944 16346
rect 7648 16292 7704 16294
rect 7728 16292 7784 16294
rect 7808 16292 7864 16294
rect 7888 16292 7944 16294
rect 7648 15258 7704 15260
rect 7728 15258 7784 15260
rect 7808 15258 7864 15260
rect 7888 15258 7944 15260
rect 7648 15206 7694 15258
rect 7694 15206 7704 15258
rect 7728 15206 7758 15258
rect 7758 15206 7770 15258
rect 7770 15206 7784 15258
rect 7808 15206 7822 15258
rect 7822 15206 7834 15258
rect 7834 15206 7864 15258
rect 7888 15206 7898 15258
rect 7898 15206 7944 15258
rect 7648 15204 7704 15206
rect 7728 15204 7784 15206
rect 7808 15204 7864 15206
rect 7888 15204 7944 15206
rect 4302 10362 4358 10364
rect 4382 10362 4438 10364
rect 4462 10362 4518 10364
rect 4542 10362 4598 10364
rect 4302 10310 4348 10362
rect 4348 10310 4358 10362
rect 4382 10310 4412 10362
rect 4412 10310 4424 10362
rect 4424 10310 4438 10362
rect 4462 10310 4476 10362
rect 4476 10310 4488 10362
rect 4488 10310 4518 10362
rect 4542 10310 4552 10362
rect 4552 10310 4598 10362
rect 4302 10308 4358 10310
rect 4382 10308 4438 10310
rect 4462 10308 4518 10310
rect 4542 10308 4598 10310
rect 4302 9274 4358 9276
rect 4382 9274 4438 9276
rect 4462 9274 4518 9276
rect 4542 9274 4598 9276
rect 4302 9222 4348 9274
rect 4348 9222 4358 9274
rect 4382 9222 4412 9274
rect 4412 9222 4424 9274
rect 4424 9222 4438 9274
rect 4462 9222 4476 9274
rect 4476 9222 4488 9274
rect 4488 9222 4518 9274
rect 4542 9222 4552 9274
rect 4552 9222 4598 9274
rect 4302 9220 4358 9222
rect 4382 9220 4438 9222
rect 4462 9220 4518 9222
rect 4542 9220 4598 9222
rect 4302 8186 4358 8188
rect 4382 8186 4438 8188
rect 4462 8186 4518 8188
rect 4542 8186 4598 8188
rect 4302 8134 4348 8186
rect 4348 8134 4358 8186
rect 4382 8134 4412 8186
rect 4412 8134 4424 8186
rect 4424 8134 4438 8186
rect 4462 8134 4476 8186
rect 4476 8134 4488 8186
rect 4488 8134 4518 8186
rect 4542 8134 4552 8186
rect 4552 8134 4598 8186
rect 4302 8132 4358 8134
rect 4382 8132 4438 8134
rect 4462 8132 4518 8134
rect 4542 8132 4598 8134
rect 4302 7098 4358 7100
rect 4382 7098 4438 7100
rect 4462 7098 4518 7100
rect 4542 7098 4598 7100
rect 4302 7046 4348 7098
rect 4348 7046 4358 7098
rect 4382 7046 4412 7098
rect 4412 7046 4424 7098
rect 4424 7046 4438 7098
rect 4462 7046 4476 7098
rect 4476 7046 4488 7098
rect 4488 7046 4518 7098
rect 4542 7046 4552 7098
rect 4552 7046 4598 7098
rect 4302 7044 4358 7046
rect 4382 7044 4438 7046
rect 4462 7044 4518 7046
rect 4542 7044 4598 7046
rect 4302 6010 4358 6012
rect 4382 6010 4438 6012
rect 4462 6010 4518 6012
rect 4542 6010 4598 6012
rect 4302 5958 4348 6010
rect 4348 5958 4358 6010
rect 4382 5958 4412 6010
rect 4412 5958 4424 6010
rect 4424 5958 4438 6010
rect 4462 5958 4476 6010
rect 4476 5958 4488 6010
rect 4488 5958 4518 6010
rect 4542 5958 4552 6010
rect 4552 5958 4598 6010
rect 4302 5956 4358 5958
rect 4382 5956 4438 5958
rect 4462 5956 4518 5958
rect 4542 5956 4598 5958
rect 4302 4922 4358 4924
rect 4382 4922 4438 4924
rect 4462 4922 4518 4924
rect 4542 4922 4598 4924
rect 4302 4870 4348 4922
rect 4348 4870 4358 4922
rect 4382 4870 4412 4922
rect 4412 4870 4424 4922
rect 4424 4870 4438 4922
rect 4462 4870 4476 4922
rect 4476 4870 4488 4922
rect 4488 4870 4518 4922
rect 4542 4870 4552 4922
rect 4552 4870 4598 4922
rect 4302 4868 4358 4870
rect 4382 4868 4438 4870
rect 4462 4868 4518 4870
rect 4542 4868 4598 4870
rect 4302 3834 4358 3836
rect 4382 3834 4438 3836
rect 4462 3834 4518 3836
rect 4542 3834 4598 3836
rect 4302 3782 4348 3834
rect 4348 3782 4358 3834
rect 4382 3782 4412 3834
rect 4412 3782 4424 3834
rect 4424 3782 4438 3834
rect 4462 3782 4476 3834
rect 4476 3782 4488 3834
rect 4488 3782 4518 3834
rect 4542 3782 4552 3834
rect 4552 3782 4598 3834
rect 4302 3780 4358 3782
rect 4382 3780 4438 3782
rect 4462 3780 4518 3782
rect 4542 3780 4598 3782
rect 7648 14170 7704 14172
rect 7728 14170 7784 14172
rect 7808 14170 7864 14172
rect 7888 14170 7944 14172
rect 7648 14118 7694 14170
rect 7694 14118 7704 14170
rect 7728 14118 7758 14170
rect 7758 14118 7770 14170
rect 7770 14118 7784 14170
rect 7808 14118 7822 14170
rect 7822 14118 7834 14170
rect 7834 14118 7864 14170
rect 7888 14118 7898 14170
rect 7898 14118 7944 14170
rect 7648 14116 7704 14118
rect 7728 14116 7784 14118
rect 7808 14116 7864 14118
rect 7888 14116 7944 14118
rect 7648 13082 7704 13084
rect 7728 13082 7784 13084
rect 7808 13082 7864 13084
rect 7888 13082 7944 13084
rect 7648 13030 7694 13082
rect 7694 13030 7704 13082
rect 7728 13030 7758 13082
rect 7758 13030 7770 13082
rect 7770 13030 7784 13082
rect 7808 13030 7822 13082
rect 7822 13030 7834 13082
rect 7834 13030 7864 13082
rect 7888 13030 7898 13082
rect 7898 13030 7944 13082
rect 7648 13028 7704 13030
rect 7728 13028 7784 13030
rect 7808 13028 7864 13030
rect 7888 13028 7944 13030
rect 7648 11994 7704 11996
rect 7728 11994 7784 11996
rect 7808 11994 7864 11996
rect 7888 11994 7944 11996
rect 7648 11942 7694 11994
rect 7694 11942 7704 11994
rect 7728 11942 7758 11994
rect 7758 11942 7770 11994
rect 7770 11942 7784 11994
rect 7808 11942 7822 11994
rect 7822 11942 7834 11994
rect 7834 11942 7864 11994
rect 7888 11942 7898 11994
rect 7898 11942 7944 11994
rect 7648 11940 7704 11942
rect 7728 11940 7784 11942
rect 7808 11940 7864 11942
rect 7888 11940 7944 11942
rect 7648 10906 7704 10908
rect 7728 10906 7784 10908
rect 7808 10906 7864 10908
rect 7888 10906 7944 10908
rect 7648 10854 7694 10906
rect 7694 10854 7704 10906
rect 7728 10854 7758 10906
rect 7758 10854 7770 10906
rect 7770 10854 7784 10906
rect 7808 10854 7822 10906
rect 7822 10854 7834 10906
rect 7834 10854 7864 10906
rect 7888 10854 7898 10906
rect 7898 10854 7944 10906
rect 7648 10852 7704 10854
rect 7728 10852 7784 10854
rect 7808 10852 7864 10854
rect 7888 10852 7944 10854
rect 7648 9818 7704 9820
rect 7728 9818 7784 9820
rect 7808 9818 7864 9820
rect 7888 9818 7944 9820
rect 7648 9766 7694 9818
rect 7694 9766 7704 9818
rect 7728 9766 7758 9818
rect 7758 9766 7770 9818
rect 7770 9766 7784 9818
rect 7808 9766 7822 9818
rect 7822 9766 7834 9818
rect 7834 9766 7864 9818
rect 7888 9766 7898 9818
rect 7898 9766 7944 9818
rect 7648 9764 7704 9766
rect 7728 9764 7784 9766
rect 7808 9764 7864 9766
rect 7888 9764 7944 9766
rect 7648 8730 7704 8732
rect 7728 8730 7784 8732
rect 7808 8730 7864 8732
rect 7888 8730 7944 8732
rect 7648 8678 7694 8730
rect 7694 8678 7704 8730
rect 7728 8678 7758 8730
rect 7758 8678 7770 8730
rect 7770 8678 7784 8730
rect 7808 8678 7822 8730
rect 7822 8678 7834 8730
rect 7834 8678 7864 8730
rect 7888 8678 7898 8730
rect 7898 8678 7944 8730
rect 7648 8676 7704 8678
rect 7728 8676 7784 8678
rect 7808 8676 7864 8678
rect 7888 8676 7944 8678
rect 7648 7642 7704 7644
rect 7728 7642 7784 7644
rect 7808 7642 7864 7644
rect 7888 7642 7944 7644
rect 7648 7590 7694 7642
rect 7694 7590 7704 7642
rect 7728 7590 7758 7642
rect 7758 7590 7770 7642
rect 7770 7590 7784 7642
rect 7808 7590 7822 7642
rect 7822 7590 7834 7642
rect 7834 7590 7864 7642
rect 7888 7590 7898 7642
rect 7898 7590 7944 7642
rect 7648 7588 7704 7590
rect 7728 7588 7784 7590
rect 7808 7588 7864 7590
rect 7888 7588 7944 7590
rect 7648 6554 7704 6556
rect 7728 6554 7784 6556
rect 7808 6554 7864 6556
rect 7888 6554 7944 6556
rect 7648 6502 7694 6554
rect 7694 6502 7704 6554
rect 7728 6502 7758 6554
rect 7758 6502 7770 6554
rect 7770 6502 7784 6554
rect 7808 6502 7822 6554
rect 7822 6502 7834 6554
rect 7834 6502 7864 6554
rect 7888 6502 7898 6554
rect 7898 6502 7944 6554
rect 7648 6500 7704 6502
rect 7728 6500 7784 6502
rect 7808 6500 7864 6502
rect 7888 6500 7944 6502
rect 7648 5466 7704 5468
rect 7728 5466 7784 5468
rect 7808 5466 7864 5468
rect 7888 5466 7944 5468
rect 7648 5414 7694 5466
rect 7694 5414 7704 5466
rect 7728 5414 7758 5466
rect 7758 5414 7770 5466
rect 7770 5414 7784 5466
rect 7808 5414 7822 5466
rect 7822 5414 7834 5466
rect 7834 5414 7864 5466
rect 7888 5414 7898 5466
rect 7898 5414 7944 5466
rect 7648 5412 7704 5414
rect 7728 5412 7784 5414
rect 7808 5412 7864 5414
rect 7888 5412 7944 5414
rect 9310 13232 9366 13288
rect 10994 23418 11050 23420
rect 11074 23418 11130 23420
rect 11154 23418 11210 23420
rect 11234 23418 11290 23420
rect 10994 23366 11040 23418
rect 11040 23366 11050 23418
rect 11074 23366 11104 23418
rect 11104 23366 11116 23418
rect 11116 23366 11130 23418
rect 11154 23366 11168 23418
rect 11168 23366 11180 23418
rect 11180 23366 11210 23418
rect 11234 23366 11244 23418
rect 11244 23366 11290 23418
rect 10994 23364 11050 23366
rect 11074 23364 11130 23366
rect 11154 23364 11210 23366
rect 11234 23364 11290 23366
rect 10994 22330 11050 22332
rect 11074 22330 11130 22332
rect 11154 22330 11210 22332
rect 11234 22330 11290 22332
rect 10994 22278 11040 22330
rect 11040 22278 11050 22330
rect 11074 22278 11104 22330
rect 11104 22278 11116 22330
rect 11116 22278 11130 22330
rect 11154 22278 11168 22330
rect 11168 22278 11180 22330
rect 11180 22278 11210 22330
rect 11234 22278 11244 22330
rect 11244 22278 11290 22330
rect 10994 22276 11050 22278
rect 11074 22276 11130 22278
rect 11154 22276 11210 22278
rect 11234 22276 11290 22278
rect 10994 21242 11050 21244
rect 11074 21242 11130 21244
rect 11154 21242 11210 21244
rect 11234 21242 11290 21244
rect 10994 21190 11040 21242
rect 11040 21190 11050 21242
rect 11074 21190 11104 21242
rect 11104 21190 11116 21242
rect 11116 21190 11130 21242
rect 11154 21190 11168 21242
rect 11168 21190 11180 21242
rect 11180 21190 11210 21242
rect 11234 21190 11244 21242
rect 11244 21190 11290 21242
rect 10994 21188 11050 21190
rect 11074 21188 11130 21190
rect 11154 21188 11210 21190
rect 11234 21188 11290 21190
rect 10994 20154 11050 20156
rect 11074 20154 11130 20156
rect 11154 20154 11210 20156
rect 11234 20154 11290 20156
rect 10994 20102 11040 20154
rect 11040 20102 11050 20154
rect 11074 20102 11104 20154
rect 11104 20102 11116 20154
rect 11116 20102 11130 20154
rect 11154 20102 11168 20154
rect 11168 20102 11180 20154
rect 11180 20102 11210 20154
rect 11234 20102 11244 20154
rect 11244 20102 11290 20154
rect 10994 20100 11050 20102
rect 11074 20100 11130 20102
rect 11154 20100 11210 20102
rect 11234 20100 11290 20102
rect 10994 19066 11050 19068
rect 11074 19066 11130 19068
rect 11154 19066 11210 19068
rect 11234 19066 11290 19068
rect 10994 19014 11040 19066
rect 11040 19014 11050 19066
rect 11074 19014 11104 19066
rect 11104 19014 11116 19066
rect 11116 19014 11130 19066
rect 11154 19014 11168 19066
rect 11168 19014 11180 19066
rect 11180 19014 11210 19066
rect 11234 19014 11244 19066
rect 11244 19014 11290 19066
rect 10994 19012 11050 19014
rect 11074 19012 11130 19014
rect 11154 19012 11210 19014
rect 11234 19012 11290 19014
rect 10994 17978 11050 17980
rect 11074 17978 11130 17980
rect 11154 17978 11210 17980
rect 11234 17978 11290 17980
rect 10994 17926 11040 17978
rect 11040 17926 11050 17978
rect 11074 17926 11104 17978
rect 11104 17926 11116 17978
rect 11116 17926 11130 17978
rect 11154 17926 11168 17978
rect 11168 17926 11180 17978
rect 11180 17926 11210 17978
rect 11234 17926 11244 17978
rect 11244 17926 11290 17978
rect 10994 17924 11050 17926
rect 11074 17924 11130 17926
rect 11154 17924 11210 17926
rect 11234 17924 11290 17926
rect 14340 26138 14396 26140
rect 14420 26138 14476 26140
rect 14500 26138 14556 26140
rect 14580 26138 14636 26140
rect 14340 26086 14386 26138
rect 14386 26086 14396 26138
rect 14420 26086 14450 26138
rect 14450 26086 14462 26138
rect 14462 26086 14476 26138
rect 14500 26086 14514 26138
rect 14514 26086 14526 26138
rect 14526 26086 14556 26138
rect 14580 26086 14590 26138
rect 14590 26086 14636 26138
rect 14340 26084 14396 26086
rect 14420 26084 14476 26086
rect 14500 26084 14556 26086
rect 14580 26084 14636 26086
rect 14340 25050 14396 25052
rect 14420 25050 14476 25052
rect 14500 25050 14556 25052
rect 14580 25050 14636 25052
rect 14340 24998 14386 25050
rect 14386 24998 14396 25050
rect 14420 24998 14450 25050
rect 14450 24998 14462 25050
rect 14462 24998 14476 25050
rect 14500 24998 14514 25050
rect 14514 24998 14526 25050
rect 14526 24998 14556 25050
rect 14580 24998 14590 25050
rect 14590 24998 14636 25050
rect 14340 24996 14396 24998
rect 14420 24996 14476 24998
rect 14500 24996 14556 24998
rect 14580 24996 14636 24998
rect 14340 23962 14396 23964
rect 14420 23962 14476 23964
rect 14500 23962 14556 23964
rect 14580 23962 14636 23964
rect 14340 23910 14386 23962
rect 14386 23910 14396 23962
rect 14420 23910 14450 23962
rect 14450 23910 14462 23962
rect 14462 23910 14476 23962
rect 14500 23910 14514 23962
rect 14514 23910 14526 23962
rect 14526 23910 14556 23962
rect 14580 23910 14590 23962
rect 14590 23910 14636 23962
rect 14340 23908 14396 23910
rect 14420 23908 14476 23910
rect 14500 23908 14556 23910
rect 14580 23908 14636 23910
rect 14340 22874 14396 22876
rect 14420 22874 14476 22876
rect 14500 22874 14556 22876
rect 14580 22874 14636 22876
rect 14340 22822 14386 22874
rect 14386 22822 14396 22874
rect 14420 22822 14450 22874
rect 14450 22822 14462 22874
rect 14462 22822 14476 22874
rect 14500 22822 14514 22874
rect 14514 22822 14526 22874
rect 14526 22822 14556 22874
rect 14580 22822 14590 22874
rect 14590 22822 14636 22874
rect 14340 22820 14396 22822
rect 14420 22820 14476 22822
rect 14500 22820 14556 22822
rect 14580 22820 14636 22822
rect 10994 16890 11050 16892
rect 11074 16890 11130 16892
rect 11154 16890 11210 16892
rect 11234 16890 11290 16892
rect 10994 16838 11040 16890
rect 11040 16838 11050 16890
rect 11074 16838 11104 16890
rect 11104 16838 11116 16890
rect 11116 16838 11130 16890
rect 11154 16838 11168 16890
rect 11168 16838 11180 16890
rect 11180 16838 11210 16890
rect 11234 16838 11244 16890
rect 11244 16838 11290 16890
rect 10994 16836 11050 16838
rect 11074 16836 11130 16838
rect 11154 16836 11210 16838
rect 11234 16836 11290 16838
rect 10994 15802 11050 15804
rect 11074 15802 11130 15804
rect 11154 15802 11210 15804
rect 11234 15802 11290 15804
rect 10994 15750 11040 15802
rect 11040 15750 11050 15802
rect 11074 15750 11104 15802
rect 11104 15750 11116 15802
rect 11116 15750 11130 15802
rect 11154 15750 11168 15802
rect 11168 15750 11180 15802
rect 11180 15750 11210 15802
rect 11234 15750 11244 15802
rect 11244 15750 11290 15802
rect 10994 15748 11050 15750
rect 11074 15748 11130 15750
rect 11154 15748 11210 15750
rect 11234 15748 11290 15750
rect 10994 14714 11050 14716
rect 11074 14714 11130 14716
rect 11154 14714 11210 14716
rect 11234 14714 11290 14716
rect 10994 14662 11040 14714
rect 11040 14662 11050 14714
rect 11074 14662 11104 14714
rect 11104 14662 11116 14714
rect 11116 14662 11130 14714
rect 11154 14662 11168 14714
rect 11168 14662 11180 14714
rect 11180 14662 11210 14714
rect 11234 14662 11244 14714
rect 11244 14662 11290 14714
rect 10994 14660 11050 14662
rect 11074 14660 11130 14662
rect 11154 14660 11210 14662
rect 11234 14660 11290 14662
rect 10994 13626 11050 13628
rect 11074 13626 11130 13628
rect 11154 13626 11210 13628
rect 11234 13626 11290 13628
rect 10994 13574 11040 13626
rect 11040 13574 11050 13626
rect 11074 13574 11104 13626
rect 11104 13574 11116 13626
rect 11116 13574 11130 13626
rect 11154 13574 11168 13626
rect 11168 13574 11180 13626
rect 11180 13574 11210 13626
rect 11234 13574 11244 13626
rect 11244 13574 11290 13626
rect 10994 13572 11050 13574
rect 11074 13572 11130 13574
rect 11154 13572 11210 13574
rect 11234 13572 11290 13574
rect 10994 12538 11050 12540
rect 11074 12538 11130 12540
rect 11154 12538 11210 12540
rect 11234 12538 11290 12540
rect 10994 12486 11040 12538
rect 11040 12486 11050 12538
rect 11074 12486 11104 12538
rect 11104 12486 11116 12538
rect 11116 12486 11130 12538
rect 11154 12486 11168 12538
rect 11168 12486 11180 12538
rect 11180 12486 11210 12538
rect 11234 12486 11244 12538
rect 11244 12486 11290 12538
rect 10994 12484 11050 12486
rect 11074 12484 11130 12486
rect 11154 12484 11210 12486
rect 11234 12484 11290 12486
rect 10994 11450 11050 11452
rect 11074 11450 11130 11452
rect 11154 11450 11210 11452
rect 11234 11450 11290 11452
rect 10994 11398 11040 11450
rect 11040 11398 11050 11450
rect 11074 11398 11104 11450
rect 11104 11398 11116 11450
rect 11116 11398 11130 11450
rect 11154 11398 11168 11450
rect 11168 11398 11180 11450
rect 11180 11398 11210 11450
rect 11234 11398 11244 11450
rect 11244 11398 11290 11450
rect 10994 11396 11050 11398
rect 11074 11396 11130 11398
rect 11154 11396 11210 11398
rect 11234 11396 11290 11398
rect 10994 10362 11050 10364
rect 11074 10362 11130 10364
rect 11154 10362 11210 10364
rect 11234 10362 11290 10364
rect 10994 10310 11040 10362
rect 11040 10310 11050 10362
rect 11074 10310 11104 10362
rect 11104 10310 11116 10362
rect 11116 10310 11130 10362
rect 11154 10310 11168 10362
rect 11168 10310 11180 10362
rect 11180 10310 11210 10362
rect 11234 10310 11244 10362
rect 11244 10310 11290 10362
rect 10994 10308 11050 10310
rect 11074 10308 11130 10310
rect 11154 10308 11210 10310
rect 11234 10308 11290 10310
rect 10994 9274 11050 9276
rect 11074 9274 11130 9276
rect 11154 9274 11210 9276
rect 11234 9274 11290 9276
rect 10994 9222 11040 9274
rect 11040 9222 11050 9274
rect 11074 9222 11104 9274
rect 11104 9222 11116 9274
rect 11116 9222 11130 9274
rect 11154 9222 11168 9274
rect 11168 9222 11180 9274
rect 11180 9222 11210 9274
rect 11234 9222 11244 9274
rect 11244 9222 11290 9274
rect 10994 9220 11050 9222
rect 11074 9220 11130 9222
rect 11154 9220 11210 9222
rect 11234 9220 11290 9222
rect 14340 21786 14396 21788
rect 14420 21786 14476 21788
rect 14500 21786 14556 21788
rect 14580 21786 14636 21788
rect 14340 21734 14386 21786
rect 14386 21734 14396 21786
rect 14420 21734 14450 21786
rect 14450 21734 14462 21786
rect 14462 21734 14476 21786
rect 14500 21734 14514 21786
rect 14514 21734 14526 21786
rect 14526 21734 14556 21786
rect 14580 21734 14590 21786
rect 14590 21734 14636 21786
rect 14340 21732 14396 21734
rect 14420 21732 14476 21734
rect 14500 21732 14556 21734
rect 14580 21732 14636 21734
rect 12438 13676 12440 13696
rect 12440 13676 12492 13696
rect 12492 13676 12494 13696
rect 11886 13132 11888 13152
rect 11888 13132 11940 13152
rect 11940 13132 11942 13152
rect 11886 13096 11942 13132
rect 12438 13640 12494 13676
rect 12438 13524 12494 13560
rect 12438 13504 12440 13524
rect 12440 13504 12492 13524
rect 12492 13504 12494 13524
rect 12070 12960 12126 13016
rect 12714 17040 12770 17096
rect 14340 20698 14396 20700
rect 14420 20698 14476 20700
rect 14500 20698 14556 20700
rect 14580 20698 14636 20700
rect 14340 20646 14386 20698
rect 14386 20646 14396 20698
rect 14420 20646 14450 20698
rect 14450 20646 14462 20698
rect 14462 20646 14476 20698
rect 14500 20646 14514 20698
rect 14514 20646 14526 20698
rect 14526 20646 14556 20698
rect 14580 20646 14590 20698
rect 14590 20646 14636 20698
rect 14340 20644 14396 20646
rect 14420 20644 14476 20646
rect 14500 20644 14556 20646
rect 14580 20644 14636 20646
rect 17686 26682 17742 26684
rect 17766 26682 17822 26684
rect 17846 26682 17902 26684
rect 17926 26682 17982 26684
rect 17686 26630 17732 26682
rect 17732 26630 17742 26682
rect 17766 26630 17796 26682
rect 17796 26630 17808 26682
rect 17808 26630 17822 26682
rect 17846 26630 17860 26682
rect 17860 26630 17872 26682
rect 17872 26630 17902 26682
rect 17926 26630 17936 26682
rect 17936 26630 17982 26682
rect 17686 26628 17742 26630
rect 17766 26628 17822 26630
rect 17846 26628 17902 26630
rect 17926 26628 17982 26630
rect 24378 26682 24434 26684
rect 24458 26682 24514 26684
rect 24538 26682 24594 26684
rect 24618 26682 24674 26684
rect 24378 26630 24424 26682
rect 24424 26630 24434 26682
rect 24458 26630 24488 26682
rect 24488 26630 24500 26682
rect 24500 26630 24514 26682
rect 24538 26630 24552 26682
rect 24552 26630 24564 26682
rect 24564 26630 24594 26682
rect 24618 26630 24628 26682
rect 24628 26630 24674 26682
rect 24378 26628 24434 26630
rect 24458 26628 24514 26630
rect 24538 26628 24594 26630
rect 24618 26628 24674 26630
rect 17686 25594 17742 25596
rect 17766 25594 17822 25596
rect 17846 25594 17902 25596
rect 17926 25594 17982 25596
rect 17686 25542 17732 25594
rect 17732 25542 17742 25594
rect 17766 25542 17796 25594
rect 17796 25542 17808 25594
rect 17808 25542 17822 25594
rect 17846 25542 17860 25594
rect 17860 25542 17872 25594
rect 17872 25542 17902 25594
rect 17926 25542 17936 25594
rect 17936 25542 17982 25594
rect 17686 25540 17742 25542
rect 17766 25540 17822 25542
rect 17846 25540 17902 25542
rect 17926 25540 17982 25542
rect 14340 19610 14396 19612
rect 14420 19610 14476 19612
rect 14500 19610 14556 19612
rect 14580 19610 14636 19612
rect 14340 19558 14386 19610
rect 14386 19558 14396 19610
rect 14420 19558 14450 19610
rect 14450 19558 14462 19610
rect 14462 19558 14476 19610
rect 14500 19558 14514 19610
rect 14514 19558 14526 19610
rect 14526 19558 14556 19610
rect 14580 19558 14590 19610
rect 14590 19558 14636 19610
rect 14340 19556 14396 19558
rect 14420 19556 14476 19558
rect 14500 19556 14556 19558
rect 14580 19556 14636 19558
rect 14340 18522 14396 18524
rect 14420 18522 14476 18524
rect 14500 18522 14556 18524
rect 14580 18522 14636 18524
rect 14340 18470 14386 18522
rect 14386 18470 14396 18522
rect 14420 18470 14450 18522
rect 14450 18470 14462 18522
rect 14462 18470 14476 18522
rect 14500 18470 14514 18522
rect 14514 18470 14526 18522
rect 14526 18470 14556 18522
rect 14580 18470 14590 18522
rect 14590 18470 14636 18522
rect 14340 18468 14396 18470
rect 14420 18468 14476 18470
rect 14500 18468 14556 18470
rect 14580 18468 14636 18470
rect 13910 17060 13966 17096
rect 13910 17040 13912 17060
rect 13912 17040 13964 17060
rect 13964 17040 13966 17060
rect 12714 13524 12770 13560
rect 12714 13504 12716 13524
rect 12716 13504 12768 13524
rect 12768 13504 12770 13524
rect 10994 8186 11050 8188
rect 11074 8186 11130 8188
rect 11154 8186 11210 8188
rect 11234 8186 11290 8188
rect 10994 8134 11040 8186
rect 11040 8134 11050 8186
rect 11074 8134 11104 8186
rect 11104 8134 11116 8186
rect 11116 8134 11130 8186
rect 11154 8134 11168 8186
rect 11168 8134 11180 8186
rect 11180 8134 11210 8186
rect 11234 8134 11244 8186
rect 11244 8134 11290 8186
rect 10994 8132 11050 8134
rect 11074 8132 11130 8134
rect 11154 8132 11210 8134
rect 11234 8132 11290 8134
rect 10994 7098 11050 7100
rect 11074 7098 11130 7100
rect 11154 7098 11210 7100
rect 11234 7098 11290 7100
rect 10994 7046 11040 7098
rect 11040 7046 11050 7098
rect 11074 7046 11104 7098
rect 11104 7046 11116 7098
rect 11116 7046 11130 7098
rect 11154 7046 11168 7098
rect 11168 7046 11180 7098
rect 11180 7046 11210 7098
rect 11234 7046 11244 7098
rect 11244 7046 11290 7098
rect 10994 7044 11050 7046
rect 11074 7044 11130 7046
rect 11154 7044 11210 7046
rect 11234 7044 11290 7046
rect 10994 6010 11050 6012
rect 11074 6010 11130 6012
rect 11154 6010 11210 6012
rect 11234 6010 11290 6012
rect 10994 5958 11040 6010
rect 11040 5958 11050 6010
rect 11074 5958 11104 6010
rect 11104 5958 11116 6010
rect 11116 5958 11130 6010
rect 11154 5958 11168 6010
rect 11168 5958 11180 6010
rect 11180 5958 11210 6010
rect 11234 5958 11244 6010
rect 11244 5958 11290 6010
rect 10994 5956 11050 5958
rect 11074 5956 11130 5958
rect 11154 5956 11210 5958
rect 11234 5956 11290 5958
rect 12898 12552 12954 12608
rect 14340 17434 14396 17436
rect 14420 17434 14476 17436
rect 14500 17434 14556 17436
rect 14580 17434 14636 17436
rect 14340 17382 14386 17434
rect 14386 17382 14396 17434
rect 14420 17382 14450 17434
rect 14450 17382 14462 17434
rect 14462 17382 14476 17434
rect 14500 17382 14514 17434
rect 14514 17382 14526 17434
rect 14526 17382 14556 17434
rect 14580 17382 14590 17434
rect 14590 17382 14636 17434
rect 14340 17380 14396 17382
rect 14420 17380 14476 17382
rect 14500 17380 14556 17382
rect 14580 17380 14636 17382
rect 14340 16346 14396 16348
rect 14420 16346 14476 16348
rect 14500 16346 14556 16348
rect 14580 16346 14636 16348
rect 14340 16294 14386 16346
rect 14386 16294 14396 16346
rect 14420 16294 14450 16346
rect 14450 16294 14462 16346
rect 14462 16294 14476 16346
rect 14500 16294 14514 16346
rect 14514 16294 14526 16346
rect 14526 16294 14556 16346
rect 14580 16294 14590 16346
rect 14590 16294 14636 16346
rect 14340 16292 14396 16294
rect 14420 16292 14476 16294
rect 14500 16292 14556 16294
rect 14580 16292 14636 16294
rect 13726 12960 13782 13016
rect 13542 12844 13598 12880
rect 13542 12824 13544 12844
rect 13544 12824 13596 12844
rect 13596 12824 13598 12844
rect 14094 13640 14150 13696
rect 14002 13096 14058 13152
rect 14738 15952 14794 16008
rect 14340 15258 14396 15260
rect 14420 15258 14476 15260
rect 14500 15258 14556 15260
rect 14580 15258 14636 15260
rect 14340 15206 14386 15258
rect 14386 15206 14396 15258
rect 14420 15206 14450 15258
rect 14450 15206 14462 15258
rect 14462 15206 14476 15258
rect 14500 15206 14514 15258
rect 14514 15206 14526 15258
rect 14526 15206 14556 15258
rect 14580 15206 14590 15258
rect 14590 15206 14636 15258
rect 14340 15204 14396 15206
rect 14420 15204 14476 15206
rect 14500 15204 14556 15206
rect 14580 15204 14636 15206
rect 14340 14170 14396 14172
rect 14420 14170 14476 14172
rect 14500 14170 14556 14172
rect 14580 14170 14636 14172
rect 14340 14118 14386 14170
rect 14386 14118 14396 14170
rect 14420 14118 14450 14170
rect 14450 14118 14462 14170
rect 14462 14118 14476 14170
rect 14500 14118 14514 14170
rect 14514 14118 14526 14170
rect 14526 14118 14556 14170
rect 14580 14118 14590 14170
rect 14590 14118 14636 14170
rect 14340 14116 14396 14118
rect 14420 14116 14476 14118
rect 14500 14116 14556 14118
rect 14580 14116 14636 14118
rect 14922 16496 14978 16552
rect 14340 13082 14396 13084
rect 14420 13082 14476 13084
rect 14500 13082 14556 13084
rect 14580 13082 14636 13084
rect 14340 13030 14386 13082
rect 14386 13030 14396 13082
rect 14420 13030 14450 13082
rect 14450 13030 14462 13082
rect 14462 13030 14476 13082
rect 14500 13030 14514 13082
rect 14514 13030 14526 13082
rect 14526 13030 14556 13082
rect 14580 13030 14590 13082
rect 14590 13030 14636 13082
rect 14340 13028 14396 13030
rect 14420 13028 14476 13030
rect 14500 13028 14556 13030
rect 14580 13028 14636 13030
rect 14554 12552 14610 12608
rect 14340 11994 14396 11996
rect 14420 11994 14476 11996
rect 14500 11994 14556 11996
rect 14580 11994 14636 11996
rect 14340 11942 14386 11994
rect 14386 11942 14396 11994
rect 14420 11942 14450 11994
rect 14450 11942 14462 11994
rect 14462 11942 14476 11994
rect 14500 11942 14514 11994
rect 14514 11942 14526 11994
rect 14526 11942 14556 11994
rect 14580 11942 14590 11994
rect 14590 11942 14636 11994
rect 14340 11940 14396 11942
rect 14420 11940 14476 11942
rect 14500 11940 14556 11942
rect 14580 11940 14636 11942
rect 17686 24506 17742 24508
rect 17766 24506 17822 24508
rect 17846 24506 17902 24508
rect 17926 24506 17982 24508
rect 17686 24454 17732 24506
rect 17732 24454 17742 24506
rect 17766 24454 17796 24506
rect 17796 24454 17808 24506
rect 17808 24454 17822 24506
rect 17846 24454 17860 24506
rect 17860 24454 17872 24506
rect 17872 24454 17902 24506
rect 17926 24454 17936 24506
rect 17936 24454 17982 24506
rect 17686 24452 17742 24454
rect 17766 24452 17822 24454
rect 17846 24452 17902 24454
rect 17926 24452 17982 24454
rect 17686 23418 17742 23420
rect 17766 23418 17822 23420
rect 17846 23418 17902 23420
rect 17926 23418 17982 23420
rect 17686 23366 17732 23418
rect 17732 23366 17742 23418
rect 17766 23366 17796 23418
rect 17796 23366 17808 23418
rect 17808 23366 17822 23418
rect 17846 23366 17860 23418
rect 17860 23366 17872 23418
rect 17872 23366 17902 23418
rect 17926 23366 17936 23418
rect 17936 23366 17982 23418
rect 17686 23364 17742 23366
rect 17766 23364 17822 23366
rect 17846 23364 17902 23366
rect 17926 23364 17982 23366
rect 17686 22330 17742 22332
rect 17766 22330 17822 22332
rect 17846 22330 17902 22332
rect 17926 22330 17982 22332
rect 17686 22278 17732 22330
rect 17732 22278 17742 22330
rect 17766 22278 17796 22330
rect 17796 22278 17808 22330
rect 17808 22278 17822 22330
rect 17846 22278 17860 22330
rect 17860 22278 17872 22330
rect 17872 22278 17902 22330
rect 17926 22278 17936 22330
rect 17936 22278 17982 22330
rect 17686 22276 17742 22278
rect 17766 22276 17822 22278
rect 17846 22276 17902 22278
rect 17926 22276 17982 22278
rect 17686 21242 17742 21244
rect 17766 21242 17822 21244
rect 17846 21242 17902 21244
rect 17926 21242 17982 21244
rect 17686 21190 17732 21242
rect 17732 21190 17742 21242
rect 17766 21190 17796 21242
rect 17796 21190 17808 21242
rect 17808 21190 17822 21242
rect 17846 21190 17860 21242
rect 17860 21190 17872 21242
rect 17872 21190 17902 21242
rect 17926 21190 17936 21242
rect 17936 21190 17982 21242
rect 17686 21188 17742 21190
rect 17766 21188 17822 21190
rect 17846 21188 17902 21190
rect 17926 21188 17982 21190
rect 17686 20154 17742 20156
rect 17766 20154 17822 20156
rect 17846 20154 17902 20156
rect 17926 20154 17982 20156
rect 17686 20102 17732 20154
rect 17732 20102 17742 20154
rect 17766 20102 17796 20154
rect 17796 20102 17808 20154
rect 17808 20102 17822 20154
rect 17846 20102 17860 20154
rect 17860 20102 17872 20154
rect 17872 20102 17902 20154
rect 17926 20102 17936 20154
rect 17936 20102 17982 20154
rect 17686 20100 17742 20102
rect 17766 20100 17822 20102
rect 17846 20100 17902 20102
rect 17926 20100 17982 20102
rect 17686 19066 17742 19068
rect 17766 19066 17822 19068
rect 17846 19066 17902 19068
rect 17926 19066 17982 19068
rect 17686 19014 17732 19066
rect 17732 19014 17742 19066
rect 17766 19014 17796 19066
rect 17796 19014 17808 19066
rect 17808 19014 17822 19066
rect 17846 19014 17860 19066
rect 17860 19014 17872 19066
rect 17872 19014 17902 19066
rect 17926 19014 17936 19066
rect 17936 19014 17982 19066
rect 17686 19012 17742 19014
rect 17766 19012 17822 19014
rect 17846 19012 17902 19014
rect 17926 19012 17982 19014
rect 17686 17978 17742 17980
rect 17766 17978 17822 17980
rect 17846 17978 17902 17980
rect 17926 17978 17982 17980
rect 17686 17926 17732 17978
rect 17732 17926 17742 17978
rect 17766 17926 17796 17978
rect 17796 17926 17808 17978
rect 17808 17926 17822 17978
rect 17846 17926 17860 17978
rect 17860 17926 17872 17978
rect 17872 17926 17902 17978
rect 17926 17926 17936 17978
rect 17936 17926 17982 17978
rect 17686 17924 17742 17926
rect 17766 17924 17822 17926
rect 17846 17924 17902 17926
rect 17926 17924 17982 17926
rect 14340 10906 14396 10908
rect 14420 10906 14476 10908
rect 14500 10906 14556 10908
rect 14580 10906 14636 10908
rect 14340 10854 14386 10906
rect 14386 10854 14396 10906
rect 14420 10854 14450 10906
rect 14450 10854 14462 10906
rect 14462 10854 14476 10906
rect 14500 10854 14514 10906
rect 14514 10854 14526 10906
rect 14526 10854 14556 10906
rect 14580 10854 14590 10906
rect 14590 10854 14636 10906
rect 14340 10852 14396 10854
rect 14420 10852 14476 10854
rect 14500 10852 14556 10854
rect 14580 10852 14636 10854
rect 14340 9818 14396 9820
rect 14420 9818 14476 9820
rect 14500 9818 14556 9820
rect 14580 9818 14636 9820
rect 14340 9766 14386 9818
rect 14386 9766 14396 9818
rect 14420 9766 14450 9818
rect 14450 9766 14462 9818
rect 14462 9766 14476 9818
rect 14500 9766 14514 9818
rect 14514 9766 14526 9818
rect 14526 9766 14556 9818
rect 14580 9766 14590 9818
rect 14590 9766 14636 9818
rect 14340 9764 14396 9766
rect 14420 9764 14476 9766
rect 14500 9764 14556 9766
rect 14580 9764 14636 9766
rect 17686 16890 17742 16892
rect 17766 16890 17822 16892
rect 17846 16890 17902 16892
rect 17926 16890 17982 16892
rect 17686 16838 17732 16890
rect 17732 16838 17742 16890
rect 17766 16838 17796 16890
rect 17796 16838 17808 16890
rect 17808 16838 17822 16890
rect 17846 16838 17860 16890
rect 17860 16838 17872 16890
rect 17872 16838 17902 16890
rect 17926 16838 17936 16890
rect 17936 16838 17982 16890
rect 17686 16836 17742 16838
rect 17766 16836 17822 16838
rect 17846 16836 17902 16838
rect 17926 16836 17982 16838
rect 17686 15802 17742 15804
rect 17766 15802 17822 15804
rect 17846 15802 17902 15804
rect 17926 15802 17982 15804
rect 17686 15750 17732 15802
rect 17732 15750 17742 15802
rect 17766 15750 17796 15802
rect 17796 15750 17808 15802
rect 17808 15750 17822 15802
rect 17846 15750 17860 15802
rect 17860 15750 17872 15802
rect 17872 15750 17902 15802
rect 17926 15750 17936 15802
rect 17936 15750 17982 15802
rect 17686 15748 17742 15750
rect 17766 15748 17822 15750
rect 17846 15748 17902 15750
rect 17926 15748 17982 15750
rect 17686 14714 17742 14716
rect 17766 14714 17822 14716
rect 17846 14714 17902 14716
rect 17926 14714 17982 14716
rect 17686 14662 17732 14714
rect 17732 14662 17742 14714
rect 17766 14662 17796 14714
rect 17796 14662 17808 14714
rect 17808 14662 17822 14714
rect 17846 14662 17860 14714
rect 17860 14662 17872 14714
rect 17872 14662 17902 14714
rect 17926 14662 17936 14714
rect 17936 14662 17982 14714
rect 17686 14660 17742 14662
rect 17766 14660 17822 14662
rect 17846 14660 17902 14662
rect 17926 14660 17982 14662
rect 17498 13252 17554 13288
rect 17498 13232 17500 13252
rect 17500 13232 17552 13252
rect 17552 13232 17554 13252
rect 14340 8730 14396 8732
rect 14420 8730 14476 8732
rect 14500 8730 14556 8732
rect 14580 8730 14636 8732
rect 14340 8678 14386 8730
rect 14386 8678 14396 8730
rect 14420 8678 14450 8730
rect 14450 8678 14462 8730
rect 14462 8678 14476 8730
rect 14500 8678 14514 8730
rect 14514 8678 14526 8730
rect 14526 8678 14556 8730
rect 14580 8678 14590 8730
rect 14590 8678 14636 8730
rect 14340 8676 14396 8678
rect 14420 8676 14476 8678
rect 14500 8676 14556 8678
rect 14580 8676 14636 8678
rect 17686 13626 17742 13628
rect 17766 13626 17822 13628
rect 17846 13626 17902 13628
rect 17926 13626 17982 13628
rect 17686 13574 17732 13626
rect 17732 13574 17742 13626
rect 17766 13574 17796 13626
rect 17796 13574 17808 13626
rect 17808 13574 17822 13626
rect 17846 13574 17860 13626
rect 17860 13574 17872 13626
rect 17872 13574 17902 13626
rect 17926 13574 17936 13626
rect 17936 13574 17982 13626
rect 17686 13572 17742 13574
rect 17766 13572 17822 13574
rect 17846 13572 17902 13574
rect 17926 13572 17982 13574
rect 21032 26138 21088 26140
rect 21112 26138 21168 26140
rect 21192 26138 21248 26140
rect 21272 26138 21328 26140
rect 21032 26086 21078 26138
rect 21078 26086 21088 26138
rect 21112 26086 21142 26138
rect 21142 26086 21154 26138
rect 21154 26086 21168 26138
rect 21192 26086 21206 26138
rect 21206 26086 21218 26138
rect 21218 26086 21248 26138
rect 21272 26086 21282 26138
rect 21282 26086 21328 26138
rect 21032 26084 21088 26086
rect 21112 26084 21168 26086
rect 21192 26084 21248 26086
rect 21272 26084 21328 26086
rect 21032 25050 21088 25052
rect 21112 25050 21168 25052
rect 21192 25050 21248 25052
rect 21272 25050 21328 25052
rect 21032 24998 21078 25050
rect 21078 24998 21088 25050
rect 21112 24998 21142 25050
rect 21142 24998 21154 25050
rect 21154 24998 21168 25050
rect 21192 24998 21206 25050
rect 21206 24998 21218 25050
rect 21218 24998 21248 25050
rect 21272 24998 21282 25050
rect 21282 24998 21328 25050
rect 21032 24996 21088 24998
rect 21112 24996 21168 24998
rect 21192 24996 21248 24998
rect 21272 24996 21328 24998
rect 21032 23962 21088 23964
rect 21112 23962 21168 23964
rect 21192 23962 21248 23964
rect 21272 23962 21328 23964
rect 21032 23910 21078 23962
rect 21078 23910 21088 23962
rect 21112 23910 21142 23962
rect 21142 23910 21154 23962
rect 21154 23910 21168 23962
rect 21192 23910 21206 23962
rect 21206 23910 21218 23962
rect 21218 23910 21248 23962
rect 21272 23910 21282 23962
rect 21282 23910 21328 23962
rect 21032 23908 21088 23910
rect 21112 23908 21168 23910
rect 21192 23908 21248 23910
rect 21272 23908 21328 23910
rect 21032 22874 21088 22876
rect 21112 22874 21168 22876
rect 21192 22874 21248 22876
rect 21272 22874 21328 22876
rect 21032 22822 21078 22874
rect 21078 22822 21088 22874
rect 21112 22822 21142 22874
rect 21142 22822 21154 22874
rect 21154 22822 21168 22874
rect 21192 22822 21206 22874
rect 21206 22822 21218 22874
rect 21218 22822 21248 22874
rect 21272 22822 21282 22874
rect 21282 22822 21328 22874
rect 21032 22820 21088 22822
rect 21112 22820 21168 22822
rect 21192 22820 21248 22822
rect 21272 22820 21328 22822
rect 21032 21786 21088 21788
rect 21112 21786 21168 21788
rect 21192 21786 21248 21788
rect 21272 21786 21328 21788
rect 21032 21734 21078 21786
rect 21078 21734 21088 21786
rect 21112 21734 21142 21786
rect 21142 21734 21154 21786
rect 21154 21734 21168 21786
rect 21192 21734 21206 21786
rect 21206 21734 21218 21786
rect 21218 21734 21248 21786
rect 21272 21734 21282 21786
rect 21282 21734 21328 21786
rect 21032 21732 21088 21734
rect 21112 21732 21168 21734
rect 21192 21732 21248 21734
rect 21272 21732 21328 21734
rect 21032 20698 21088 20700
rect 21112 20698 21168 20700
rect 21192 20698 21248 20700
rect 21272 20698 21328 20700
rect 21032 20646 21078 20698
rect 21078 20646 21088 20698
rect 21112 20646 21142 20698
rect 21142 20646 21154 20698
rect 21154 20646 21168 20698
rect 21192 20646 21206 20698
rect 21206 20646 21218 20698
rect 21218 20646 21248 20698
rect 21272 20646 21282 20698
rect 21282 20646 21328 20698
rect 21032 20644 21088 20646
rect 21112 20644 21168 20646
rect 21192 20644 21248 20646
rect 21272 20644 21328 20646
rect 24378 25594 24434 25596
rect 24458 25594 24514 25596
rect 24538 25594 24594 25596
rect 24618 25594 24674 25596
rect 24378 25542 24424 25594
rect 24424 25542 24434 25594
rect 24458 25542 24488 25594
rect 24488 25542 24500 25594
rect 24500 25542 24514 25594
rect 24538 25542 24552 25594
rect 24552 25542 24564 25594
rect 24564 25542 24594 25594
rect 24618 25542 24628 25594
rect 24628 25542 24674 25594
rect 24378 25540 24434 25542
rect 24458 25540 24514 25542
rect 24538 25540 24594 25542
rect 24618 25540 24674 25542
rect 24378 24506 24434 24508
rect 24458 24506 24514 24508
rect 24538 24506 24594 24508
rect 24618 24506 24674 24508
rect 24378 24454 24424 24506
rect 24424 24454 24434 24506
rect 24458 24454 24488 24506
rect 24488 24454 24500 24506
rect 24500 24454 24514 24506
rect 24538 24454 24552 24506
rect 24552 24454 24564 24506
rect 24564 24454 24594 24506
rect 24618 24454 24628 24506
rect 24628 24454 24674 24506
rect 24378 24452 24434 24454
rect 24458 24452 24514 24454
rect 24538 24452 24594 24454
rect 24618 24452 24674 24454
rect 24378 23418 24434 23420
rect 24458 23418 24514 23420
rect 24538 23418 24594 23420
rect 24618 23418 24674 23420
rect 24378 23366 24424 23418
rect 24424 23366 24434 23418
rect 24458 23366 24488 23418
rect 24488 23366 24500 23418
rect 24500 23366 24514 23418
rect 24538 23366 24552 23418
rect 24552 23366 24564 23418
rect 24564 23366 24594 23418
rect 24618 23366 24628 23418
rect 24628 23366 24674 23418
rect 24378 23364 24434 23366
rect 24458 23364 24514 23366
rect 24538 23364 24594 23366
rect 24618 23364 24674 23366
rect 24378 22330 24434 22332
rect 24458 22330 24514 22332
rect 24538 22330 24594 22332
rect 24618 22330 24674 22332
rect 24378 22278 24424 22330
rect 24424 22278 24434 22330
rect 24458 22278 24488 22330
rect 24488 22278 24500 22330
rect 24500 22278 24514 22330
rect 24538 22278 24552 22330
rect 24552 22278 24564 22330
rect 24564 22278 24594 22330
rect 24618 22278 24628 22330
rect 24628 22278 24674 22330
rect 24378 22276 24434 22278
rect 24458 22276 24514 22278
rect 24538 22276 24594 22278
rect 24618 22276 24674 22278
rect 27724 26138 27780 26140
rect 27804 26138 27860 26140
rect 27884 26138 27940 26140
rect 27964 26138 28020 26140
rect 27724 26086 27770 26138
rect 27770 26086 27780 26138
rect 27804 26086 27834 26138
rect 27834 26086 27846 26138
rect 27846 26086 27860 26138
rect 27884 26086 27898 26138
rect 27898 26086 27910 26138
rect 27910 26086 27940 26138
rect 27964 26086 27974 26138
rect 27974 26086 28020 26138
rect 27724 26084 27780 26086
rect 27804 26084 27860 26086
rect 27884 26084 27940 26086
rect 27964 26084 28020 26086
rect 27724 25050 27780 25052
rect 27804 25050 27860 25052
rect 27884 25050 27940 25052
rect 27964 25050 28020 25052
rect 27724 24998 27770 25050
rect 27770 24998 27780 25050
rect 27804 24998 27834 25050
rect 27834 24998 27846 25050
rect 27846 24998 27860 25050
rect 27884 24998 27898 25050
rect 27898 24998 27910 25050
rect 27910 24998 27940 25050
rect 27964 24998 27974 25050
rect 27974 24998 28020 25050
rect 27724 24996 27780 24998
rect 27804 24996 27860 24998
rect 27884 24996 27940 24998
rect 27964 24996 28020 24998
rect 27724 23962 27780 23964
rect 27804 23962 27860 23964
rect 27884 23962 27940 23964
rect 27964 23962 28020 23964
rect 27724 23910 27770 23962
rect 27770 23910 27780 23962
rect 27804 23910 27834 23962
rect 27834 23910 27846 23962
rect 27846 23910 27860 23962
rect 27884 23910 27898 23962
rect 27898 23910 27910 23962
rect 27910 23910 27940 23962
rect 27964 23910 27974 23962
rect 27974 23910 28020 23962
rect 27724 23908 27780 23910
rect 27804 23908 27860 23910
rect 27884 23908 27940 23910
rect 27964 23908 28020 23910
rect 27724 22874 27780 22876
rect 27804 22874 27860 22876
rect 27884 22874 27940 22876
rect 27964 22874 28020 22876
rect 27724 22822 27770 22874
rect 27770 22822 27780 22874
rect 27804 22822 27834 22874
rect 27834 22822 27846 22874
rect 27846 22822 27860 22874
rect 27884 22822 27898 22874
rect 27898 22822 27910 22874
rect 27910 22822 27940 22874
rect 27964 22822 27974 22874
rect 27974 22822 28020 22874
rect 27724 22820 27780 22822
rect 27804 22820 27860 22822
rect 27884 22820 27940 22822
rect 27964 22820 28020 22822
rect 27724 21786 27780 21788
rect 27804 21786 27860 21788
rect 27884 21786 27940 21788
rect 27964 21786 28020 21788
rect 27724 21734 27770 21786
rect 27770 21734 27780 21786
rect 27804 21734 27834 21786
rect 27834 21734 27846 21786
rect 27846 21734 27860 21786
rect 27884 21734 27898 21786
rect 27898 21734 27910 21786
rect 27910 21734 27940 21786
rect 27964 21734 27974 21786
rect 27974 21734 28020 21786
rect 27724 21732 27780 21734
rect 27804 21732 27860 21734
rect 27884 21732 27940 21734
rect 27964 21732 28020 21734
rect 24378 21242 24434 21244
rect 24458 21242 24514 21244
rect 24538 21242 24594 21244
rect 24618 21242 24674 21244
rect 24378 21190 24424 21242
rect 24424 21190 24434 21242
rect 24458 21190 24488 21242
rect 24488 21190 24500 21242
rect 24500 21190 24514 21242
rect 24538 21190 24552 21242
rect 24552 21190 24564 21242
rect 24564 21190 24594 21242
rect 24618 21190 24628 21242
rect 24628 21190 24674 21242
rect 24378 21188 24434 21190
rect 24458 21188 24514 21190
rect 24538 21188 24594 21190
rect 24618 21188 24674 21190
rect 27724 20698 27780 20700
rect 27804 20698 27860 20700
rect 27884 20698 27940 20700
rect 27964 20698 28020 20700
rect 27724 20646 27770 20698
rect 27770 20646 27780 20698
rect 27804 20646 27834 20698
rect 27834 20646 27846 20698
rect 27846 20646 27860 20698
rect 27884 20646 27898 20698
rect 27898 20646 27910 20698
rect 27910 20646 27940 20698
rect 27964 20646 27974 20698
rect 27974 20646 28020 20698
rect 27724 20644 27780 20646
rect 27804 20644 27860 20646
rect 27884 20644 27940 20646
rect 27964 20644 28020 20646
rect 17686 12538 17742 12540
rect 17766 12538 17822 12540
rect 17846 12538 17902 12540
rect 17926 12538 17982 12540
rect 17686 12486 17732 12538
rect 17732 12486 17742 12538
rect 17766 12486 17796 12538
rect 17796 12486 17808 12538
rect 17808 12486 17822 12538
rect 17846 12486 17860 12538
rect 17860 12486 17872 12538
rect 17872 12486 17902 12538
rect 17926 12486 17936 12538
rect 17936 12486 17982 12538
rect 17686 12484 17742 12486
rect 17766 12484 17822 12486
rect 17846 12484 17902 12486
rect 17926 12484 17982 12486
rect 17686 11450 17742 11452
rect 17766 11450 17822 11452
rect 17846 11450 17902 11452
rect 17926 11450 17982 11452
rect 17686 11398 17732 11450
rect 17732 11398 17742 11450
rect 17766 11398 17796 11450
rect 17796 11398 17808 11450
rect 17808 11398 17822 11450
rect 17846 11398 17860 11450
rect 17860 11398 17872 11450
rect 17872 11398 17902 11450
rect 17926 11398 17936 11450
rect 17936 11398 17982 11450
rect 17686 11396 17742 11398
rect 17766 11396 17822 11398
rect 17846 11396 17902 11398
rect 17926 11396 17982 11398
rect 17686 10362 17742 10364
rect 17766 10362 17822 10364
rect 17846 10362 17902 10364
rect 17926 10362 17982 10364
rect 17686 10310 17732 10362
rect 17732 10310 17742 10362
rect 17766 10310 17796 10362
rect 17796 10310 17808 10362
rect 17808 10310 17822 10362
rect 17846 10310 17860 10362
rect 17860 10310 17872 10362
rect 17872 10310 17902 10362
rect 17926 10310 17936 10362
rect 17936 10310 17982 10362
rect 17686 10308 17742 10310
rect 17766 10308 17822 10310
rect 17846 10308 17902 10310
rect 17926 10308 17982 10310
rect 17686 9274 17742 9276
rect 17766 9274 17822 9276
rect 17846 9274 17902 9276
rect 17926 9274 17982 9276
rect 17686 9222 17732 9274
rect 17732 9222 17742 9274
rect 17766 9222 17796 9274
rect 17796 9222 17808 9274
rect 17808 9222 17822 9274
rect 17846 9222 17860 9274
rect 17860 9222 17872 9274
rect 17872 9222 17902 9274
rect 17926 9222 17936 9274
rect 17936 9222 17982 9274
rect 17686 9220 17742 9222
rect 17766 9220 17822 9222
rect 17846 9220 17902 9222
rect 17926 9220 17982 9222
rect 14340 7642 14396 7644
rect 14420 7642 14476 7644
rect 14500 7642 14556 7644
rect 14580 7642 14636 7644
rect 14340 7590 14386 7642
rect 14386 7590 14396 7642
rect 14420 7590 14450 7642
rect 14450 7590 14462 7642
rect 14462 7590 14476 7642
rect 14500 7590 14514 7642
rect 14514 7590 14526 7642
rect 14526 7590 14556 7642
rect 14580 7590 14590 7642
rect 14590 7590 14636 7642
rect 14340 7588 14396 7590
rect 14420 7588 14476 7590
rect 14500 7588 14556 7590
rect 14580 7588 14636 7590
rect 14340 6554 14396 6556
rect 14420 6554 14476 6556
rect 14500 6554 14556 6556
rect 14580 6554 14636 6556
rect 14340 6502 14386 6554
rect 14386 6502 14396 6554
rect 14420 6502 14450 6554
rect 14450 6502 14462 6554
rect 14462 6502 14476 6554
rect 14500 6502 14514 6554
rect 14514 6502 14526 6554
rect 14526 6502 14556 6554
rect 14580 6502 14590 6554
rect 14590 6502 14636 6554
rect 14340 6500 14396 6502
rect 14420 6500 14476 6502
rect 14500 6500 14556 6502
rect 14580 6500 14636 6502
rect 17686 8186 17742 8188
rect 17766 8186 17822 8188
rect 17846 8186 17902 8188
rect 17926 8186 17982 8188
rect 17686 8134 17732 8186
rect 17732 8134 17742 8186
rect 17766 8134 17796 8186
rect 17796 8134 17808 8186
rect 17808 8134 17822 8186
rect 17846 8134 17860 8186
rect 17860 8134 17872 8186
rect 17872 8134 17902 8186
rect 17926 8134 17936 8186
rect 17936 8134 17982 8186
rect 17686 8132 17742 8134
rect 17766 8132 17822 8134
rect 17846 8132 17902 8134
rect 17926 8132 17982 8134
rect 21032 19610 21088 19612
rect 21112 19610 21168 19612
rect 21192 19610 21248 19612
rect 21272 19610 21328 19612
rect 21032 19558 21078 19610
rect 21078 19558 21088 19610
rect 21112 19558 21142 19610
rect 21142 19558 21154 19610
rect 21154 19558 21168 19610
rect 21192 19558 21206 19610
rect 21206 19558 21218 19610
rect 21218 19558 21248 19610
rect 21272 19558 21282 19610
rect 21282 19558 21328 19610
rect 21032 19556 21088 19558
rect 21112 19556 21168 19558
rect 21192 19556 21248 19558
rect 21272 19556 21328 19558
rect 21032 18522 21088 18524
rect 21112 18522 21168 18524
rect 21192 18522 21248 18524
rect 21272 18522 21328 18524
rect 21032 18470 21078 18522
rect 21078 18470 21088 18522
rect 21112 18470 21142 18522
rect 21142 18470 21154 18522
rect 21154 18470 21168 18522
rect 21192 18470 21206 18522
rect 21206 18470 21218 18522
rect 21218 18470 21248 18522
rect 21272 18470 21282 18522
rect 21282 18470 21328 18522
rect 21032 18468 21088 18470
rect 21112 18468 21168 18470
rect 21192 18468 21248 18470
rect 21272 18468 21328 18470
rect 20442 12844 20498 12880
rect 20442 12824 20444 12844
rect 20444 12824 20496 12844
rect 20496 12824 20498 12844
rect 17686 7098 17742 7100
rect 17766 7098 17822 7100
rect 17846 7098 17902 7100
rect 17926 7098 17982 7100
rect 17686 7046 17732 7098
rect 17732 7046 17742 7098
rect 17766 7046 17796 7098
rect 17796 7046 17808 7098
rect 17808 7046 17822 7098
rect 17846 7046 17860 7098
rect 17860 7046 17872 7098
rect 17872 7046 17902 7098
rect 17926 7046 17936 7098
rect 17936 7046 17982 7098
rect 17686 7044 17742 7046
rect 17766 7044 17822 7046
rect 17846 7044 17902 7046
rect 17926 7044 17982 7046
rect 14340 5466 14396 5468
rect 14420 5466 14476 5468
rect 14500 5466 14556 5468
rect 14580 5466 14636 5468
rect 14340 5414 14386 5466
rect 14386 5414 14396 5466
rect 14420 5414 14450 5466
rect 14450 5414 14462 5466
rect 14462 5414 14476 5466
rect 14500 5414 14514 5466
rect 14514 5414 14526 5466
rect 14526 5414 14556 5466
rect 14580 5414 14590 5466
rect 14590 5414 14636 5466
rect 14340 5412 14396 5414
rect 14420 5412 14476 5414
rect 14500 5412 14556 5414
rect 14580 5412 14636 5414
rect 17686 6010 17742 6012
rect 17766 6010 17822 6012
rect 17846 6010 17902 6012
rect 17926 6010 17982 6012
rect 17686 5958 17732 6010
rect 17732 5958 17742 6010
rect 17766 5958 17796 6010
rect 17796 5958 17808 6010
rect 17808 5958 17822 6010
rect 17846 5958 17860 6010
rect 17860 5958 17872 6010
rect 17872 5958 17902 6010
rect 17926 5958 17936 6010
rect 17936 5958 17982 6010
rect 17686 5956 17742 5958
rect 17766 5956 17822 5958
rect 17846 5956 17902 5958
rect 17926 5956 17982 5958
rect 21032 17434 21088 17436
rect 21112 17434 21168 17436
rect 21192 17434 21248 17436
rect 21272 17434 21328 17436
rect 21032 17382 21078 17434
rect 21078 17382 21088 17434
rect 21112 17382 21142 17434
rect 21142 17382 21154 17434
rect 21154 17382 21168 17434
rect 21192 17382 21206 17434
rect 21206 17382 21218 17434
rect 21218 17382 21248 17434
rect 21272 17382 21282 17434
rect 21282 17382 21328 17434
rect 21032 17380 21088 17382
rect 21112 17380 21168 17382
rect 21192 17380 21248 17382
rect 21272 17380 21328 17382
rect 21032 16346 21088 16348
rect 21112 16346 21168 16348
rect 21192 16346 21248 16348
rect 21272 16346 21328 16348
rect 21032 16294 21078 16346
rect 21078 16294 21088 16346
rect 21112 16294 21142 16346
rect 21142 16294 21154 16346
rect 21154 16294 21168 16346
rect 21192 16294 21206 16346
rect 21206 16294 21218 16346
rect 21218 16294 21248 16346
rect 21272 16294 21282 16346
rect 21282 16294 21328 16346
rect 21032 16292 21088 16294
rect 21112 16292 21168 16294
rect 21192 16292 21248 16294
rect 21272 16292 21328 16294
rect 24378 20154 24434 20156
rect 24458 20154 24514 20156
rect 24538 20154 24594 20156
rect 24618 20154 24674 20156
rect 24378 20102 24424 20154
rect 24424 20102 24434 20154
rect 24458 20102 24488 20154
rect 24488 20102 24500 20154
rect 24500 20102 24514 20154
rect 24538 20102 24552 20154
rect 24552 20102 24564 20154
rect 24564 20102 24594 20154
rect 24618 20102 24628 20154
rect 24628 20102 24674 20154
rect 24378 20100 24434 20102
rect 24458 20100 24514 20102
rect 24538 20100 24594 20102
rect 24618 20100 24674 20102
rect 24378 19066 24434 19068
rect 24458 19066 24514 19068
rect 24538 19066 24594 19068
rect 24618 19066 24674 19068
rect 24378 19014 24424 19066
rect 24424 19014 24434 19066
rect 24458 19014 24488 19066
rect 24488 19014 24500 19066
rect 24500 19014 24514 19066
rect 24538 19014 24552 19066
rect 24552 19014 24564 19066
rect 24564 19014 24594 19066
rect 24618 19014 24628 19066
rect 24628 19014 24674 19066
rect 24378 19012 24434 19014
rect 24458 19012 24514 19014
rect 24538 19012 24594 19014
rect 24618 19012 24674 19014
rect 24378 17978 24434 17980
rect 24458 17978 24514 17980
rect 24538 17978 24594 17980
rect 24618 17978 24674 17980
rect 24378 17926 24424 17978
rect 24424 17926 24434 17978
rect 24458 17926 24488 17978
rect 24488 17926 24500 17978
rect 24500 17926 24514 17978
rect 24538 17926 24552 17978
rect 24552 17926 24564 17978
rect 24564 17926 24594 17978
rect 24618 17926 24628 17978
rect 24628 17926 24674 17978
rect 24378 17924 24434 17926
rect 24458 17924 24514 17926
rect 24538 17924 24594 17926
rect 24618 17924 24674 17926
rect 21032 15258 21088 15260
rect 21112 15258 21168 15260
rect 21192 15258 21248 15260
rect 21272 15258 21328 15260
rect 21032 15206 21078 15258
rect 21078 15206 21088 15258
rect 21112 15206 21142 15258
rect 21142 15206 21154 15258
rect 21154 15206 21168 15258
rect 21192 15206 21206 15258
rect 21206 15206 21218 15258
rect 21218 15206 21248 15258
rect 21272 15206 21282 15258
rect 21282 15206 21328 15258
rect 21032 15204 21088 15206
rect 21112 15204 21168 15206
rect 21192 15204 21248 15206
rect 21272 15204 21328 15206
rect 21032 14170 21088 14172
rect 21112 14170 21168 14172
rect 21192 14170 21248 14172
rect 21272 14170 21328 14172
rect 21032 14118 21078 14170
rect 21078 14118 21088 14170
rect 21112 14118 21142 14170
rect 21142 14118 21154 14170
rect 21154 14118 21168 14170
rect 21192 14118 21206 14170
rect 21206 14118 21218 14170
rect 21218 14118 21248 14170
rect 21272 14118 21282 14170
rect 21282 14118 21328 14170
rect 21032 14116 21088 14118
rect 21112 14116 21168 14118
rect 21192 14116 21248 14118
rect 21272 14116 21328 14118
rect 21032 13082 21088 13084
rect 21112 13082 21168 13084
rect 21192 13082 21248 13084
rect 21272 13082 21328 13084
rect 21032 13030 21078 13082
rect 21078 13030 21088 13082
rect 21112 13030 21142 13082
rect 21142 13030 21154 13082
rect 21154 13030 21168 13082
rect 21192 13030 21206 13082
rect 21206 13030 21218 13082
rect 21218 13030 21248 13082
rect 21272 13030 21282 13082
rect 21282 13030 21328 13082
rect 21032 13028 21088 13030
rect 21112 13028 21168 13030
rect 21192 13028 21248 13030
rect 21272 13028 21328 13030
rect 21032 11994 21088 11996
rect 21112 11994 21168 11996
rect 21192 11994 21248 11996
rect 21272 11994 21328 11996
rect 21032 11942 21078 11994
rect 21078 11942 21088 11994
rect 21112 11942 21142 11994
rect 21142 11942 21154 11994
rect 21154 11942 21168 11994
rect 21192 11942 21206 11994
rect 21206 11942 21218 11994
rect 21218 11942 21248 11994
rect 21272 11942 21282 11994
rect 21282 11942 21328 11994
rect 21032 11940 21088 11942
rect 21112 11940 21168 11942
rect 21192 11940 21248 11942
rect 21272 11940 21328 11942
rect 21032 10906 21088 10908
rect 21112 10906 21168 10908
rect 21192 10906 21248 10908
rect 21272 10906 21328 10908
rect 21032 10854 21078 10906
rect 21078 10854 21088 10906
rect 21112 10854 21142 10906
rect 21142 10854 21154 10906
rect 21154 10854 21168 10906
rect 21192 10854 21206 10906
rect 21206 10854 21218 10906
rect 21218 10854 21248 10906
rect 21272 10854 21282 10906
rect 21282 10854 21328 10906
rect 21032 10852 21088 10854
rect 21112 10852 21168 10854
rect 21192 10852 21248 10854
rect 21272 10852 21328 10854
rect 24378 16890 24434 16892
rect 24458 16890 24514 16892
rect 24538 16890 24594 16892
rect 24618 16890 24674 16892
rect 24378 16838 24424 16890
rect 24424 16838 24434 16890
rect 24458 16838 24488 16890
rect 24488 16838 24500 16890
rect 24500 16838 24514 16890
rect 24538 16838 24552 16890
rect 24552 16838 24564 16890
rect 24564 16838 24594 16890
rect 24618 16838 24628 16890
rect 24628 16838 24674 16890
rect 24378 16836 24434 16838
rect 24458 16836 24514 16838
rect 24538 16836 24594 16838
rect 24618 16836 24674 16838
rect 24378 15802 24434 15804
rect 24458 15802 24514 15804
rect 24538 15802 24594 15804
rect 24618 15802 24674 15804
rect 24378 15750 24424 15802
rect 24424 15750 24434 15802
rect 24458 15750 24488 15802
rect 24488 15750 24500 15802
rect 24500 15750 24514 15802
rect 24538 15750 24552 15802
rect 24552 15750 24564 15802
rect 24564 15750 24594 15802
rect 24618 15750 24628 15802
rect 24628 15750 24674 15802
rect 24378 15748 24434 15750
rect 24458 15748 24514 15750
rect 24538 15748 24594 15750
rect 24618 15748 24674 15750
rect 27724 19610 27780 19612
rect 27804 19610 27860 19612
rect 27884 19610 27940 19612
rect 27964 19610 28020 19612
rect 27724 19558 27770 19610
rect 27770 19558 27780 19610
rect 27804 19558 27834 19610
rect 27834 19558 27846 19610
rect 27846 19558 27860 19610
rect 27884 19558 27898 19610
rect 27898 19558 27910 19610
rect 27910 19558 27940 19610
rect 27964 19558 27974 19610
rect 27974 19558 28020 19610
rect 27724 19556 27780 19558
rect 27804 19556 27860 19558
rect 27884 19556 27940 19558
rect 27964 19556 28020 19558
rect 27724 18522 27780 18524
rect 27804 18522 27860 18524
rect 27884 18522 27940 18524
rect 27964 18522 28020 18524
rect 27724 18470 27770 18522
rect 27770 18470 27780 18522
rect 27804 18470 27834 18522
rect 27834 18470 27846 18522
rect 27846 18470 27860 18522
rect 27884 18470 27898 18522
rect 27898 18470 27910 18522
rect 27910 18470 27940 18522
rect 27964 18470 27974 18522
rect 27974 18470 28020 18522
rect 27724 18468 27780 18470
rect 27804 18468 27860 18470
rect 27884 18468 27940 18470
rect 27964 18468 28020 18470
rect 27724 17434 27780 17436
rect 27804 17434 27860 17436
rect 27884 17434 27940 17436
rect 27964 17434 28020 17436
rect 27724 17382 27770 17434
rect 27770 17382 27780 17434
rect 27804 17382 27834 17434
rect 27834 17382 27846 17434
rect 27846 17382 27860 17434
rect 27884 17382 27898 17434
rect 27898 17382 27910 17434
rect 27910 17382 27940 17434
rect 27964 17382 27974 17434
rect 27974 17382 28020 17434
rect 27724 17380 27780 17382
rect 27804 17380 27860 17382
rect 27884 17380 27940 17382
rect 27964 17380 28020 17382
rect 27724 16346 27780 16348
rect 27804 16346 27860 16348
rect 27884 16346 27940 16348
rect 27964 16346 28020 16348
rect 27724 16294 27770 16346
rect 27770 16294 27780 16346
rect 27804 16294 27834 16346
rect 27834 16294 27846 16346
rect 27846 16294 27860 16346
rect 27884 16294 27898 16346
rect 27898 16294 27910 16346
rect 27910 16294 27940 16346
rect 27964 16294 27974 16346
rect 27974 16294 28020 16346
rect 27724 16292 27780 16294
rect 27804 16292 27860 16294
rect 27884 16292 27940 16294
rect 27964 16292 28020 16294
rect 27724 15258 27780 15260
rect 27804 15258 27860 15260
rect 27884 15258 27940 15260
rect 27964 15258 28020 15260
rect 27724 15206 27770 15258
rect 27770 15206 27780 15258
rect 27804 15206 27834 15258
rect 27834 15206 27846 15258
rect 27846 15206 27860 15258
rect 27884 15206 27898 15258
rect 27898 15206 27910 15258
rect 27910 15206 27940 15258
rect 27964 15206 27974 15258
rect 27974 15206 28020 15258
rect 27724 15204 27780 15206
rect 27804 15204 27860 15206
rect 27884 15204 27940 15206
rect 27964 15204 28020 15206
rect 24378 14714 24434 14716
rect 24458 14714 24514 14716
rect 24538 14714 24594 14716
rect 24618 14714 24674 14716
rect 24378 14662 24424 14714
rect 24424 14662 24434 14714
rect 24458 14662 24488 14714
rect 24488 14662 24500 14714
rect 24500 14662 24514 14714
rect 24538 14662 24552 14714
rect 24552 14662 24564 14714
rect 24564 14662 24594 14714
rect 24618 14662 24628 14714
rect 24628 14662 24674 14714
rect 24378 14660 24434 14662
rect 24458 14660 24514 14662
rect 24538 14660 24594 14662
rect 24618 14660 24674 14662
rect 24378 13626 24434 13628
rect 24458 13626 24514 13628
rect 24538 13626 24594 13628
rect 24618 13626 24674 13628
rect 24378 13574 24424 13626
rect 24424 13574 24434 13626
rect 24458 13574 24488 13626
rect 24488 13574 24500 13626
rect 24500 13574 24514 13626
rect 24538 13574 24552 13626
rect 24552 13574 24564 13626
rect 24564 13574 24594 13626
rect 24618 13574 24628 13626
rect 24628 13574 24674 13626
rect 24378 13572 24434 13574
rect 24458 13572 24514 13574
rect 24538 13572 24594 13574
rect 24618 13572 24674 13574
rect 21032 9818 21088 9820
rect 21112 9818 21168 9820
rect 21192 9818 21248 9820
rect 21272 9818 21328 9820
rect 21032 9766 21078 9818
rect 21078 9766 21088 9818
rect 21112 9766 21142 9818
rect 21142 9766 21154 9818
rect 21154 9766 21168 9818
rect 21192 9766 21206 9818
rect 21206 9766 21218 9818
rect 21218 9766 21248 9818
rect 21272 9766 21282 9818
rect 21282 9766 21328 9818
rect 21032 9764 21088 9766
rect 21112 9764 21168 9766
rect 21192 9764 21248 9766
rect 21272 9764 21328 9766
rect 21032 8730 21088 8732
rect 21112 8730 21168 8732
rect 21192 8730 21248 8732
rect 21272 8730 21328 8732
rect 21032 8678 21078 8730
rect 21078 8678 21088 8730
rect 21112 8678 21142 8730
rect 21142 8678 21154 8730
rect 21154 8678 21168 8730
rect 21192 8678 21206 8730
rect 21206 8678 21218 8730
rect 21218 8678 21248 8730
rect 21272 8678 21282 8730
rect 21282 8678 21328 8730
rect 21032 8676 21088 8678
rect 21112 8676 21168 8678
rect 21192 8676 21248 8678
rect 21272 8676 21328 8678
rect 10994 4922 11050 4924
rect 11074 4922 11130 4924
rect 11154 4922 11210 4924
rect 11234 4922 11290 4924
rect 10994 4870 11040 4922
rect 11040 4870 11050 4922
rect 11074 4870 11104 4922
rect 11104 4870 11116 4922
rect 11116 4870 11130 4922
rect 11154 4870 11168 4922
rect 11168 4870 11180 4922
rect 11180 4870 11210 4922
rect 11234 4870 11244 4922
rect 11244 4870 11290 4922
rect 10994 4868 11050 4870
rect 11074 4868 11130 4870
rect 11154 4868 11210 4870
rect 11234 4868 11290 4870
rect 17686 4922 17742 4924
rect 17766 4922 17822 4924
rect 17846 4922 17902 4924
rect 17926 4922 17982 4924
rect 17686 4870 17732 4922
rect 17732 4870 17742 4922
rect 17766 4870 17796 4922
rect 17796 4870 17808 4922
rect 17808 4870 17822 4922
rect 17846 4870 17860 4922
rect 17860 4870 17872 4922
rect 17872 4870 17902 4922
rect 17926 4870 17936 4922
rect 17936 4870 17982 4922
rect 17686 4868 17742 4870
rect 17766 4868 17822 4870
rect 17846 4868 17902 4870
rect 17926 4868 17982 4870
rect 7648 4378 7704 4380
rect 7728 4378 7784 4380
rect 7808 4378 7864 4380
rect 7888 4378 7944 4380
rect 7648 4326 7694 4378
rect 7694 4326 7704 4378
rect 7728 4326 7758 4378
rect 7758 4326 7770 4378
rect 7770 4326 7784 4378
rect 7808 4326 7822 4378
rect 7822 4326 7834 4378
rect 7834 4326 7864 4378
rect 7888 4326 7898 4378
rect 7898 4326 7944 4378
rect 7648 4324 7704 4326
rect 7728 4324 7784 4326
rect 7808 4324 7864 4326
rect 7888 4324 7944 4326
rect 14340 4378 14396 4380
rect 14420 4378 14476 4380
rect 14500 4378 14556 4380
rect 14580 4378 14636 4380
rect 14340 4326 14386 4378
rect 14386 4326 14396 4378
rect 14420 4326 14450 4378
rect 14450 4326 14462 4378
rect 14462 4326 14476 4378
rect 14500 4326 14514 4378
rect 14514 4326 14526 4378
rect 14526 4326 14556 4378
rect 14580 4326 14590 4378
rect 14590 4326 14636 4378
rect 14340 4324 14396 4326
rect 14420 4324 14476 4326
rect 14500 4324 14556 4326
rect 14580 4324 14636 4326
rect 21032 7642 21088 7644
rect 21112 7642 21168 7644
rect 21192 7642 21248 7644
rect 21272 7642 21328 7644
rect 21032 7590 21078 7642
rect 21078 7590 21088 7642
rect 21112 7590 21142 7642
rect 21142 7590 21154 7642
rect 21154 7590 21168 7642
rect 21192 7590 21206 7642
rect 21206 7590 21218 7642
rect 21218 7590 21248 7642
rect 21272 7590 21282 7642
rect 21282 7590 21328 7642
rect 21032 7588 21088 7590
rect 21112 7588 21168 7590
rect 21192 7588 21248 7590
rect 21272 7588 21328 7590
rect 24378 12538 24434 12540
rect 24458 12538 24514 12540
rect 24538 12538 24594 12540
rect 24618 12538 24674 12540
rect 24378 12486 24424 12538
rect 24424 12486 24434 12538
rect 24458 12486 24488 12538
rect 24488 12486 24500 12538
rect 24500 12486 24514 12538
rect 24538 12486 24552 12538
rect 24552 12486 24564 12538
rect 24564 12486 24594 12538
rect 24618 12486 24628 12538
rect 24628 12486 24674 12538
rect 24378 12484 24434 12486
rect 24458 12484 24514 12486
rect 24538 12484 24594 12486
rect 24618 12484 24674 12486
rect 24378 11450 24434 11452
rect 24458 11450 24514 11452
rect 24538 11450 24594 11452
rect 24618 11450 24674 11452
rect 24378 11398 24424 11450
rect 24424 11398 24434 11450
rect 24458 11398 24488 11450
rect 24488 11398 24500 11450
rect 24500 11398 24514 11450
rect 24538 11398 24552 11450
rect 24552 11398 24564 11450
rect 24564 11398 24594 11450
rect 24618 11398 24628 11450
rect 24628 11398 24674 11450
rect 24378 11396 24434 11398
rect 24458 11396 24514 11398
rect 24538 11396 24594 11398
rect 24618 11396 24674 11398
rect 24378 10362 24434 10364
rect 24458 10362 24514 10364
rect 24538 10362 24594 10364
rect 24618 10362 24674 10364
rect 24378 10310 24424 10362
rect 24424 10310 24434 10362
rect 24458 10310 24488 10362
rect 24488 10310 24500 10362
rect 24500 10310 24514 10362
rect 24538 10310 24552 10362
rect 24552 10310 24564 10362
rect 24564 10310 24594 10362
rect 24618 10310 24628 10362
rect 24628 10310 24674 10362
rect 24378 10308 24434 10310
rect 24458 10308 24514 10310
rect 24538 10308 24594 10310
rect 24618 10308 24674 10310
rect 27724 14170 27780 14172
rect 27804 14170 27860 14172
rect 27884 14170 27940 14172
rect 27964 14170 28020 14172
rect 27724 14118 27770 14170
rect 27770 14118 27780 14170
rect 27804 14118 27834 14170
rect 27834 14118 27846 14170
rect 27846 14118 27860 14170
rect 27884 14118 27898 14170
rect 27898 14118 27910 14170
rect 27910 14118 27940 14170
rect 27964 14118 27974 14170
rect 27974 14118 28020 14170
rect 27724 14116 27780 14118
rect 27804 14116 27860 14118
rect 27884 14116 27940 14118
rect 27964 14116 28020 14118
rect 27724 13082 27780 13084
rect 27804 13082 27860 13084
rect 27884 13082 27940 13084
rect 27964 13082 28020 13084
rect 27724 13030 27770 13082
rect 27770 13030 27780 13082
rect 27804 13030 27834 13082
rect 27834 13030 27846 13082
rect 27846 13030 27860 13082
rect 27884 13030 27898 13082
rect 27898 13030 27910 13082
rect 27910 13030 27940 13082
rect 27964 13030 27974 13082
rect 27974 13030 28020 13082
rect 27724 13028 27780 13030
rect 27804 13028 27860 13030
rect 27884 13028 27940 13030
rect 27964 13028 28020 13030
rect 27724 11994 27780 11996
rect 27804 11994 27860 11996
rect 27884 11994 27940 11996
rect 27964 11994 28020 11996
rect 27724 11942 27770 11994
rect 27770 11942 27780 11994
rect 27804 11942 27834 11994
rect 27834 11942 27846 11994
rect 27846 11942 27860 11994
rect 27884 11942 27898 11994
rect 27898 11942 27910 11994
rect 27910 11942 27940 11994
rect 27964 11942 27974 11994
rect 27974 11942 28020 11994
rect 27724 11940 27780 11942
rect 27804 11940 27860 11942
rect 27884 11940 27940 11942
rect 27964 11940 28020 11942
rect 27724 10906 27780 10908
rect 27804 10906 27860 10908
rect 27884 10906 27940 10908
rect 27964 10906 28020 10908
rect 27724 10854 27770 10906
rect 27770 10854 27780 10906
rect 27804 10854 27834 10906
rect 27834 10854 27846 10906
rect 27846 10854 27860 10906
rect 27884 10854 27898 10906
rect 27898 10854 27910 10906
rect 27910 10854 27940 10906
rect 27964 10854 27974 10906
rect 27974 10854 28020 10906
rect 27724 10852 27780 10854
rect 27804 10852 27860 10854
rect 27884 10852 27940 10854
rect 27964 10852 28020 10854
rect 24378 9274 24434 9276
rect 24458 9274 24514 9276
rect 24538 9274 24594 9276
rect 24618 9274 24674 9276
rect 24378 9222 24424 9274
rect 24424 9222 24434 9274
rect 24458 9222 24488 9274
rect 24488 9222 24500 9274
rect 24500 9222 24514 9274
rect 24538 9222 24552 9274
rect 24552 9222 24564 9274
rect 24564 9222 24594 9274
rect 24618 9222 24628 9274
rect 24628 9222 24674 9274
rect 24378 9220 24434 9222
rect 24458 9220 24514 9222
rect 24538 9220 24594 9222
rect 24618 9220 24674 9222
rect 27724 9818 27780 9820
rect 27804 9818 27860 9820
rect 27884 9818 27940 9820
rect 27964 9818 28020 9820
rect 27724 9766 27770 9818
rect 27770 9766 27780 9818
rect 27804 9766 27834 9818
rect 27834 9766 27846 9818
rect 27846 9766 27860 9818
rect 27884 9766 27898 9818
rect 27898 9766 27910 9818
rect 27910 9766 27940 9818
rect 27964 9766 27974 9818
rect 27974 9766 28020 9818
rect 27724 9764 27780 9766
rect 27804 9764 27860 9766
rect 27884 9764 27940 9766
rect 27964 9764 28020 9766
rect 24378 8186 24434 8188
rect 24458 8186 24514 8188
rect 24538 8186 24594 8188
rect 24618 8186 24674 8188
rect 24378 8134 24424 8186
rect 24424 8134 24434 8186
rect 24458 8134 24488 8186
rect 24488 8134 24500 8186
rect 24500 8134 24514 8186
rect 24538 8134 24552 8186
rect 24552 8134 24564 8186
rect 24564 8134 24594 8186
rect 24618 8134 24628 8186
rect 24628 8134 24674 8186
rect 24378 8132 24434 8134
rect 24458 8132 24514 8134
rect 24538 8132 24594 8134
rect 24618 8132 24674 8134
rect 27724 8730 27780 8732
rect 27804 8730 27860 8732
rect 27884 8730 27940 8732
rect 27964 8730 28020 8732
rect 27724 8678 27770 8730
rect 27770 8678 27780 8730
rect 27804 8678 27834 8730
rect 27834 8678 27846 8730
rect 27846 8678 27860 8730
rect 27884 8678 27898 8730
rect 27898 8678 27910 8730
rect 27910 8678 27940 8730
rect 27964 8678 27974 8730
rect 27974 8678 28020 8730
rect 27724 8676 27780 8678
rect 27804 8676 27860 8678
rect 27884 8676 27940 8678
rect 27964 8676 28020 8678
rect 21032 6554 21088 6556
rect 21112 6554 21168 6556
rect 21192 6554 21248 6556
rect 21272 6554 21328 6556
rect 21032 6502 21078 6554
rect 21078 6502 21088 6554
rect 21112 6502 21142 6554
rect 21142 6502 21154 6554
rect 21154 6502 21168 6554
rect 21192 6502 21206 6554
rect 21206 6502 21218 6554
rect 21218 6502 21248 6554
rect 21272 6502 21282 6554
rect 21282 6502 21328 6554
rect 21032 6500 21088 6502
rect 21112 6500 21168 6502
rect 21192 6500 21248 6502
rect 21272 6500 21328 6502
rect 24378 7098 24434 7100
rect 24458 7098 24514 7100
rect 24538 7098 24594 7100
rect 24618 7098 24674 7100
rect 24378 7046 24424 7098
rect 24424 7046 24434 7098
rect 24458 7046 24488 7098
rect 24488 7046 24500 7098
rect 24500 7046 24514 7098
rect 24538 7046 24552 7098
rect 24552 7046 24564 7098
rect 24564 7046 24594 7098
rect 24618 7046 24628 7098
rect 24628 7046 24674 7098
rect 24378 7044 24434 7046
rect 24458 7044 24514 7046
rect 24538 7044 24594 7046
rect 24618 7044 24674 7046
rect 27724 7642 27780 7644
rect 27804 7642 27860 7644
rect 27884 7642 27940 7644
rect 27964 7642 28020 7644
rect 27724 7590 27770 7642
rect 27770 7590 27780 7642
rect 27804 7590 27834 7642
rect 27834 7590 27846 7642
rect 27846 7590 27860 7642
rect 27884 7590 27898 7642
rect 27898 7590 27910 7642
rect 27910 7590 27940 7642
rect 27964 7590 27974 7642
rect 27974 7590 28020 7642
rect 27724 7588 27780 7590
rect 27804 7588 27860 7590
rect 27884 7588 27940 7590
rect 27964 7588 28020 7590
rect 27724 6554 27780 6556
rect 27804 6554 27860 6556
rect 27884 6554 27940 6556
rect 27964 6554 28020 6556
rect 27724 6502 27770 6554
rect 27770 6502 27780 6554
rect 27804 6502 27834 6554
rect 27834 6502 27846 6554
rect 27846 6502 27860 6554
rect 27884 6502 27898 6554
rect 27898 6502 27910 6554
rect 27910 6502 27940 6554
rect 27964 6502 27974 6554
rect 27974 6502 28020 6554
rect 27724 6500 27780 6502
rect 27804 6500 27860 6502
rect 27884 6500 27940 6502
rect 27964 6500 28020 6502
rect 24378 6010 24434 6012
rect 24458 6010 24514 6012
rect 24538 6010 24594 6012
rect 24618 6010 24674 6012
rect 24378 5958 24424 6010
rect 24424 5958 24434 6010
rect 24458 5958 24488 6010
rect 24488 5958 24500 6010
rect 24500 5958 24514 6010
rect 24538 5958 24552 6010
rect 24552 5958 24564 6010
rect 24564 5958 24594 6010
rect 24618 5958 24628 6010
rect 24628 5958 24674 6010
rect 24378 5956 24434 5958
rect 24458 5956 24514 5958
rect 24538 5956 24594 5958
rect 24618 5956 24674 5958
rect 21032 5466 21088 5468
rect 21112 5466 21168 5468
rect 21192 5466 21248 5468
rect 21272 5466 21328 5468
rect 21032 5414 21078 5466
rect 21078 5414 21088 5466
rect 21112 5414 21142 5466
rect 21142 5414 21154 5466
rect 21154 5414 21168 5466
rect 21192 5414 21206 5466
rect 21206 5414 21218 5466
rect 21218 5414 21248 5466
rect 21272 5414 21282 5466
rect 21282 5414 21328 5466
rect 21032 5412 21088 5414
rect 21112 5412 21168 5414
rect 21192 5412 21248 5414
rect 21272 5412 21328 5414
rect 27724 5466 27780 5468
rect 27804 5466 27860 5468
rect 27884 5466 27940 5468
rect 27964 5466 28020 5468
rect 27724 5414 27770 5466
rect 27770 5414 27780 5466
rect 27804 5414 27834 5466
rect 27834 5414 27846 5466
rect 27846 5414 27860 5466
rect 27884 5414 27898 5466
rect 27898 5414 27910 5466
rect 27910 5414 27940 5466
rect 27964 5414 27974 5466
rect 27974 5414 28020 5466
rect 27724 5412 27780 5414
rect 27804 5412 27860 5414
rect 27884 5412 27940 5414
rect 27964 5412 28020 5414
rect 24378 4922 24434 4924
rect 24458 4922 24514 4924
rect 24538 4922 24594 4924
rect 24618 4922 24674 4924
rect 24378 4870 24424 4922
rect 24424 4870 24434 4922
rect 24458 4870 24488 4922
rect 24488 4870 24500 4922
rect 24500 4870 24514 4922
rect 24538 4870 24552 4922
rect 24552 4870 24564 4922
rect 24564 4870 24594 4922
rect 24618 4870 24628 4922
rect 24628 4870 24674 4922
rect 24378 4868 24434 4870
rect 24458 4868 24514 4870
rect 24538 4868 24594 4870
rect 24618 4868 24674 4870
rect 21032 4378 21088 4380
rect 21112 4378 21168 4380
rect 21192 4378 21248 4380
rect 21272 4378 21328 4380
rect 21032 4326 21078 4378
rect 21078 4326 21088 4378
rect 21112 4326 21142 4378
rect 21142 4326 21154 4378
rect 21154 4326 21168 4378
rect 21192 4326 21206 4378
rect 21206 4326 21218 4378
rect 21218 4326 21248 4378
rect 21272 4326 21282 4378
rect 21282 4326 21328 4378
rect 21032 4324 21088 4326
rect 21112 4324 21168 4326
rect 21192 4324 21248 4326
rect 21272 4324 21328 4326
rect 27724 4378 27780 4380
rect 27804 4378 27860 4380
rect 27884 4378 27940 4380
rect 27964 4378 28020 4380
rect 27724 4326 27770 4378
rect 27770 4326 27780 4378
rect 27804 4326 27834 4378
rect 27834 4326 27846 4378
rect 27846 4326 27860 4378
rect 27884 4326 27898 4378
rect 27898 4326 27910 4378
rect 27910 4326 27940 4378
rect 27964 4326 27974 4378
rect 27974 4326 28020 4378
rect 27724 4324 27780 4326
rect 27804 4324 27860 4326
rect 27884 4324 27940 4326
rect 27964 4324 28020 4326
rect 7648 3290 7704 3292
rect 7728 3290 7784 3292
rect 7808 3290 7864 3292
rect 7888 3290 7944 3292
rect 7648 3238 7694 3290
rect 7694 3238 7704 3290
rect 7728 3238 7758 3290
rect 7758 3238 7770 3290
rect 7770 3238 7784 3290
rect 7808 3238 7822 3290
rect 7822 3238 7834 3290
rect 7834 3238 7864 3290
rect 7888 3238 7898 3290
rect 7898 3238 7944 3290
rect 7648 3236 7704 3238
rect 7728 3236 7784 3238
rect 7808 3236 7864 3238
rect 7888 3236 7944 3238
rect 4302 2746 4358 2748
rect 4382 2746 4438 2748
rect 4462 2746 4518 2748
rect 4542 2746 4598 2748
rect 4302 2694 4348 2746
rect 4348 2694 4358 2746
rect 4382 2694 4412 2746
rect 4412 2694 4424 2746
rect 4424 2694 4438 2746
rect 4462 2694 4476 2746
rect 4476 2694 4488 2746
rect 4488 2694 4518 2746
rect 4542 2694 4552 2746
rect 4552 2694 4598 2746
rect 4302 2692 4358 2694
rect 4382 2692 4438 2694
rect 4462 2692 4518 2694
rect 4542 2692 4598 2694
rect 10994 3834 11050 3836
rect 11074 3834 11130 3836
rect 11154 3834 11210 3836
rect 11234 3834 11290 3836
rect 10994 3782 11040 3834
rect 11040 3782 11050 3834
rect 11074 3782 11104 3834
rect 11104 3782 11116 3834
rect 11116 3782 11130 3834
rect 11154 3782 11168 3834
rect 11168 3782 11180 3834
rect 11180 3782 11210 3834
rect 11234 3782 11244 3834
rect 11244 3782 11290 3834
rect 10994 3780 11050 3782
rect 11074 3780 11130 3782
rect 11154 3780 11210 3782
rect 11234 3780 11290 3782
rect 17686 3834 17742 3836
rect 17766 3834 17822 3836
rect 17846 3834 17902 3836
rect 17926 3834 17982 3836
rect 17686 3782 17732 3834
rect 17732 3782 17742 3834
rect 17766 3782 17796 3834
rect 17796 3782 17808 3834
rect 17808 3782 17822 3834
rect 17846 3782 17860 3834
rect 17860 3782 17872 3834
rect 17872 3782 17902 3834
rect 17926 3782 17936 3834
rect 17936 3782 17982 3834
rect 17686 3780 17742 3782
rect 17766 3780 17822 3782
rect 17846 3780 17902 3782
rect 17926 3780 17982 3782
rect 24378 3834 24434 3836
rect 24458 3834 24514 3836
rect 24538 3834 24594 3836
rect 24618 3834 24674 3836
rect 24378 3782 24424 3834
rect 24424 3782 24434 3834
rect 24458 3782 24488 3834
rect 24488 3782 24500 3834
rect 24500 3782 24514 3834
rect 24538 3782 24552 3834
rect 24552 3782 24564 3834
rect 24564 3782 24594 3834
rect 24618 3782 24628 3834
rect 24628 3782 24674 3834
rect 24378 3780 24434 3782
rect 24458 3780 24514 3782
rect 24538 3780 24594 3782
rect 24618 3780 24674 3782
rect 14340 3290 14396 3292
rect 14420 3290 14476 3292
rect 14500 3290 14556 3292
rect 14580 3290 14636 3292
rect 14340 3238 14386 3290
rect 14386 3238 14396 3290
rect 14420 3238 14450 3290
rect 14450 3238 14462 3290
rect 14462 3238 14476 3290
rect 14500 3238 14514 3290
rect 14514 3238 14526 3290
rect 14526 3238 14556 3290
rect 14580 3238 14590 3290
rect 14590 3238 14636 3290
rect 14340 3236 14396 3238
rect 14420 3236 14476 3238
rect 14500 3236 14556 3238
rect 14580 3236 14636 3238
rect 21032 3290 21088 3292
rect 21112 3290 21168 3292
rect 21192 3290 21248 3292
rect 21272 3290 21328 3292
rect 21032 3238 21078 3290
rect 21078 3238 21088 3290
rect 21112 3238 21142 3290
rect 21142 3238 21154 3290
rect 21154 3238 21168 3290
rect 21192 3238 21206 3290
rect 21206 3238 21218 3290
rect 21218 3238 21248 3290
rect 21272 3238 21282 3290
rect 21282 3238 21328 3290
rect 21032 3236 21088 3238
rect 21112 3236 21168 3238
rect 21192 3236 21248 3238
rect 21272 3236 21328 3238
rect 27724 3290 27780 3292
rect 27804 3290 27860 3292
rect 27884 3290 27940 3292
rect 27964 3290 28020 3292
rect 27724 3238 27770 3290
rect 27770 3238 27780 3290
rect 27804 3238 27834 3290
rect 27834 3238 27846 3290
rect 27846 3238 27860 3290
rect 27884 3238 27898 3290
rect 27898 3238 27910 3290
rect 27910 3238 27940 3290
rect 27964 3238 27974 3290
rect 27974 3238 28020 3290
rect 27724 3236 27780 3238
rect 27804 3236 27860 3238
rect 27884 3236 27940 3238
rect 27964 3236 28020 3238
rect 10994 2746 11050 2748
rect 11074 2746 11130 2748
rect 11154 2746 11210 2748
rect 11234 2746 11290 2748
rect 10994 2694 11040 2746
rect 11040 2694 11050 2746
rect 11074 2694 11104 2746
rect 11104 2694 11116 2746
rect 11116 2694 11130 2746
rect 11154 2694 11168 2746
rect 11168 2694 11180 2746
rect 11180 2694 11210 2746
rect 11234 2694 11244 2746
rect 11244 2694 11290 2746
rect 10994 2692 11050 2694
rect 11074 2692 11130 2694
rect 11154 2692 11210 2694
rect 11234 2692 11290 2694
rect 17686 2746 17742 2748
rect 17766 2746 17822 2748
rect 17846 2746 17902 2748
rect 17926 2746 17982 2748
rect 17686 2694 17732 2746
rect 17732 2694 17742 2746
rect 17766 2694 17796 2746
rect 17796 2694 17808 2746
rect 17808 2694 17822 2746
rect 17846 2694 17860 2746
rect 17860 2694 17872 2746
rect 17872 2694 17902 2746
rect 17926 2694 17936 2746
rect 17936 2694 17982 2746
rect 17686 2692 17742 2694
rect 17766 2692 17822 2694
rect 17846 2692 17902 2694
rect 17926 2692 17982 2694
rect 24378 2746 24434 2748
rect 24458 2746 24514 2748
rect 24538 2746 24594 2748
rect 24618 2746 24674 2748
rect 24378 2694 24424 2746
rect 24424 2694 24434 2746
rect 24458 2694 24488 2746
rect 24488 2694 24500 2746
rect 24500 2694 24514 2746
rect 24538 2694 24552 2746
rect 24552 2694 24564 2746
rect 24564 2694 24594 2746
rect 24618 2694 24628 2746
rect 24628 2694 24674 2746
rect 24378 2692 24434 2694
rect 24458 2692 24514 2694
rect 24538 2692 24594 2694
rect 24618 2692 24674 2694
rect 7648 2202 7704 2204
rect 7728 2202 7784 2204
rect 7808 2202 7864 2204
rect 7888 2202 7944 2204
rect 7648 2150 7694 2202
rect 7694 2150 7704 2202
rect 7728 2150 7758 2202
rect 7758 2150 7770 2202
rect 7770 2150 7784 2202
rect 7808 2150 7822 2202
rect 7822 2150 7834 2202
rect 7834 2150 7864 2202
rect 7888 2150 7898 2202
rect 7898 2150 7944 2202
rect 7648 2148 7704 2150
rect 7728 2148 7784 2150
rect 7808 2148 7864 2150
rect 7888 2148 7944 2150
rect 14340 2202 14396 2204
rect 14420 2202 14476 2204
rect 14500 2202 14556 2204
rect 14580 2202 14636 2204
rect 14340 2150 14386 2202
rect 14386 2150 14396 2202
rect 14420 2150 14450 2202
rect 14450 2150 14462 2202
rect 14462 2150 14476 2202
rect 14500 2150 14514 2202
rect 14514 2150 14526 2202
rect 14526 2150 14556 2202
rect 14580 2150 14590 2202
rect 14590 2150 14636 2202
rect 14340 2148 14396 2150
rect 14420 2148 14476 2150
rect 14500 2148 14556 2150
rect 14580 2148 14636 2150
rect 21032 2202 21088 2204
rect 21112 2202 21168 2204
rect 21192 2202 21248 2204
rect 21272 2202 21328 2204
rect 21032 2150 21078 2202
rect 21078 2150 21088 2202
rect 21112 2150 21142 2202
rect 21142 2150 21154 2202
rect 21154 2150 21168 2202
rect 21192 2150 21206 2202
rect 21206 2150 21218 2202
rect 21218 2150 21248 2202
rect 21272 2150 21282 2202
rect 21282 2150 21328 2202
rect 21032 2148 21088 2150
rect 21112 2148 21168 2150
rect 21192 2148 21248 2150
rect 21272 2148 21328 2150
rect 27724 2202 27780 2204
rect 27804 2202 27860 2204
rect 27884 2202 27940 2204
rect 27964 2202 28020 2204
rect 27724 2150 27770 2202
rect 27770 2150 27780 2202
rect 27804 2150 27834 2202
rect 27834 2150 27846 2202
rect 27846 2150 27860 2202
rect 27884 2150 27898 2202
rect 27898 2150 27910 2202
rect 27910 2150 27940 2202
rect 27964 2150 27974 2202
rect 27974 2150 28020 2202
rect 27724 2148 27780 2150
rect 27804 2148 27860 2150
rect 27884 2148 27940 2150
rect 27964 2148 28020 2150
rect 3238 2080 3294 2136
<< metal3 >>
rect 0 26890 800 26920
rect 1669 26890 1735 26893
rect 0 26888 1735 26890
rect 0 26832 1674 26888
rect 1730 26832 1735 26888
rect 0 26830 1735 26832
rect 0 26800 800 26830
rect 1669 26827 1735 26830
rect 4292 26688 4608 26689
rect 4292 26624 4298 26688
rect 4362 26624 4378 26688
rect 4442 26624 4458 26688
rect 4522 26624 4538 26688
rect 4602 26624 4608 26688
rect 4292 26623 4608 26624
rect 10984 26688 11300 26689
rect 10984 26624 10990 26688
rect 11054 26624 11070 26688
rect 11134 26624 11150 26688
rect 11214 26624 11230 26688
rect 11294 26624 11300 26688
rect 10984 26623 11300 26624
rect 17676 26688 17992 26689
rect 17676 26624 17682 26688
rect 17746 26624 17762 26688
rect 17826 26624 17842 26688
rect 17906 26624 17922 26688
rect 17986 26624 17992 26688
rect 17676 26623 17992 26624
rect 24368 26688 24684 26689
rect 24368 26624 24374 26688
rect 24438 26624 24454 26688
rect 24518 26624 24534 26688
rect 24598 26624 24614 26688
rect 24678 26624 24684 26688
rect 24368 26623 24684 26624
rect 7638 26144 7954 26145
rect 7638 26080 7644 26144
rect 7708 26080 7724 26144
rect 7788 26080 7804 26144
rect 7868 26080 7884 26144
rect 7948 26080 7954 26144
rect 7638 26079 7954 26080
rect 14330 26144 14646 26145
rect 14330 26080 14336 26144
rect 14400 26080 14416 26144
rect 14480 26080 14496 26144
rect 14560 26080 14576 26144
rect 14640 26080 14646 26144
rect 14330 26079 14646 26080
rect 21022 26144 21338 26145
rect 21022 26080 21028 26144
rect 21092 26080 21108 26144
rect 21172 26080 21188 26144
rect 21252 26080 21268 26144
rect 21332 26080 21338 26144
rect 21022 26079 21338 26080
rect 27714 26144 28030 26145
rect 27714 26080 27720 26144
rect 27784 26080 27800 26144
rect 27864 26080 27880 26144
rect 27944 26080 27960 26144
rect 28024 26080 28030 26144
rect 27714 26079 28030 26080
rect 4292 25600 4608 25601
rect 4292 25536 4298 25600
rect 4362 25536 4378 25600
rect 4442 25536 4458 25600
rect 4522 25536 4538 25600
rect 4602 25536 4608 25600
rect 4292 25535 4608 25536
rect 10984 25600 11300 25601
rect 10984 25536 10990 25600
rect 11054 25536 11070 25600
rect 11134 25536 11150 25600
rect 11214 25536 11230 25600
rect 11294 25536 11300 25600
rect 10984 25535 11300 25536
rect 17676 25600 17992 25601
rect 17676 25536 17682 25600
rect 17746 25536 17762 25600
rect 17826 25536 17842 25600
rect 17906 25536 17922 25600
rect 17986 25536 17992 25600
rect 17676 25535 17992 25536
rect 24368 25600 24684 25601
rect 24368 25536 24374 25600
rect 24438 25536 24454 25600
rect 24518 25536 24534 25600
rect 24598 25536 24614 25600
rect 24678 25536 24684 25600
rect 24368 25535 24684 25536
rect 7638 25056 7954 25057
rect 7638 24992 7644 25056
rect 7708 24992 7724 25056
rect 7788 24992 7804 25056
rect 7868 24992 7884 25056
rect 7948 24992 7954 25056
rect 7638 24991 7954 24992
rect 14330 25056 14646 25057
rect 14330 24992 14336 25056
rect 14400 24992 14416 25056
rect 14480 24992 14496 25056
rect 14560 24992 14576 25056
rect 14640 24992 14646 25056
rect 14330 24991 14646 24992
rect 21022 25056 21338 25057
rect 21022 24992 21028 25056
rect 21092 24992 21108 25056
rect 21172 24992 21188 25056
rect 21252 24992 21268 25056
rect 21332 24992 21338 25056
rect 21022 24991 21338 24992
rect 27714 25056 28030 25057
rect 27714 24992 27720 25056
rect 27784 24992 27800 25056
rect 27864 24992 27880 25056
rect 27944 24992 27960 25056
rect 28024 24992 28030 25056
rect 27714 24991 28030 24992
rect 4292 24512 4608 24513
rect 4292 24448 4298 24512
rect 4362 24448 4378 24512
rect 4442 24448 4458 24512
rect 4522 24448 4538 24512
rect 4602 24448 4608 24512
rect 4292 24447 4608 24448
rect 10984 24512 11300 24513
rect 10984 24448 10990 24512
rect 11054 24448 11070 24512
rect 11134 24448 11150 24512
rect 11214 24448 11230 24512
rect 11294 24448 11300 24512
rect 10984 24447 11300 24448
rect 17676 24512 17992 24513
rect 17676 24448 17682 24512
rect 17746 24448 17762 24512
rect 17826 24448 17842 24512
rect 17906 24448 17922 24512
rect 17986 24448 17992 24512
rect 17676 24447 17992 24448
rect 24368 24512 24684 24513
rect 24368 24448 24374 24512
rect 24438 24448 24454 24512
rect 24518 24448 24534 24512
rect 24598 24448 24614 24512
rect 24678 24448 24684 24512
rect 24368 24447 24684 24448
rect 7638 23968 7954 23969
rect 7638 23904 7644 23968
rect 7708 23904 7724 23968
rect 7788 23904 7804 23968
rect 7868 23904 7884 23968
rect 7948 23904 7954 23968
rect 7638 23903 7954 23904
rect 14330 23968 14646 23969
rect 14330 23904 14336 23968
rect 14400 23904 14416 23968
rect 14480 23904 14496 23968
rect 14560 23904 14576 23968
rect 14640 23904 14646 23968
rect 14330 23903 14646 23904
rect 21022 23968 21338 23969
rect 21022 23904 21028 23968
rect 21092 23904 21108 23968
rect 21172 23904 21188 23968
rect 21252 23904 21268 23968
rect 21332 23904 21338 23968
rect 21022 23903 21338 23904
rect 27714 23968 28030 23969
rect 27714 23904 27720 23968
rect 27784 23904 27800 23968
rect 27864 23904 27880 23968
rect 27944 23904 27960 23968
rect 28024 23904 28030 23968
rect 27714 23903 28030 23904
rect 4292 23424 4608 23425
rect 0 23354 800 23384
rect 4292 23360 4298 23424
rect 4362 23360 4378 23424
rect 4442 23360 4458 23424
rect 4522 23360 4538 23424
rect 4602 23360 4608 23424
rect 4292 23359 4608 23360
rect 10984 23424 11300 23425
rect 10984 23360 10990 23424
rect 11054 23360 11070 23424
rect 11134 23360 11150 23424
rect 11214 23360 11230 23424
rect 11294 23360 11300 23424
rect 10984 23359 11300 23360
rect 17676 23424 17992 23425
rect 17676 23360 17682 23424
rect 17746 23360 17762 23424
rect 17826 23360 17842 23424
rect 17906 23360 17922 23424
rect 17986 23360 17992 23424
rect 17676 23359 17992 23360
rect 24368 23424 24684 23425
rect 24368 23360 24374 23424
rect 24438 23360 24454 23424
rect 24518 23360 24534 23424
rect 24598 23360 24614 23424
rect 24678 23360 24684 23424
rect 24368 23359 24684 23360
rect 3509 23354 3575 23357
rect 0 23352 3575 23354
rect 0 23296 3514 23352
rect 3570 23296 3575 23352
rect 0 23294 3575 23296
rect 0 23264 800 23294
rect 3509 23291 3575 23294
rect 7638 22880 7954 22881
rect 7638 22816 7644 22880
rect 7708 22816 7724 22880
rect 7788 22816 7804 22880
rect 7868 22816 7884 22880
rect 7948 22816 7954 22880
rect 7638 22815 7954 22816
rect 14330 22880 14646 22881
rect 14330 22816 14336 22880
rect 14400 22816 14416 22880
rect 14480 22816 14496 22880
rect 14560 22816 14576 22880
rect 14640 22816 14646 22880
rect 14330 22815 14646 22816
rect 21022 22880 21338 22881
rect 21022 22816 21028 22880
rect 21092 22816 21108 22880
rect 21172 22816 21188 22880
rect 21252 22816 21268 22880
rect 21332 22816 21338 22880
rect 21022 22815 21338 22816
rect 27714 22880 28030 22881
rect 27714 22816 27720 22880
rect 27784 22816 27800 22880
rect 27864 22816 27880 22880
rect 27944 22816 27960 22880
rect 28024 22816 28030 22880
rect 27714 22815 28030 22816
rect 4292 22336 4608 22337
rect 4292 22272 4298 22336
rect 4362 22272 4378 22336
rect 4442 22272 4458 22336
rect 4522 22272 4538 22336
rect 4602 22272 4608 22336
rect 4292 22271 4608 22272
rect 10984 22336 11300 22337
rect 10984 22272 10990 22336
rect 11054 22272 11070 22336
rect 11134 22272 11150 22336
rect 11214 22272 11230 22336
rect 11294 22272 11300 22336
rect 10984 22271 11300 22272
rect 17676 22336 17992 22337
rect 17676 22272 17682 22336
rect 17746 22272 17762 22336
rect 17826 22272 17842 22336
rect 17906 22272 17922 22336
rect 17986 22272 17992 22336
rect 17676 22271 17992 22272
rect 24368 22336 24684 22337
rect 24368 22272 24374 22336
rect 24438 22272 24454 22336
rect 24518 22272 24534 22336
rect 24598 22272 24614 22336
rect 24678 22272 24684 22336
rect 24368 22271 24684 22272
rect 7638 21792 7954 21793
rect 7638 21728 7644 21792
rect 7708 21728 7724 21792
rect 7788 21728 7804 21792
rect 7868 21728 7884 21792
rect 7948 21728 7954 21792
rect 7638 21727 7954 21728
rect 14330 21792 14646 21793
rect 14330 21728 14336 21792
rect 14400 21728 14416 21792
rect 14480 21728 14496 21792
rect 14560 21728 14576 21792
rect 14640 21728 14646 21792
rect 14330 21727 14646 21728
rect 21022 21792 21338 21793
rect 21022 21728 21028 21792
rect 21092 21728 21108 21792
rect 21172 21728 21188 21792
rect 21252 21728 21268 21792
rect 21332 21728 21338 21792
rect 21022 21727 21338 21728
rect 27714 21792 28030 21793
rect 27714 21728 27720 21792
rect 27784 21728 27800 21792
rect 27864 21728 27880 21792
rect 27944 21728 27960 21792
rect 28024 21728 28030 21792
rect 27714 21727 28030 21728
rect 4292 21248 4608 21249
rect 4292 21184 4298 21248
rect 4362 21184 4378 21248
rect 4442 21184 4458 21248
rect 4522 21184 4538 21248
rect 4602 21184 4608 21248
rect 4292 21183 4608 21184
rect 10984 21248 11300 21249
rect 10984 21184 10990 21248
rect 11054 21184 11070 21248
rect 11134 21184 11150 21248
rect 11214 21184 11230 21248
rect 11294 21184 11300 21248
rect 10984 21183 11300 21184
rect 17676 21248 17992 21249
rect 17676 21184 17682 21248
rect 17746 21184 17762 21248
rect 17826 21184 17842 21248
rect 17906 21184 17922 21248
rect 17986 21184 17992 21248
rect 17676 21183 17992 21184
rect 24368 21248 24684 21249
rect 24368 21184 24374 21248
rect 24438 21184 24454 21248
rect 24518 21184 24534 21248
rect 24598 21184 24614 21248
rect 24678 21184 24684 21248
rect 24368 21183 24684 21184
rect 7638 20704 7954 20705
rect 7638 20640 7644 20704
rect 7708 20640 7724 20704
rect 7788 20640 7804 20704
rect 7868 20640 7884 20704
rect 7948 20640 7954 20704
rect 7638 20639 7954 20640
rect 14330 20704 14646 20705
rect 14330 20640 14336 20704
rect 14400 20640 14416 20704
rect 14480 20640 14496 20704
rect 14560 20640 14576 20704
rect 14640 20640 14646 20704
rect 14330 20639 14646 20640
rect 21022 20704 21338 20705
rect 21022 20640 21028 20704
rect 21092 20640 21108 20704
rect 21172 20640 21188 20704
rect 21252 20640 21268 20704
rect 21332 20640 21338 20704
rect 21022 20639 21338 20640
rect 27714 20704 28030 20705
rect 27714 20640 27720 20704
rect 27784 20640 27800 20704
rect 27864 20640 27880 20704
rect 27944 20640 27960 20704
rect 28024 20640 28030 20704
rect 27714 20639 28030 20640
rect 4292 20160 4608 20161
rect 4292 20096 4298 20160
rect 4362 20096 4378 20160
rect 4442 20096 4458 20160
rect 4522 20096 4538 20160
rect 4602 20096 4608 20160
rect 4292 20095 4608 20096
rect 10984 20160 11300 20161
rect 10984 20096 10990 20160
rect 11054 20096 11070 20160
rect 11134 20096 11150 20160
rect 11214 20096 11230 20160
rect 11294 20096 11300 20160
rect 10984 20095 11300 20096
rect 17676 20160 17992 20161
rect 17676 20096 17682 20160
rect 17746 20096 17762 20160
rect 17826 20096 17842 20160
rect 17906 20096 17922 20160
rect 17986 20096 17992 20160
rect 17676 20095 17992 20096
rect 24368 20160 24684 20161
rect 24368 20096 24374 20160
rect 24438 20096 24454 20160
rect 24518 20096 24534 20160
rect 24598 20096 24614 20160
rect 24678 20096 24684 20160
rect 24368 20095 24684 20096
rect 0 19818 800 19848
rect 1669 19818 1735 19821
rect 0 19816 1735 19818
rect 0 19760 1674 19816
rect 1730 19760 1735 19816
rect 0 19758 1735 19760
rect 0 19728 800 19758
rect 1669 19755 1735 19758
rect 7638 19616 7954 19617
rect 7638 19552 7644 19616
rect 7708 19552 7724 19616
rect 7788 19552 7804 19616
rect 7868 19552 7884 19616
rect 7948 19552 7954 19616
rect 7638 19551 7954 19552
rect 14330 19616 14646 19617
rect 14330 19552 14336 19616
rect 14400 19552 14416 19616
rect 14480 19552 14496 19616
rect 14560 19552 14576 19616
rect 14640 19552 14646 19616
rect 14330 19551 14646 19552
rect 21022 19616 21338 19617
rect 21022 19552 21028 19616
rect 21092 19552 21108 19616
rect 21172 19552 21188 19616
rect 21252 19552 21268 19616
rect 21332 19552 21338 19616
rect 21022 19551 21338 19552
rect 27714 19616 28030 19617
rect 27714 19552 27720 19616
rect 27784 19552 27800 19616
rect 27864 19552 27880 19616
rect 27944 19552 27960 19616
rect 28024 19552 28030 19616
rect 27714 19551 28030 19552
rect 4292 19072 4608 19073
rect 4292 19008 4298 19072
rect 4362 19008 4378 19072
rect 4442 19008 4458 19072
rect 4522 19008 4538 19072
rect 4602 19008 4608 19072
rect 4292 19007 4608 19008
rect 10984 19072 11300 19073
rect 10984 19008 10990 19072
rect 11054 19008 11070 19072
rect 11134 19008 11150 19072
rect 11214 19008 11230 19072
rect 11294 19008 11300 19072
rect 10984 19007 11300 19008
rect 17676 19072 17992 19073
rect 17676 19008 17682 19072
rect 17746 19008 17762 19072
rect 17826 19008 17842 19072
rect 17906 19008 17922 19072
rect 17986 19008 17992 19072
rect 17676 19007 17992 19008
rect 24368 19072 24684 19073
rect 24368 19008 24374 19072
rect 24438 19008 24454 19072
rect 24518 19008 24534 19072
rect 24598 19008 24614 19072
rect 24678 19008 24684 19072
rect 24368 19007 24684 19008
rect 7638 18528 7954 18529
rect 7638 18464 7644 18528
rect 7708 18464 7724 18528
rect 7788 18464 7804 18528
rect 7868 18464 7884 18528
rect 7948 18464 7954 18528
rect 7638 18463 7954 18464
rect 14330 18528 14646 18529
rect 14330 18464 14336 18528
rect 14400 18464 14416 18528
rect 14480 18464 14496 18528
rect 14560 18464 14576 18528
rect 14640 18464 14646 18528
rect 14330 18463 14646 18464
rect 21022 18528 21338 18529
rect 21022 18464 21028 18528
rect 21092 18464 21108 18528
rect 21172 18464 21188 18528
rect 21252 18464 21268 18528
rect 21332 18464 21338 18528
rect 21022 18463 21338 18464
rect 27714 18528 28030 18529
rect 27714 18464 27720 18528
rect 27784 18464 27800 18528
rect 27864 18464 27880 18528
rect 27944 18464 27960 18528
rect 28024 18464 28030 18528
rect 27714 18463 28030 18464
rect 4292 17984 4608 17985
rect 4292 17920 4298 17984
rect 4362 17920 4378 17984
rect 4442 17920 4458 17984
rect 4522 17920 4538 17984
rect 4602 17920 4608 17984
rect 4292 17919 4608 17920
rect 10984 17984 11300 17985
rect 10984 17920 10990 17984
rect 11054 17920 11070 17984
rect 11134 17920 11150 17984
rect 11214 17920 11230 17984
rect 11294 17920 11300 17984
rect 10984 17919 11300 17920
rect 17676 17984 17992 17985
rect 17676 17920 17682 17984
rect 17746 17920 17762 17984
rect 17826 17920 17842 17984
rect 17906 17920 17922 17984
rect 17986 17920 17992 17984
rect 17676 17919 17992 17920
rect 24368 17984 24684 17985
rect 24368 17920 24374 17984
rect 24438 17920 24454 17984
rect 24518 17920 24534 17984
rect 24598 17920 24614 17984
rect 24678 17920 24684 17984
rect 24368 17919 24684 17920
rect 7638 17440 7954 17441
rect 7638 17376 7644 17440
rect 7708 17376 7724 17440
rect 7788 17376 7804 17440
rect 7868 17376 7884 17440
rect 7948 17376 7954 17440
rect 7638 17375 7954 17376
rect 14330 17440 14646 17441
rect 14330 17376 14336 17440
rect 14400 17376 14416 17440
rect 14480 17376 14496 17440
rect 14560 17376 14576 17440
rect 14640 17376 14646 17440
rect 14330 17375 14646 17376
rect 21022 17440 21338 17441
rect 21022 17376 21028 17440
rect 21092 17376 21108 17440
rect 21172 17376 21188 17440
rect 21252 17376 21268 17440
rect 21332 17376 21338 17440
rect 21022 17375 21338 17376
rect 27714 17440 28030 17441
rect 27714 17376 27720 17440
rect 27784 17376 27800 17440
rect 27864 17376 27880 17440
rect 27944 17376 27960 17440
rect 28024 17376 28030 17440
rect 27714 17375 28030 17376
rect 12709 17098 12775 17101
rect 13905 17098 13971 17101
rect 12709 17096 13971 17098
rect 12709 17040 12714 17096
rect 12770 17040 13910 17096
rect 13966 17040 13971 17096
rect 12709 17038 13971 17040
rect 12709 17035 12775 17038
rect 13905 17035 13971 17038
rect 4292 16896 4608 16897
rect 4292 16832 4298 16896
rect 4362 16832 4378 16896
rect 4442 16832 4458 16896
rect 4522 16832 4538 16896
rect 4602 16832 4608 16896
rect 4292 16831 4608 16832
rect 10984 16896 11300 16897
rect 10984 16832 10990 16896
rect 11054 16832 11070 16896
rect 11134 16832 11150 16896
rect 11214 16832 11230 16896
rect 11294 16832 11300 16896
rect 10984 16831 11300 16832
rect 17676 16896 17992 16897
rect 17676 16832 17682 16896
rect 17746 16832 17762 16896
rect 17826 16832 17842 16896
rect 17906 16832 17922 16896
rect 17986 16832 17992 16896
rect 17676 16831 17992 16832
rect 24368 16896 24684 16897
rect 24368 16832 24374 16896
rect 24438 16832 24454 16896
rect 24518 16832 24534 16896
rect 24598 16832 24614 16896
rect 24678 16832 24684 16896
rect 24368 16831 24684 16832
rect 14917 16554 14983 16557
rect 14782 16552 14983 16554
rect 14782 16496 14922 16552
rect 14978 16496 14983 16552
rect 14782 16494 14983 16496
rect 7638 16352 7954 16353
rect 0 16282 800 16312
rect 7638 16288 7644 16352
rect 7708 16288 7724 16352
rect 7788 16288 7804 16352
rect 7868 16288 7884 16352
rect 7948 16288 7954 16352
rect 7638 16287 7954 16288
rect 14330 16352 14646 16353
rect 14330 16288 14336 16352
rect 14400 16288 14416 16352
rect 14480 16288 14496 16352
rect 14560 16288 14576 16352
rect 14640 16288 14646 16352
rect 14330 16287 14646 16288
rect 1577 16282 1643 16285
rect 0 16280 1643 16282
rect 0 16224 1582 16280
rect 1638 16224 1643 16280
rect 0 16222 1643 16224
rect 0 16192 800 16222
rect 1577 16219 1643 16222
rect 14782 16013 14842 16494
rect 14917 16491 14983 16494
rect 21022 16352 21338 16353
rect 21022 16288 21028 16352
rect 21092 16288 21108 16352
rect 21172 16288 21188 16352
rect 21252 16288 21268 16352
rect 21332 16288 21338 16352
rect 21022 16287 21338 16288
rect 27714 16352 28030 16353
rect 27714 16288 27720 16352
rect 27784 16288 27800 16352
rect 27864 16288 27880 16352
rect 27944 16288 27960 16352
rect 28024 16288 28030 16352
rect 27714 16287 28030 16288
rect 14733 16008 14842 16013
rect 14733 15952 14738 16008
rect 14794 15952 14842 16008
rect 14733 15950 14842 15952
rect 14733 15947 14799 15950
rect 4292 15808 4608 15809
rect 4292 15744 4298 15808
rect 4362 15744 4378 15808
rect 4442 15744 4458 15808
rect 4522 15744 4538 15808
rect 4602 15744 4608 15808
rect 4292 15743 4608 15744
rect 10984 15808 11300 15809
rect 10984 15744 10990 15808
rect 11054 15744 11070 15808
rect 11134 15744 11150 15808
rect 11214 15744 11230 15808
rect 11294 15744 11300 15808
rect 10984 15743 11300 15744
rect 17676 15808 17992 15809
rect 17676 15744 17682 15808
rect 17746 15744 17762 15808
rect 17826 15744 17842 15808
rect 17906 15744 17922 15808
rect 17986 15744 17992 15808
rect 17676 15743 17992 15744
rect 24368 15808 24684 15809
rect 24368 15744 24374 15808
rect 24438 15744 24454 15808
rect 24518 15744 24534 15808
rect 24598 15744 24614 15808
rect 24678 15744 24684 15808
rect 24368 15743 24684 15744
rect 7638 15264 7954 15265
rect 7638 15200 7644 15264
rect 7708 15200 7724 15264
rect 7788 15200 7804 15264
rect 7868 15200 7884 15264
rect 7948 15200 7954 15264
rect 7638 15199 7954 15200
rect 14330 15264 14646 15265
rect 14330 15200 14336 15264
rect 14400 15200 14416 15264
rect 14480 15200 14496 15264
rect 14560 15200 14576 15264
rect 14640 15200 14646 15264
rect 14330 15199 14646 15200
rect 21022 15264 21338 15265
rect 21022 15200 21028 15264
rect 21092 15200 21108 15264
rect 21172 15200 21188 15264
rect 21252 15200 21268 15264
rect 21332 15200 21338 15264
rect 21022 15199 21338 15200
rect 27714 15264 28030 15265
rect 27714 15200 27720 15264
rect 27784 15200 27800 15264
rect 27864 15200 27880 15264
rect 27944 15200 27960 15264
rect 28024 15200 28030 15264
rect 27714 15199 28030 15200
rect 4292 14720 4608 14721
rect 4292 14656 4298 14720
rect 4362 14656 4378 14720
rect 4442 14656 4458 14720
rect 4522 14656 4538 14720
rect 4602 14656 4608 14720
rect 4292 14655 4608 14656
rect 10984 14720 11300 14721
rect 10984 14656 10990 14720
rect 11054 14656 11070 14720
rect 11134 14656 11150 14720
rect 11214 14656 11230 14720
rect 11294 14656 11300 14720
rect 10984 14655 11300 14656
rect 17676 14720 17992 14721
rect 17676 14656 17682 14720
rect 17746 14656 17762 14720
rect 17826 14656 17842 14720
rect 17906 14656 17922 14720
rect 17986 14656 17992 14720
rect 17676 14655 17992 14656
rect 24368 14720 24684 14721
rect 24368 14656 24374 14720
rect 24438 14656 24454 14720
rect 24518 14656 24534 14720
rect 24598 14656 24614 14720
rect 24678 14656 24684 14720
rect 24368 14655 24684 14656
rect 7638 14176 7954 14177
rect 7638 14112 7644 14176
rect 7708 14112 7724 14176
rect 7788 14112 7804 14176
rect 7868 14112 7884 14176
rect 7948 14112 7954 14176
rect 7638 14111 7954 14112
rect 14330 14176 14646 14177
rect 14330 14112 14336 14176
rect 14400 14112 14416 14176
rect 14480 14112 14496 14176
rect 14560 14112 14576 14176
rect 14640 14112 14646 14176
rect 14330 14111 14646 14112
rect 21022 14176 21338 14177
rect 21022 14112 21028 14176
rect 21092 14112 21108 14176
rect 21172 14112 21188 14176
rect 21252 14112 21268 14176
rect 21332 14112 21338 14176
rect 21022 14111 21338 14112
rect 27714 14176 28030 14177
rect 27714 14112 27720 14176
rect 27784 14112 27800 14176
rect 27864 14112 27880 14176
rect 27944 14112 27960 14176
rect 28024 14112 28030 14176
rect 27714 14111 28030 14112
rect 12433 13698 12499 13701
rect 14089 13698 14155 13701
rect 12433 13696 14155 13698
rect 12433 13640 12438 13696
rect 12494 13640 14094 13696
rect 14150 13640 14155 13696
rect 12433 13638 14155 13640
rect 12433 13635 12499 13638
rect 14089 13635 14155 13638
rect 4292 13632 4608 13633
rect 4292 13568 4298 13632
rect 4362 13568 4378 13632
rect 4442 13568 4458 13632
rect 4522 13568 4538 13632
rect 4602 13568 4608 13632
rect 4292 13567 4608 13568
rect 10984 13632 11300 13633
rect 10984 13568 10990 13632
rect 11054 13568 11070 13632
rect 11134 13568 11150 13632
rect 11214 13568 11230 13632
rect 11294 13568 11300 13632
rect 10984 13567 11300 13568
rect 17676 13632 17992 13633
rect 17676 13568 17682 13632
rect 17746 13568 17762 13632
rect 17826 13568 17842 13632
rect 17906 13568 17922 13632
rect 17986 13568 17992 13632
rect 17676 13567 17992 13568
rect 24368 13632 24684 13633
rect 24368 13568 24374 13632
rect 24438 13568 24454 13632
rect 24518 13568 24534 13632
rect 24598 13568 24614 13632
rect 24678 13568 24684 13632
rect 24368 13567 24684 13568
rect 12433 13562 12499 13565
rect 12709 13562 12775 13565
rect 12433 13560 12775 13562
rect 12433 13504 12438 13560
rect 12494 13504 12714 13560
rect 12770 13504 12775 13560
rect 12433 13502 12775 13504
rect 12433 13499 12499 13502
rect 12709 13499 12775 13502
rect 9305 13290 9371 13293
rect 17493 13290 17559 13293
rect 9305 13288 17559 13290
rect 9305 13232 9310 13288
rect 9366 13232 17498 13288
rect 17554 13232 17559 13288
rect 9305 13230 17559 13232
rect 9305 13227 9371 13230
rect 17493 13227 17559 13230
rect 11881 13154 11947 13157
rect 13997 13154 14063 13157
rect 11881 13152 14063 13154
rect 11881 13096 11886 13152
rect 11942 13096 14002 13152
rect 14058 13096 14063 13152
rect 11881 13094 14063 13096
rect 11881 13091 11947 13094
rect 13997 13091 14063 13094
rect 7638 13088 7954 13089
rect 7638 13024 7644 13088
rect 7708 13024 7724 13088
rect 7788 13024 7804 13088
rect 7868 13024 7884 13088
rect 7948 13024 7954 13088
rect 7638 13023 7954 13024
rect 14330 13088 14646 13089
rect 14330 13024 14336 13088
rect 14400 13024 14416 13088
rect 14480 13024 14496 13088
rect 14560 13024 14576 13088
rect 14640 13024 14646 13088
rect 14330 13023 14646 13024
rect 21022 13088 21338 13089
rect 21022 13024 21028 13088
rect 21092 13024 21108 13088
rect 21172 13024 21188 13088
rect 21252 13024 21268 13088
rect 21332 13024 21338 13088
rect 21022 13023 21338 13024
rect 27714 13088 28030 13089
rect 27714 13024 27720 13088
rect 27784 13024 27800 13088
rect 27864 13024 27880 13088
rect 27944 13024 27960 13088
rect 28024 13024 28030 13088
rect 27714 13023 28030 13024
rect 12065 13018 12131 13021
rect 13721 13018 13787 13021
rect 12065 13016 13787 13018
rect 12065 12960 12070 13016
rect 12126 12960 13726 13016
rect 13782 12960 13787 13016
rect 12065 12958 13787 12960
rect 12065 12955 12131 12958
rect 13721 12955 13787 12958
rect 13537 12882 13603 12885
rect 20437 12882 20503 12885
rect 13537 12880 20503 12882
rect 13537 12824 13542 12880
rect 13598 12824 20442 12880
rect 20498 12824 20503 12880
rect 13537 12822 20503 12824
rect 13537 12819 13603 12822
rect 20437 12819 20503 12822
rect 0 12746 800 12776
rect 1577 12746 1643 12749
rect 0 12744 1643 12746
rect 0 12688 1582 12744
rect 1638 12688 1643 12744
rect 0 12686 1643 12688
rect 0 12656 800 12686
rect 1577 12683 1643 12686
rect 12893 12610 12959 12613
rect 14549 12610 14615 12613
rect 12893 12608 14615 12610
rect 12893 12552 12898 12608
rect 12954 12552 14554 12608
rect 14610 12552 14615 12608
rect 12893 12550 14615 12552
rect 12893 12547 12959 12550
rect 14549 12547 14615 12550
rect 4292 12544 4608 12545
rect 4292 12480 4298 12544
rect 4362 12480 4378 12544
rect 4442 12480 4458 12544
rect 4522 12480 4538 12544
rect 4602 12480 4608 12544
rect 4292 12479 4608 12480
rect 10984 12544 11300 12545
rect 10984 12480 10990 12544
rect 11054 12480 11070 12544
rect 11134 12480 11150 12544
rect 11214 12480 11230 12544
rect 11294 12480 11300 12544
rect 10984 12479 11300 12480
rect 17676 12544 17992 12545
rect 17676 12480 17682 12544
rect 17746 12480 17762 12544
rect 17826 12480 17842 12544
rect 17906 12480 17922 12544
rect 17986 12480 17992 12544
rect 17676 12479 17992 12480
rect 24368 12544 24684 12545
rect 24368 12480 24374 12544
rect 24438 12480 24454 12544
rect 24518 12480 24534 12544
rect 24598 12480 24614 12544
rect 24678 12480 24684 12544
rect 24368 12479 24684 12480
rect 7638 12000 7954 12001
rect 7638 11936 7644 12000
rect 7708 11936 7724 12000
rect 7788 11936 7804 12000
rect 7868 11936 7884 12000
rect 7948 11936 7954 12000
rect 7638 11935 7954 11936
rect 14330 12000 14646 12001
rect 14330 11936 14336 12000
rect 14400 11936 14416 12000
rect 14480 11936 14496 12000
rect 14560 11936 14576 12000
rect 14640 11936 14646 12000
rect 14330 11935 14646 11936
rect 21022 12000 21338 12001
rect 21022 11936 21028 12000
rect 21092 11936 21108 12000
rect 21172 11936 21188 12000
rect 21252 11936 21268 12000
rect 21332 11936 21338 12000
rect 21022 11935 21338 11936
rect 27714 12000 28030 12001
rect 27714 11936 27720 12000
rect 27784 11936 27800 12000
rect 27864 11936 27880 12000
rect 27944 11936 27960 12000
rect 28024 11936 28030 12000
rect 27714 11935 28030 11936
rect 4292 11456 4608 11457
rect 4292 11392 4298 11456
rect 4362 11392 4378 11456
rect 4442 11392 4458 11456
rect 4522 11392 4538 11456
rect 4602 11392 4608 11456
rect 4292 11391 4608 11392
rect 10984 11456 11300 11457
rect 10984 11392 10990 11456
rect 11054 11392 11070 11456
rect 11134 11392 11150 11456
rect 11214 11392 11230 11456
rect 11294 11392 11300 11456
rect 10984 11391 11300 11392
rect 17676 11456 17992 11457
rect 17676 11392 17682 11456
rect 17746 11392 17762 11456
rect 17826 11392 17842 11456
rect 17906 11392 17922 11456
rect 17986 11392 17992 11456
rect 17676 11391 17992 11392
rect 24368 11456 24684 11457
rect 24368 11392 24374 11456
rect 24438 11392 24454 11456
rect 24518 11392 24534 11456
rect 24598 11392 24614 11456
rect 24678 11392 24684 11456
rect 24368 11391 24684 11392
rect 7638 10912 7954 10913
rect 7638 10848 7644 10912
rect 7708 10848 7724 10912
rect 7788 10848 7804 10912
rect 7868 10848 7884 10912
rect 7948 10848 7954 10912
rect 7638 10847 7954 10848
rect 14330 10912 14646 10913
rect 14330 10848 14336 10912
rect 14400 10848 14416 10912
rect 14480 10848 14496 10912
rect 14560 10848 14576 10912
rect 14640 10848 14646 10912
rect 14330 10847 14646 10848
rect 21022 10912 21338 10913
rect 21022 10848 21028 10912
rect 21092 10848 21108 10912
rect 21172 10848 21188 10912
rect 21252 10848 21268 10912
rect 21332 10848 21338 10912
rect 21022 10847 21338 10848
rect 27714 10912 28030 10913
rect 27714 10848 27720 10912
rect 27784 10848 27800 10912
rect 27864 10848 27880 10912
rect 27944 10848 27960 10912
rect 28024 10848 28030 10912
rect 27714 10847 28030 10848
rect 4292 10368 4608 10369
rect 4292 10304 4298 10368
rect 4362 10304 4378 10368
rect 4442 10304 4458 10368
rect 4522 10304 4538 10368
rect 4602 10304 4608 10368
rect 4292 10303 4608 10304
rect 10984 10368 11300 10369
rect 10984 10304 10990 10368
rect 11054 10304 11070 10368
rect 11134 10304 11150 10368
rect 11214 10304 11230 10368
rect 11294 10304 11300 10368
rect 10984 10303 11300 10304
rect 17676 10368 17992 10369
rect 17676 10304 17682 10368
rect 17746 10304 17762 10368
rect 17826 10304 17842 10368
rect 17906 10304 17922 10368
rect 17986 10304 17992 10368
rect 17676 10303 17992 10304
rect 24368 10368 24684 10369
rect 24368 10304 24374 10368
rect 24438 10304 24454 10368
rect 24518 10304 24534 10368
rect 24598 10304 24614 10368
rect 24678 10304 24684 10368
rect 24368 10303 24684 10304
rect 7638 9824 7954 9825
rect 7638 9760 7644 9824
rect 7708 9760 7724 9824
rect 7788 9760 7804 9824
rect 7868 9760 7884 9824
rect 7948 9760 7954 9824
rect 7638 9759 7954 9760
rect 14330 9824 14646 9825
rect 14330 9760 14336 9824
rect 14400 9760 14416 9824
rect 14480 9760 14496 9824
rect 14560 9760 14576 9824
rect 14640 9760 14646 9824
rect 14330 9759 14646 9760
rect 21022 9824 21338 9825
rect 21022 9760 21028 9824
rect 21092 9760 21108 9824
rect 21172 9760 21188 9824
rect 21252 9760 21268 9824
rect 21332 9760 21338 9824
rect 21022 9759 21338 9760
rect 27714 9824 28030 9825
rect 27714 9760 27720 9824
rect 27784 9760 27800 9824
rect 27864 9760 27880 9824
rect 27944 9760 27960 9824
rect 28024 9760 28030 9824
rect 27714 9759 28030 9760
rect 4292 9280 4608 9281
rect 0 9210 800 9240
rect 4292 9216 4298 9280
rect 4362 9216 4378 9280
rect 4442 9216 4458 9280
rect 4522 9216 4538 9280
rect 4602 9216 4608 9280
rect 4292 9215 4608 9216
rect 10984 9280 11300 9281
rect 10984 9216 10990 9280
rect 11054 9216 11070 9280
rect 11134 9216 11150 9280
rect 11214 9216 11230 9280
rect 11294 9216 11300 9280
rect 10984 9215 11300 9216
rect 17676 9280 17992 9281
rect 17676 9216 17682 9280
rect 17746 9216 17762 9280
rect 17826 9216 17842 9280
rect 17906 9216 17922 9280
rect 17986 9216 17992 9280
rect 17676 9215 17992 9216
rect 24368 9280 24684 9281
rect 24368 9216 24374 9280
rect 24438 9216 24454 9280
rect 24518 9216 24534 9280
rect 24598 9216 24614 9280
rect 24678 9216 24684 9280
rect 24368 9215 24684 9216
rect 2957 9210 3023 9213
rect 0 9208 3023 9210
rect 0 9152 2962 9208
rect 3018 9152 3023 9208
rect 0 9150 3023 9152
rect 0 9120 800 9150
rect 2957 9147 3023 9150
rect 7638 8736 7954 8737
rect 7638 8672 7644 8736
rect 7708 8672 7724 8736
rect 7788 8672 7804 8736
rect 7868 8672 7884 8736
rect 7948 8672 7954 8736
rect 7638 8671 7954 8672
rect 14330 8736 14646 8737
rect 14330 8672 14336 8736
rect 14400 8672 14416 8736
rect 14480 8672 14496 8736
rect 14560 8672 14576 8736
rect 14640 8672 14646 8736
rect 14330 8671 14646 8672
rect 21022 8736 21338 8737
rect 21022 8672 21028 8736
rect 21092 8672 21108 8736
rect 21172 8672 21188 8736
rect 21252 8672 21268 8736
rect 21332 8672 21338 8736
rect 21022 8671 21338 8672
rect 27714 8736 28030 8737
rect 27714 8672 27720 8736
rect 27784 8672 27800 8736
rect 27864 8672 27880 8736
rect 27944 8672 27960 8736
rect 28024 8672 28030 8736
rect 27714 8671 28030 8672
rect 4292 8192 4608 8193
rect 4292 8128 4298 8192
rect 4362 8128 4378 8192
rect 4442 8128 4458 8192
rect 4522 8128 4538 8192
rect 4602 8128 4608 8192
rect 4292 8127 4608 8128
rect 10984 8192 11300 8193
rect 10984 8128 10990 8192
rect 11054 8128 11070 8192
rect 11134 8128 11150 8192
rect 11214 8128 11230 8192
rect 11294 8128 11300 8192
rect 10984 8127 11300 8128
rect 17676 8192 17992 8193
rect 17676 8128 17682 8192
rect 17746 8128 17762 8192
rect 17826 8128 17842 8192
rect 17906 8128 17922 8192
rect 17986 8128 17992 8192
rect 17676 8127 17992 8128
rect 24368 8192 24684 8193
rect 24368 8128 24374 8192
rect 24438 8128 24454 8192
rect 24518 8128 24534 8192
rect 24598 8128 24614 8192
rect 24678 8128 24684 8192
rect 24368 8127 24684 8128
rect 7638 7648 7954 7649
rect 7638 7584 7644 7648
rect 7708 7584 7724 7648
rect 7788 7584 7804 7648
rect 7868 7584 7884 7648
rect 7948 7584 7954 7648
rect 7638 7583 7954 7584
rect 14330 7648 14646 7649
rect 14330 7584 14336 7648
rect 14400 7584 14416 7648
rect 14480 7584 14496 7648
rect 14560 7584 14576 7648
rect 14640 7584 14646 7648
rect 14330 7583 14646 7584
rect 21022 7648 21338 7649
rect 21022 7584 21028 7648
rect 21092 7584 21108 7648
rect 21172 7584 21188 7648
rect 21252 7584 21268 7648
rect 21332 7584 21338 7648
rect 21022 7583 21338 7584
rect 27714 7648 28030 7649
rect 27714 7584 27720 7648
rect 27784 7584 27800 7648
rect 27864 7584 27880 7648
rect 27944 7584 27960 7648
rect 28024 7584 28030 7648
rect 27714 7583 28030 7584
rect 4292 7104 4608 7105
rect 4292 7040 4298 7104
rect 4362 7040 4378 7104
rect 4442 7040 4458 7104
rect 4522 7040 4538 7104
rect 4602 7040 4608 7104
rect 4292 7039 4608 7040
rect 10984 7104 11300 7105
rect 10984 7040 10990 7104
rect 11054 7040 11070 7104
rect 11134 7040 11150 7104
rect 11214 7040 11230 7104
rect 11294 7040 11300 7104
rect 10984 7039 11300 7040
rect 17676 7104 17992 7105
rect 17676 7040 17682 7104
rect 17746 7040 17762 7104
rect 17826 7040 17842 7104
rect 17906 7040 17922 7104
rect 17986 7040 17992 7104
rect 17676 7039 17992 7040
rect 24368 7104 24684 7105
rect 24368 7040 24374 7104
rect 24438 7040 24454 7104
rect 24518 7040 24534 7104
rect 24598 7040 24614 7104
rect 24678 7040 24684 7104
rect 24368 7039 24684 7040
rect 7638 6560 7954 6561
rect 7638 6496 7644 6560
rect 7708 6496 7724 6560
rect 7788 6496 7804 6560
rect 7868 6496 7884 6560
rect 7948 6496 7954 6560
rect 7638 6495 7954 6496
rect 14330 6560 14646 6561
rect 14330 6496 14336 6560
rect 14400 6496 14416 6560
rect 14480 6496 14496 6560
rect 14560 6496 14576 6560
rect 14640 6496 14646 6560
rect 14330 6495 14646 6496
rect 21022 6560 21338 6561
rect 21022 6496 21028 6560
rect 21092 6496 21108 6560
rect 21172 6496 21188 6560
rect 21252 6496 21268 6560
rect 21332 6496 21338 6560
rect 21022 6495 21338 6496
rect 27714 6560 28030 6561
rect 27714 6496 27720 6560
rect 27784 6496 27800 6560
rect 27864 6496 27880 6560
rect 27944 6496 27960 6560
rect 28024 6496 28030 6560
rect 27714 6495 28030 6496
rect 4292 6016 4608 6017
rect 4292 5952 4298 6016
rect 4362 5952 4378 6016
rect 4442 5952 4458 6016
rect 4522 5952 4538 6016
rect 4602 5952 4608 6016
rect 4292 5951 4608 5952
rect 10984 6016 11300 6017
rect 10984 5952 10990 6016
rect 11054 5952 11070 6016
rect 11134 5952 11150 6016
rect 11214 5952 11230 6016
rect 11294 5952 11300 6016
rect 10984 5951 11300 5952
rect 17676 6016 17992 6017
rect 17676 5952 17682 6016
rect 17746 5952 17762 6016
rect 17826 5952 17842 6016
rect 17906 5952 17922 6016
rect 17986 5952 17992 6016
rect 17676 5951 17992 5952
rect 24368 6016 24684 6017
rect 24368 5952 24374 6016
rect 24438 5952 24454 6016
rect 24518 5952 24534 6016
rect 24598 5952 24614 6016
rect 24678 5952 24684 6016
rect 24368 5951 24684 5952
rect 0 5674 800 5704
rect 1485 5674 1551 5677
rect 0 5672 1551 5674
rect 0 5616 1490 5672
rect 1546 5616 1551 5672
rect 0 5614 1551 5616
rect 0 5584 800 5614
rect 1485 5611 1551 5614
rect 7638 5472 7954 5473
rect 7638 5408 7644 5472
rect 7708 5408 7724 5472
rect 7788 5408 7804 5472
rect 7868 5408 7884 5472
rect 7948 5408 7954 5472
rect 7638 5407 7954 5408
rect 14330 5472 14646 5473
rect 14330 5408 14336 5472
rect 14400 5408 14416 5472
rect 14480 5408 14496 5472
rect 14560 5408 14576 5472
rect 14640 5408 14646 5472
rect 14330 5407 14646 5408
rect 21022 5472 21338 5473
rect 21022 5408 21028 5472
rect 21092 5408 21108 5472
rect 21172 5408 21188 5472
rect 21252 5408 21268 5472
rect 21332 5408 21338 5472
rect 21022 5407 21338 5408
rect 27714 5472 28030 5473
rect 27714 5408 27720 5472
rect 27784 5408 27800 5472
rect 27864 5408 27880 5472
rect 27944 5408 27960 5472
rect 28024 5408 28030 5472
rect 27714 5407 28030 5408
rect 4292 4928 4608 4929
rect 4292 4864 4298 4928
rect 4362 4864 4378 4928
rect 4442 4864 4458 4928
rect 4522 4864 4538 4928
rect 4602 4864 4608 4928
rect 4292 4863 4608 4864
rect 10984 4928 11300 4929
rect 10984 4864 10990 4928
rect 11054 4864 11070 4928
rect 11134 4864 11150 4928
rect 11214 4864 11230 4928
rect 11294 4864 11300 4928
rect 10984 4863 11300 4864
rect 17676 4928 17992 4929
rect 17676 4864 17682 4928
rect 17746 4864 17762 4928
rect 17826 4864 17842 4928
rect 17906 4864 17922 4928
rect 17986 4864 17992 4928
rect 17676 4863 17992 4864
rect 24368 4928 24684 4929
rect 24368 4864 24374 4928
rect 24438 4864 24454 4928
rect 24518 4864 24534 4928
rect 24598 4864 24614 4928
rect 24678 4864 24684 4928
rect 24368 4863 24684 4864
rect 7638 4384 7954 4385
rect 7638 4320 7644 4384
rect 7708 4320 7724 4384
rect 7788 4320 7804 4384
rect 7868 4320 7884 4384
rect 7948 4320 7954 4384
rect 7638 4319 7954 4320
rect 14330 4384 14646 4385
rect 14330 4320 14336 4384
rect 14400 4320 14416 4384
rect 14480 4320 14496 4384
rect 14560 4320 14576 4384
rect 14640 4320 14646 4384
rect 14330 4319 14646 4320
rect 21022 4384 21338 4385
rect 21022 4320 21028 4384
rect 21092 4320 21108 4384
rect 21172 4320 21188 4384
rect 21252 4320 21268 4384
rect 21332 4320 21338 4384
rect 21022 4319 21338 4320
rect 27714 4384 28030 4385
rect 27714 4320 27720 4384
rect 27784 4320 27800 4384
rect 27864 4320 27880 4384
rect 27944 4320 27960 4384
rect 28024 4320 28030 4384
rect 27714 4319 28030 4320
rect 4292 3840 4608 3841
rect 4292 3776 4298 3840
rect 4362 3776 4378 3840
rect 4442 3776 4458 3840
rect 4522 3776 4538 3840
rect 4602 3776 4608 3840
rect 4292 3775 4608 3776
rect 10984 3840 11300 3841
rect 10984 3776 10990 3840
rect 11054 3776 11070 3840
rect 11134 3776 11150 3840
rect 11214 3776 11230 3840
rect 11294 3776 11300 3840
rect 10984 3775 11300 3776
rect 17676 3840 17992 3841
rect 17676 3776 17682 3840
rect 17746 3776 17762 3840
rect 17826 3776 17842 3840
rect 17906 3776 17922 3840
rect 17986 3776 17992 3840
rect 17676 3775 17992 3776
rect 24368 3840 24684 3841
rect 24368 3776 24374 3840
rect 24438 3776 24454 3840
rect 24518 3776 24534 3840
rect 24598 3776 24614 3840
rect 24678 3776 24684 3840
rect 24368 3775 24684 3776
rect 7638 3296 7954 3297
rect 7638 3232 7644 3296
rect 7708 3232 7724 3296
rect 7788 3232 7804 3296
rect 7868 3232 7884 3296
rect 7948 3232 7954 3296
rect 7638 3231 7954 3232
rect 14330 3296 14646 3297
rect 14330 3232 14336 3296
rect 14400 3232 14416 3296
rect 14480 3232 14496 3296
rect 14560 3232 14576 3296
rect 14640 3232 14646 3296
rect 14330 3231 14646 3232
rect 21022 3296 21338 3297
rect 21022 3232 21028 3296
rect 21092 3232 21108 3296
rect 21172 3232 21188 3296
rect 21252 3232 21268 3296
rect 21332 3232 21338 3296
rect 21022 3231 21338 3232
rect 27714 3296 28030 3297
rect 27714 3232 27720 3296
rect 27784 3232 27800 3296
rect 27864 3232 27880 3296
rect 27944 3232 27960 3296
rect 28024 3232 28030 3296
rect 27714 3231 28030 3232
rect 4292 2752 4608 2753
rect 4292 2688 4298 2752
rect 4362 2688 4378 2752
rect 4442 2688 4458 2752
rect 4522 2688 4538 2752
rect 4602 2688 4608 2752
rect 4292 2687 4608 2688
rect 10984 2752 11300 2753
rect 10984 2688 10990 2752
rect 11054 2688 11070 2752
rect 11134 2688 11150 2752
rect 11214 2688 11230 2752
rect 11294 2688 11300 2752
rect 10984 2687 11300 2688
rect 17676 2752 17992 2753
rect 17676 2688 17682 2752
rect 17746 2688 17762 2752
rect 17826 2688 17842 2752
rect 17906 2688 17922 2752
rect 17986 2688 17992 2752
rect 17676 2687 17992 2688
rect 24368 2752 24684 2753
rect 24368 2688 24374 2752
rect 24438 2688 24454 2752
rect 24518 2688 24534 2752
rect 24598 2688 24614 2752
rect 24678 2688 24684 2752
rect 24368 2687 24684 2688
rect 7638 2208 7954 2209
rect 0 2138 800 2168
rect 7638 2144 7644 2208
rect 7708 2144 7724 2208
rect 7788 2144 7804 2208
rect 7868 2144 7884 2208
rect 7948 2144 7954 2208
rect 7638 2143 7954 2144
rect 14330 2208 14646 2209
rect 14330 2144 14336 2208
rect 14400 2144 14416 2208
rect 14480 2144 14496 2208
rect 14560 2144 14576 2208
rect 14640 2144 14646 2208
rect 14330 2143 14646 2144
rect 21022 2208 21338 2209
rect 21022 2144 21028 2208
rect 21092 2144 21108 2208
rect 21172 2144 21188 2208
rect 21252 2144 21268 2208
rect 21332 2144 21338 2208
rect 21022 2143 21338 2144
rect 27714 2208 28030 2209
rect 27714 2144 27720 2208
rect 27784 2144 27800 2208
rect 27864 2144 27880 2208
rect 27944 2144 27960 2208
rect 28024 2144 28030 2208
rect 27714 2143 28030 2144
rect 3233 2138 3299 2141
rect 0 2136 3299 2138
rect 0 2080 3238 2136
rect 3294 2080 3299 2136
rect 0 2078 3299 2080
rect 0 2048 800 2078
rect 3233 2075 3299 2078
<< via3 >>
rect 4298 26684 4362 26688
rect 4298 26628 4302 26684
rect 4302 26628 4358 26684
rect 4358 26628 4362 26684
rect 4298 26624 4362 26628
rect 4378 26684 4442 26688
rect 4378 26628 4382 26684
rect 4382 26628 4438 26684
rect 4438 26628 4442 26684
rect 4378 26624 4442 26628
rect 4458 26684 4522 26688
rect 4458 26628 4462 26684
rect 4462 26628 4518 26684
rect 4518 26628 4522 26684
rect 4458 26624 4522 26628
rect 4538 26684 4602 26688
rect 4538 26628 4542 26684
rect 4542 26628 4598 26684
rect 4598 26628 4602 26684
rect 4538 26624 4602 26628
rect 10990 26684 11054 26688
rect 10990 26628 10994 26684
rect 10994 26628 11050 26684
rect 11050 26628 11054 26684
rect 10990 26624 11054 26628
rect 11070 26684 11134 26688
rect 11070 26628 11074 26684
rect 11074 26628 11130 26684
rect 11130 26628 11134 26684
rect 11070 26624 11134 26628
rect 11150 26684 11214 26688
rect 11150 26628 11154 26684
rect 11154 26628 11210 26684
rect 11210 26628 11214 26684
rect 11150 26624 11214 26628
rect 11230 26684 11294 26688
rect 11230 26628 11234 26684
rect 11234 26628 11290 26684
rect 11290 26628 11294 26684
rect 11230 26624 11294 26628
rect 17682 26684 17746 26688
rect 17682 26628 17686 26684
rect 17686 26628 17742 26684
rect 17742 26628 17746 26684
rect 17682 26624 17746 26628
rect 17762 26684 17826 26688
rect 17762 26628 17766 26684
rect 17766 26628 17822 26684
rect 17822 26628 17826 26684
rect 17762 26624 17826 26628
rect 17842 26684 17906 26688
rect 17842 26628 17846 26684
rect 17846 26628 17902 26684
rect 17902 26628 17906 26684
rect 17842 26624 17906 26628
rect 17922 26684 17986 26688
rect 17922 26628 17926 26684
rect 17926 26628 17982 26684
rect 17982 26628 17986 26684
rect 17922 26624 17986 26628
rect 24374 26684 24438 26688
rect 24374 26628 24378 26684
rect 24378 26628 24434 26684
rect 24434 26628 24438 26684
rect 24374 26624 24438 26628
rect 24454 26684 24518 26688
rect 24454 26628 24458 26684
rect 24458 26628 24514 26684
rect 24514 26628 24518 26684
rect 24454 26624 24518 26628
rect 24534 26684 24598 26688
rect 24534 26628 24538 26684
rect 24538 26628 24594 26684
rect 24594 26628 24598 26684
rect 24534 26624 24598 26628
rect 24614 26684 24678 26688
rect 24614 26628 24618 26684
rect 24618 26628 24674 26684
rect 24674 26628 24678 26684
rect 24614 26624 24678 26628
rect 7644 26140 7708 26144
rect 7644 26084 7648 26140
rect 7648 26084 7704 26140
rect 7704 26084 7708 26140
rect 7644 26080 7708 26084
rect 7724 26140 7788 26144
rect 7724 26084 7728 26140
rect 7728 26084 7784 26140
rect 7784 26084 7788 26140
rect 7724 26080 7788 26084
rect 7804 26140 7868 26144
rect 7804 26084 7808 26140
rect 7808 26084 7864 26140
rect 7864 26084 7868 26140
rect 7804 26080 7868 26084
rect 7884 26140 7948 26144
rect 7884 26084 7888 26140
rect 7888 26084 7944 26140
rect 7944 26084 7948 26140
rect 7884 26080 7948 26084
rect 14336 26140 14400 26144
rect 14336 26084 14340 26140
rect 14340 26084 14396 26140
rect 14396 26084 14400 26140
rect 14336 26080 14400 26084
rect 14416 26140 14480 26144
rect 14416 26084 14420 26140
rect 14420 26084 14476 26140
rect 14476 26084 14480 26140
rect 14416 26080 14480 26084
rect 14496 26140 14560 26144
rect 14496 26084 14500 26140
rect 14500 26084 14556 26140
rect 14556 26084 14560 26140
rect 14496 26080 14560 26084
rect 14576 26140 14640 26144
rect 14576 26084 14580 26140
rect 14580 26084 14636 26140
rect 14636 26084 14640 26140
rect 14576 26080 14640 26084
rect 21028 26140 21092 26144
rect 21028 26084 21032 26140
rect 21032 26084 21088 26140
rect 21088 26084 21092 26140
rect 21028 26080 21092 26084
rect 21108 26140 21172 26144
rect 21108 26084 21112 26140
rect 21112 26084 21168 26140
rect 21168 26084 21172 26140
rect 21108 26080 21172 26084
rect 21188 26140 21252 26144
rect 21188 26084 21192 26140
rect 21192 26084 21248 26140
rect 21248 26084 21252 26140
rect 21188 26080 21252 26084
rect 21268 26140 21332 26144
rect 21268 26084 21272 26140
rect 21272 26084 21328 26140
rect 21328 26084 21332 26140
rect 21268 26080 21332 26084
rect 27720 26140 27784 26144
rect 27720 26084 27724 26140
rect 27724 26084 27780 26140
rect 27780 26084 27784 26140
rect 27720 26080 27784 26084
rect 27800 26140 27864 26144
rect 27800 26084 27804 26140
rect 27804 26084 27860 26140
rect 27860 26084 27864 26140
rect 27800 26080 27864 26084
rect 27880 26140 27944 26144
rect 27880 26084 27884 26140
rect 27884 26084 27940 26140
rect 27940 26084 27944 26140
rect 27880 26080 27944 26084
rect 27960 26140 28024 26144
rect 27960 26084 27964 26140
rect 27964 26084 28020 26140
rect 28020 26084 28024 26140
rect 27960 26080 28024 26084
rect 4298 25596 4362 25600
rect 4298 25540 4302 25596
rect 4302 25540 4358 25596
rect 4358 25540 4362 25596
rect 4298 25536 4362 25540
rect 4378 25596 4442 25600
rect 4378 25540 4382 25596
rect 4382 25540 4438 25596
rect 4438 25540 4442 25596
rect 4378 25536 4442 25540
rect 4458 25596 4522 25600
rect 4458 25540 4462 25596
rect 4462 25540 4518 25596
rect 4518 25540 4522 25596
rect 4458 25536 4522 25540
rect 4538 25596 4602 25600
rect 4538 25540 4542 25596
rect 4542 25540 4598 25596
rect 4598 25540 4602 25596
rect 4538 25536 4602 25540
rect 10990 25596 11054 25600
rect 10990 25540 10994 25596
rect 10994 25540 11050 25596
rect 11050 25540 11054 25596
rect 10990 25536 11054 25540
rect 11070 25596 11134 25600
rect 11070 25540 11074 25596
rect 11074 25540 11130 25596
rect 11130 25540 11134 25596
rect 11070 25536 11134 25540
rect 11150 25596 11214 25600
rect 11150 25540 11154 25596
rect 11154 25540 11210 25596
rect 11210 25540 11214 25596
rect 11150 25536 11214 25540
rect 11230 25596 11294 25600
rect 11230 25540 11234 25596
rect 11234 25540 11290 25596
rect 11290 25540 11294 25596
rect 11230 25536 11294 25540
rect 17682 25596 17746 25600
rect 17682 25540 17686 25596
rect 17686 25540 17742 25596
rect 17742 25540 17746 25596
rect 17682 25536 17746 25540
rect 17762 25596 17826 25600
rect 17762 25540 17766 25596
rect 17766 25540 17822 25596
rect 17822 25540 17826 25596
rect 17762 25536 17826 25540
rect 17842 25596 17906 25600
rect 17842 25540 17846 25596
rect 17846 25540 17902 25596
rect 17902 25540 17906 25596
rect 17842 25536 17906 25540
rect 17922 25596 17986 25600
rect 17922 25540 17926 25596
rect 17926 25540 17982 25596
rect 17982 25540 17986 25596
rect 17922 25536 17986 25540
rect 24374 25596 24438 25600
rect 24374 25540 24378 25596
rect 24378 25540 24434 25596
rect 24434 25540 24438 25596
rect 24374 25536 24438 25540
rect 24454 25596 24518 25600
rect 24454 25540 24458 25596
rect 24458 25540 24514 25596
rect 24514 25540 24518 25596
rect 24454 25536 24518 25540
rect 24534 25596 24598 25600
rect 24534 25540 24538 25596
rect 24538 25540 24594 25596
rect 24594 25540 24598 25596
rect 24534 25536 24598 25540
rect 24614 25596 24678 25600
rect 24614 25540 24618 25596
rect 24618 25540 24674 25596
rect 24674 25540 24678 25596
rect 24614 25536 24678 25540
rect 7644 25052 7708 25056
rect 7644 24996 7648 25052
rect 7648 24996 7704 25052
rect 7704 24996 7708 25052
rect 7644 24992 7708 24996
rect 7724 25052 7788 25056
rect 7724 24996 7728 25052
rect 7728 24996 7784 25052
rect 7784 24996 7788 25052
rect 7724 24992 7788 24996
rect 7804 25052 7868 25056
rect 7804 24996 7808 25052
rect 7808 24996 7864 25052
rect 7864 24996 7868 25052
rect 7804 24992 7868 24996
rect 7884 25052 7948 25056
rect 7884 24996 7888 25052
rect 7888 24996 7944 25052
rect 7944 24996 7948 25052
rect 7884 24992 7948 24996
rect 14336 25052 14400 25056
rect 14336 24996 14340 25052
rect 14340 24996 14396 25052
rect 14396 24996 14400 25052
rect 14336 24992 14400 24996
rect 14416 25052 14480 25056
rect 14416 24996 14420 25052
rect 14420 24996 14476 25052
rect 14476 24996 14480 25052
rect 14416 24992 14480 24996
rect 14496 25052 14560 25056
rect 14496 24996 14500 25052
rect 14500 24996 14556 25052
rect 14556 24996 14560 25052
rect 14496 24992 14560 24996
rect 14576 25052 14640 25056
rect 14576 24996 14580 25052
rect 14580 24996 14636 25052
rect 14636 24996 14640 25052
rect 14576 24992 14640 24996
rect 21028 25052 21092 25056
rect 21028 24996 21032 25052
rect 21032 24996 21088 25052
rect 21088 24996 21092 25052
rect 21028 24992 21092 24996
rect 21108 25052 21172 25056
rect 21108 24996 21112 25052
rect 21112 24996 21168 25052
rect 21168 24996 21172 25052
rect 21108 24992 21172 24996
rect 21188 25052 21252 25056
rect 21188 24996 21192 25052
rect 21192 24996 21248 25052
rect 21248 24996 21252 25052
rect 21188 24992 21252 24996
rect 21268 25052 21332 25056
rect 21268 24996 21272 25052
rect 21272 24996 21328 25052
rect 21328 24996 21332 25052
rect 21268 24992 21332 24996
rect 27720 25052 27784 25056
rect 27720 24996 27724 25052
rect 27724 24996 27780 25052
rect 27780 24996 27784 25052
rect 27720 24992 27784 24996
rect 27800 25052 27864 25056
rect 27800 24996 27804 25052
rect 27804 24996 27860 25052
rect 27860 24996 27864 25052
rect 27800 24992 27864 24996
rect 27880 25052 27944 25056
rect 27880 24996 27884 25052
rect 27884 24996 27940 25052
rect 27940 24996 27944 25052
rect 27880 24992 27944 24996
rect 27960 25052 28024 25056
rect 27960 24996 27964 25052
rect 27964 24996 28020 25052
rect 28020 24996 28024 25052
rect 27960 24992 28024 24996
rect 4298 24508 4362 24512
rect 4298 24452 4302 24508
rect 4302 24452 4358 24508
rect 4358 24452 4362 24508
rect 4298 24448 4362 24452
rect 4378 24508 4442 24512
rect 4378 24452 4382 24508
rect 4382 24452 4438 24508
rect 4438 24452 4442 24508
rect 4378 24448 4442 24452
rect 4458 24508 4522 24512
rect 4458 24452 4462 24508
rect 4462 24452 4518 24508
rect 4518 24452 4522 24508
rect 4458 24448 4522 24452
rect 4538 24508 4602 24512
rect 4538 24452 4542 24508
rect 4542 24452 4598 24508
rect 4598 24452 4602 24508
rect 4538 24448 4602 24452
rect 10990 24508 11054 24512
rect 10990 24452 10994 24508
rect 10994 24452 11050 24508
rect 11050 24452 11054 24508
rect 10990 24448 11054 24452
rect 11070 24508 11134 24512
rect 11070 24452 11074 24508
rect 11074 24452 11130 24508
rect 11130 24452 11134 24508
rect 11070 24448 11134 24452
rect 11150 24508 11214 24512
rect 11150 24452 11154 24508
rect 11154 24452 11210 24508
rect 11210 24452 11214 24508
rect 11150 24448 11214 24452
rect 11230 24508 11294 24512
rect 11230 24452 11234 24508
rect 11234 24452 11290 24508
rect 11290 24452 11294 24508
rect 11230 24448 11294 24452
rect 17682 24508 17746 24512
rect 17682 24452 17686 24508
rect 17686 24452 17742 24508
rect 17742 24452 17746 24508
rect 17682 24448 17746 24452
rect 17762 24508 17826 24512
rect 17762 24452 17766 24508
rect 17766 24452 17822 24508
rect 17822 24452 17826 24508
rect 17762 24448 17826 24452
rect 17842 24508 17906 24512
rect 17842 24452 17846 24508
rect 17846 24452 17902 24508
rect 17902 24452 17906 24508
rect 17842 24448 17906 24452
rect 17922 24508 17986 24512
rect 17922 24452 17926 24508
rect 17926 24452 17982 24508
rect 17982 24452 17986 24508
rect 17922 24448 17986 24452
rect 24374 24508 24438 24512
rect 24374 24452 24378 24508
rect 24378 24452 24434 24508
rect 24434 24452 24438 24508
rect 24374 24448 24438 24452
rect 24454 24508 24518 24512
rect 24454 24452 24458 24508
rect 24458 24452 24514 24508
rect 24514 24452 24518 24508
rect 24454 24448 24518 24452
rect 24534 24508 24598 24512
rect 24534 24452 24538 24508
rect 24538 24452 24594 24508
rect 24594 24452 24598 24508
rect 24534 24448 24598 24452
rect 24614 24508 24678 24512
rect 24614 24452 24618 24508
rect 24618 24452 24674 24508
rect 24674 24452 24678 24508
rect 24614 24448 24678 24452
rect 7644 23964 7708 23968
rect 7644 23908 7648 23964
rect 7648 23908 7704 23964
rect 7704 23908 7708 23964
rect 7644 23904 7708 23908
rect 7724 23964 7788 23968
rect 7724 23908 7728 23964
rect 7728 23908 7784 23964
rect 7784 23908 7788 23964
rect 7724 23904 7788 23908
rect 7804 23964 7868 23968
rect 7804 23908 7808 23964
rect 7808 23908 7864 23964
rect 7864 23908 7868 23964
rect 7804 23904 7868 23908
rect 7884 23964 7948 23968
rect 7884 23908 7888 23964
rect 7888 23908 7944 23964
rect 7944 23908 7948 23964
rect 7884 23904 7948 23908
rect 14336 23964 14400 23968
rect 14336 23908 14340 23964
rect 14340 23908 14396 23964
rect 14396 23908 14400 23964
rect 14336 23904 14400 23908
rect 14416 23964 14480 23968
rect 14416 23908 14420 23964
rect 14420 23908 14476 23964
rect 14476 23908 14480 23964
rect 14416 23904 14480 23908
rect 14496 23964 14560 23968
rect 14496 23908 14500 23964
rect 14500 23908 14556 23964
rect 14556 23908 14560 23964
rect 14496 23904 14560 23908
rect 14576 23964 14640 23968
rect 14576 23908 14580 23964
rect 14580 23908 14636 23964
rect 14636 23908 14640 23964
rect 14576 23904 14640 23908
rect 21028 23964 21092 23968
rect 21028 23908 21032 23964
rect 21032 23908 21088 23964
rect 21088 23908 21092 23964
rect 21028 23904 21092 23908
rect 21108 23964 21172 23968
rect 21108 23908 21112 23964
rect 21112 23908 21168 23964
rect 21168 23908 21172 23964
rect 21108 23904 21172 23908
rect 21188 23964 21252 23968
rect 21188 23908 21192 23964
rect 21192 23908 21248 23964
rect 21248 23908 21252 23964
rect 21188 23904 21252 23908
rect 21268 23964 21332 23968
rect 21268 23908 21272 23964
rect 21272 23908 21328 23964
rect 21328 23908 21332 23964
rect 21268 23904 21332 23908
rect 27720 23964 27784 23968
rect 27720 23908 27724 23964
rect 27724 23908 27780 23964
rect 27780 23908 27784 23964
rect 27720 23904 27784 23908
rect 27800 23964 27864 23968
rect 27800 23908 27804 23964
rect 27804 23908 27860 23964
rect 27860 23908 27864 23964
rect 27800 23904 27864 23908
rect 27880 23964 27944 23968
rect 27880 23908 27884 23964
rect 27884 23908 27940 23964
rect 27940 23908 27944 23964
rect 27880 23904 27944 23908
rect 27960 23964 28024 23968
rect 27960 23908 27964 23964
rect 27964 23908 28020 23964
rect 28020 23908 28024 23964
rect 27960 23904 28024 23908
rect 4298 23420 4362 23424
rect 4298 23364 4302 23420
rect 4302 23364 4358 23420
rect 4358 23364 4362 23420
rect 4298 23360 4362 23364
rect 4378 23420 4442 23424
rect 4378 23364 4382 23420
rect 4382 23364 4438 23420
rect 4438 23364 4442 23420
rect 4378 23360 4442 23364
rect 4458 23420 4522 23424
rect 4458 23364 4462 23420
rect 4462 23364 4518 23420
rect 4518 23364 4522 23420
rect 4458 23360 4522 23364
rect 4538 23420 4602 23424
rect 4538 23364 4542 23420
rect 4542 23364 4598 23420
rect 4598 23364 4602 23420
rect 4538 23360 4602 23364
rect 10990 23420 11054 23424
rect 10990 23364 10994 23420
rect 10994 23364 11050 23420
rect 11050 23364 11054 23420
rect 10990 23360 11054 23364
rect 11070 23420 11134 23424
rect 11070 23364 11074 23420
rect 11074 23364 11130 23420
rect 11130 23364 11134 23420
rect 11070 23360 11134 23364
rect 11150 23420 11214 23424
rect 11150 23364 11154 23420
rect 11154 23364 11210 23420
rect 11210 23364 11214 23420
rect 11150 23360 11214 23364
rect 11230 23420 11294 23424
rect 11230 23364 11234 23420
rect 11234 23364 11290 23420
rect 11290 23364 11294 23420
rect 11230 23360 11294 23364
rect 17682 23420 17746 23424
rect 17682 23364 17686 23420
rect 17686 23364 17742 23420
rect 17742 23364 17746 23420
rect 17682 23360 17746 23364
rect 17762 23420 17826 23424
rect 17762 23364 17766 23420
rect 17766 23364 17822 23420
rect 17822 23364 17826 23420
rect 17762 23360 17826 23364
rect 17842 23420 17906 23424
rect 17842 23364 17846 23420
rect 17846 23364 17902 23420
rect 17902 23364 17906 23420
rect 17842 23360 17906 23364
rect 17922 23420 17986 23424
rect 17922 23364 17926 23420
rect 17926 23364 17982 23420
rect 17982 23364 17986 23420
rect 17922 23360 17986 23364
rect 24374 23420 24438 23424
rect 24374 23364 24378 23420
rect 24378 23364 24434 23420
rect 24434 23364 24438 23420
rect 24374 23360 24438 23364
rect 24454 23420 24518 23424
rect 24454 23364 24458 23420
rect 24458 23364 24514 23420
rect 24514 23364 24518 23420
rect 24454 23360 24518 23364
rect 24534 23420 24598 23424
rect 24534 23364 24538 23420
rect 24538 23364 24594 23420
rect 24594 23364 24598 23420
rect 24534 23360 24598 23364
rect 24614 23420 24678 23424
rect 24614 23364 24618 23420
rect 24618 23364 24674 23420
rect 24674 23364 24678 23420
rect 24614 23360 24678 23364
rect 7644 22876 7708 22880
rect 7644 22820 7648 22876
rect 7648 22820 7704 22876
rect 7704 22820 7708 22876
rect 7644 22816 7708 22820
rect 7724 22876 7788 22880
rect 7724 22820 7728 22876
rect 7728 22820 7784 22876
rect 7784 22820 7788 22876
rect 7724 22816 7788 22820
rect 7804 22876 7868 22880
rect 7804 22820 7808 22876
rect 7808 22820 7864 22876
rect 7864 22820 7868 22876
rect 7804 22816 7868 22820
rect 7884 22876 7948 22880
rect 7884 22820 7888 22876
rect 7888 22820 7944 22876
rect 7944 22820 7948 22876
rect 7884 22816 7948 22820
rect 14336 22876 14400 22880
rect 14336 22820 14340 22876
rect 14340 22820 14396 22876
rect 14396 22820 14400 22876
rect 14336 22816 14400 22820
rect 14416 22876 14480 22880
rect 14416 22820 14420 22876
rect 14420 22820 14476 22876
rect 14476 22820 14480 22876
rect 14416 22816 14480 22820
rect 14496 22876 14560 22880
rect 14496 22820 14500 22876
rect 14500 22820 14556 22876
rect 14556 22820 14560 22876
rect 14496 22816 14560 22820
rect 14576 22876 14640 22880
rect 14576 22820 14580 22876
rect 14580 22820 14636 22876
rect 14636 22820 14640 22876
rect 14576 22816 14640 22820
rect 21028 22876 21092 22880
rect 21028 22820 21032 22876
rect 21032 22820 21088 22876
rect 21088 22820 21092 22876
rect 21028 22816 21092 22820
rect 21108 22876 21172 22880
rect 21108 22820 21112 22876
rect 21112 22820 21168 22876
rect 21168 22820 21172 22876
rect 21108 22816 21172 22820
rect 21188 22876 21252 22880
rect 21188 22820 21192 22876
rect 21192 22820 21248 22876
rect 21248 22820 21252 22876
rect 21188 22816 21252 22820
rect 21268 22876 21332 22880
rect 21268 22820 21272 22876
rect 21272 22820 21328 22876
rect 21328 22820 21332 22876
rect 21268 22816 21332 22820
rect 27720 22876 27784 22880
rect 27720 22820 27724 22876
rect 27724 22820 27780 22876
rect 27780 22820 27784 22876
rect 27720 22816 27784 22820
rect 27800 22876 27864 22880
rect 27800 22820 27804 22876
rect 27804 22820 27860 22876
rect 27860 22820 27864 22876
rect 27800 22816 27864 22820
rect 27880 22876 27944 22880
rect 27880 22820 27884 22876
rect 27884 22820 27940 22876
rect 27940 22820 27944 22876
rect 27880 22816 27944 22820
rect 27960 22876 28024 22880
rect 27960 22820 27964 22876
rect 27964 22820 28020 22876
rect 28020 22820 28024 22876
rect 27960 22816 28024 22820
rect 4298 22332 4362 22336
rect 4298 22276 4302 22332
rect 4302 22276 4358 22332
rect 4358 22276 4362 22332
rect 4298 22272 4362 22276
rect 4378 22332 4442 22336
rect 4378 22276 4382 22332
rect 4382 22276 4438 22332
rect 4438 22276 4442 22332
rect 4378 22272 4442 22276
rect 4458 22332 4522 22336
rect 4458 22276 4462 22332
rect 4462 22276 4518 22332
rect 4518 22276 4522 22332
rect 4458 22272 4522 22276
rect 4538 22332 4602 22336
rect 4538 22276 4542 22332
rect 4542 22276 4598 22332
rect 4598 22276 4602 22332
rect 4538 22272 4602 22276
rect 10990 22332 11054 22336
rect 10990 22276 10994 22332
rect 10994 22276 11050 22332
rect 11050 22276 11054 22332
rect 10990 22272 11054 22276
rect 11070 22332 11134 22336
rect 11070 22276 11074 22332
rect 11074 22276 11130 22332
rect 11130 22276 11134 22332
rect 11070 22272 11134 22276
rect 11150 22332 11214 22336
rect 11150 22276 11154 22332
rect 11154 22276 11210 22332
rect 11210 22276 11214 22332
rect 11150 22272 11214 22276
rect 11230 22332 11294 22336
rect 11230 22276 11234 22332
rect 11234 22276 11290 22332
rect 11290 22276 11294 22332
rect 11230 22272 11294 22276
rect 17682 22332 17746 22336
rect 17682 22276 17686 22332
rect 17686 22276 17742 22332
rect 17742 22276 17746 22332
rect 17682 22272 17746 22276
rect 17762 22332 17826 22336
rect 17762 22276 17766 22332
rect 17766 22276 17822 22332
rect 17822 22276 17826 22332
rect 17762 22272 17826 22276
rect 17842 22332 17906 22336
rect 17842 22276 17846 22332
rect 17846 22276 17902 22332
rect 17902 22276 17906 22332
rect 17842 22272 17906 22276
rect 17922 22332 17986 22336
rect 17922 22276 17926 22332
rect 17926 22276 17982 22332
rect 17982 22276 17986 22332
rect 17922 22272 17986 22276
rect 24374 22332 24438 22336
rect 24374 22276 24378 22332
rect 24378 22276 24434 22332
rect 24434 22276 24438 22332
rect 24374 22272 24438 22276
rect 24454 22332 24518 22336
rect 24454 22276 24458 22332
rect 24458 22276 24514 22332
rect 24514 22276 24518 22332
rect 24454 22272 24518 22276
rect 24534 22332 24598 22336
rect 24534 22276 24538 22332
rect 24538 22276 24594 22332
rect 24594 22276 24598 22332
rect 24534 22272 24598 22276
rect 24614 22332 24678 22336
rect 24614 22276 24618 22332
rect 24618 22276 24674 22332
rect 24674 22276 24678 22332
rect 24614 22272 24678 22276
rect 7644 21788 7708 21792
rect 7644 21732 7648 21788
rect 7648 21732 7704 21788
rect 7704 21732 7708 21788
rect 7644 21728 7708 21732
rect 7724 21788 7788 21792
rect 7724 21732 7728 21788
rect 7728 21732 7784 21788
rect 7784 21732 7788 21788
rect 7724 21728 7788 21732
rect 7804 21788 7868 21792
rect 7804 21732 7808 21788
rect 7808 21732 7864 21788
rect 7864 21732 7868 21788
rect 7804 21728 7868 21732
rect 7884 21788 7948 21792
rect 7884 21732 7888 21788
rect 7888 21732 7944 21788
rect 7944 21732 7948 21788
rect 7884 21728 7948 21732
rect 14336 21788 14400 21792
rect 14336 21732 14340 21788
rect 14340 21732 14396 21788
rect 14396 21732 14400 21788
rect 14336 21728 14400 21732
rect 14416 21788 14480 21792
rect 14416 21732 14420 21788
rect 14420 21732 14476 21788
rect 14476 21732 14480 21788
rect 14416 21728 14480 21732
rect 14496 21788 14560 21792
rect 14496 21732 14500 21788
rect 14500 21732 14556 21788
rect 14556 21732 14560 21788
rect 14496 21728 14560 21732
rect 14576 21788 14640 21792
rect 14576 21732 14580 21788
rect 14580 21732 14636 21788
rect 14636 21732 14640 21788
rect 14576 21728 14640 21732
rect 21028 21788 21092 21792
rect 21028 21732 21032 21788
rect 21032 21732 21088 21788
rect 21088 21732 21092 21788
rect 21028 21728 21092 21732
rect 21108 21788 21172 21792
rect 21108 21732 21112 21788
rect 21112 21732 21168 21788
rect 21168 21732 21172 21788
rect 21108 21728 21172 21732
rect 21188 21788 21252 21792
rect 21188 21732 21192 21788
rect 21192 21732 21248 21788
rect 21248 21732 21252 21788
rect 21188 21728 21252 21732
rect 21268 21788 21332 21792
rect 21268 21732 21272 21788
rect 21272 21732 21328 21788
rect 21328 21732 21332 21788
rect 21268 21728 21332 21732
rect 27720 21788 27784 21792
rect 27720 21732 27724 21788
rect 27724 21732 27780 21788
rect 27780 21732 27784 21788
rect 27720 21728 27784 21732
rect 27800 21788 27864 21792
rect 27800 21732 27804 21788
rect 27804 21732 27860 21788
rect 27860 21732 27864 21788
rect 27800 21728 27864 21732
rect 27880 21788 27944 21792
rect 27880 21732 27884 21788
rect 27884 21732 27940 21788
rect 27940 21732 27944 21788
rect 27880 21728 27944 21732
rect 27960 21788 28024 21792
rect 27960 21732 27964 21788
rect 27964 21732 28020 21788
rect 28020 21732 28024 21788
rect 27960 21728 28024 21732
rect 4298 21244 4362 21248
rect 4298 21188 4302 21244
rect 4302 21188 4358 21244
rect 4358 21188 4362 21244
rect 4298 21184 4362 21188
rect 4378 21244 4442 21248
rect 4378 21188 4382 21244
rect 4382 21188 4438 21244
rect 4438 21188 4442 21244
rect 4378 21184 4442 21188
rect 4458 21244 4522 21248
rect 4458 21188 4462 21244
rect 4462 21188 4518 21244
rect 4518 21188 4522 21244
rect 4458 21184 4522 21188
rect 4538 21244 4602 21248
rect 4538 21188 4542 21244
rect 4542 21188 4598 21244
rect 4598 21188 4602 21244
rect 4538 21184 4602 21188
rect 10990 21244 11054 21248
rect 10990 21188 10994 21244
rect 10994 21188 11050 21244
rect 11050 21188 11054 21244
rect 10990 21184 11054 21188
rect 11070 21244 11134 21248
rect 11070 21188 11074 21244
rect 11074 21188 11130 21244
rect 11130 21188 11134 21244
rect 11070 21184 11134 21188
rect 11150 21244 11214 21248
rect 11150 21188 11154 21244
rect 11154 21188 11210 21244
rect 11210 21188 11214 21244
rect 11150 21184 11214 21188
rect 11230 21244 11294 21248
rect 11230 21188 11234 21244
rect 11234 21188 11290 21244
rect 11290 21188 11294 21244
rect 11230 21184 11294 21188
rect 17682 21244 17746 21248
rect 17682 21188 17686 21244
rect 17686 21188 17742 21244
rect 17742 21188 17746 21244
rect 17682 21184 17746 21188
rect 17762 21244 17826 21248
rect 17762 21188 17766 21244
rect 17766 21188 17822 21244
rect 17822 21188 17826 21244
rect 17762 21184 17826 21188
rect 17842 21244 17906 21248
rect 17842 21188 17846 21244
rect 17846 21188 17902 21244
rect 17902 21188 17906 21244
rect 17842 21184 17906 21188
rect 17922 21244 17986 21248
rect 17922 21188 17926 21244
rect 17926 21188 17982 21244
rect 17982 21188 17986 21244
rect 17922 21184 17986 21188
rect 24374 21244 24438 21248
rect 24374 21188 24378 21244
rect 24378 21188 24434 21244
rect 24434 21188 24438 21244
rect 24374 21184 24438 21188
rect 24454 21244 24518 21248
rect 24454 21188 24458 21244
rect 24458 21188 24514 21244
rect 24514 21188 24518 21244
rect 24454 21184 24518 21188
rect 24534 21244 24598 21248
rect 24534 21188 24538 21244
rect 24538 21188 24594 21244
rect 24594 21188 24598 21244
rect 24534 21184 24598 21188
rect 24614 21244 24678 21248
rect 24614 21188 24618 21244
rect 24618 21188 24674 21244
rect 24674 21188 24678 21244
rect 24614 21184 24678 21188
rect 7644 20700 7708 20704
rect 7644 20644 7648 20700
rect 7648 20644 7704 20700
rect 7704 20644 7708 20700
rect 7644 20640 7708 20644
rect 7724 20700 7788 20704
rect 7724 20644 7728 20700
rect 7728 20644 7784 20700
rect 7784 20644 7788 20700
rect 7724 20640 7788 20644
rect 7804 20700 7868 20704
rect 7804 20644 7808 20700
rect 7808 20644 7864 20700
rect 7864 20644 7868 20700
rect 7804 20640 7868 20644
rect 7884 20700 7948 20704
rect 7884 20644 7888 20700
rect 7888 20644 7944 20700
rect 7944 20644 7948 20700
rect 7884 20640 7948 20644
rect 14336 20700 14400 20704
rect 14336 20644 14340 20700
rect 14340 20644 14396 20700
rect 14396 20644 14400 20700
rect 14336 20640 14400 20644
rect 14416 20700 14480 20704
rect 14416 20644 14420 20700
rect 14420 20644 14476 20700
rect 14476 20644 14480 20700
rect 14416 20640 14480 20644
rect 14496 20700 14560 20704
rect 14496 20644 14500 20700
rect 14500 20644 14556 20700
rect 14556 20644 14560 20700
rect 14496 20640 14560 20644
rect 14576 20700 14640 20704
rect 14576 20644 14580 20700
rect 14580 20644 14636 20700
rect 14636 20644 14640 20700
rect 14576 20640 14640 20644
rect 21028 20700 21092 20704
rect 21028 20644 21032 20700
rect 21032 20644 21088 20700
rect 21088 20644 21092 20700
rect 21028 20640 21092 20644
rect 21108 20700 21172 20704
rect 21108 20644 21112 20700
rect 21112 20644 21168 20700
rect 21168 20644 21172 20700
rect 21108 20640 21172 20644
rect 21188 20700 21252 20704
rect 21188 20644 21192 20700
rect 21192 20644 21248 20700
rect 21248 20644 21252 20700
rect 21188 20640 21252 20644
rect 21268 20700 21332 20704
rect 21268 20644 21272 20700
rect 21272 20644 21328 20700
rect 21328 20644 21332 20700
rect 21268 20640 21332 20644
rect 27720 20700 27784 20704
rect 27720 20644 27724 20700
rect 27724 20644 27780 20700
rect 27780 20644 27784 20700
rect 27720 20640 27784 20644
rect 27800 20700 27864 20704
rect 27800 20644 27804 20700
rect 27804 20644 27860 20700
rect 27860 20644 27864 20700
rect 27800 20640 27864 20644
rect 27880 20700 27944 20704
rect 27880 20644 27884 20700
rect 27884 20644 27940 20700
rect 27940 20644 27944 20700
rect 27880 20640 27944 20644
rect 27960 20700 28024 20704
rect 27960 20644 27964 20700
rect 27964 20644 28020 20700
rect 28020 20644 28024 20700
rect 27960 20640 28024 20644
rect 4298 20156 4362 20160
rect 4298 20100 4302 20156
rect 4302 20100 4358 20156
rect 4358 20100 4362 20156
rect 4298 20096 4362 20100
rect 4378 20156 4442 20160
rect 4378 20100 4382 20156
rect 4382 20100 4438 20156
rect 4438 20100 4442 20156
rect 4378 20096 4442 20100
rect 4458 20156 4522 20160
rect 4458 20100 4462 20156
rect 4462 20100 4518 20156
rect 4518 20100 4522 20156
rect 4458 20096 4522 20100
rect 4538 20156 4602 20160
rect 4538 20100 4542 20156
rect 4542 20100 4598 20156
rect 4598 20100 4602 20156
rect 4538 20096 4602 20100
rect 10990 20156 11054 20160
rect 10990 20100 10994 20156
rect 10994 20100 11050 20156
rect 11050 20100 11054 20156
rect 10990 20096 11054 20100
rect 11070 20156 11134 20160
rect 11070 20100 11074 20156
rect 11074 20100 11130 20156
rect 11130 20100 11134 20156
rect 11070 20096 11134 20100
rect 11150 20156 11214 20160
rect 11150 20100 11154 20156
rect 11154 20100 11210 20156
rect 11210 20100 11214 20156
rect 11150 20096 11214 20100
rect 11230 20156 11294 20160
rect 11230 20100 11234 20156
rect 11234 20100 11290 20156
rect 11290 20100 11294 20156
rect 11230 20096 11294 20100
rect 17682 20156 17746 20160
rect 17682 20100 17686 20156
rect 17686 20100 17742 20156
rect 17742 20100 17746 20156
rect 17682 20096 17746 20100
rect 17762 20156 17826 20160
rect 17762 20100 17766 20156
rect 17766 20100 17822 20156
rect 17822 20100 17826 20156
rect 17762 20096 17826 20100
rect 17842 20156 17906 20160
rect 17842 20100 17846 20156
rect 17846 20100 17902 20156
rect 17902 20100 17906 20156
rect 17842 20096 17906 20100
rect 17922 20156 17986 20160
rect 17922 20100 17926 20156
rect 17926 20100 17982 20156
rect 17982 20100 17986 20156
rect 17922 20096 17986 20100
rect 24374 20156 24438 20160
rect 24374 20100 24378 20156
rect 24378 20100 24434 20156
rect 24434 20100 24438 20156
rect 24374 20096 24438 20100
rect 24454 20156 24518 20160
rect 24454 20100 24458 20156
rect 24458 20100 24514 20156
rect 24514 20100 24518 20156
rect 24454 20096 24518 20100
rect 24534 20156 24598 20160
rect 24534 20100 24538 20156
rect 24538 20100 24594 20156
rect 24594 20100 24598 20156
rect 24534 20096 24598 20100
rect 24614 20156 24678 20160
rect 24614 20100 24618 20156
rect 24618 20100 24674 20156
rect 24674 20100 24678 20156
rect 24614 20096 24678 20100
rect 7644 19612 7708 19616
rect 7644 19556 7648 19612
rect 7648 19556 7704 19612
rect 7704 19556 7708 19612
rect 7644 19552 7708 19556
rect 7724 19612 7788 19616
rect 7724 19556 7728 19612
rect 7728 19556 7784 19612
rect 7784 19556 7788 19612
rect 7724 19552 7788 19556
rect 7804 19612 7868 19616
rect 7804 19556 7808 19612
rect 7808 19556 7864 19612
rect 7864 19556 7868 19612
rect 7804 19552 7868 19556
rect 7884 19612 7948 19616
rect 7884 19556 7888 19612
rect 7888 19556 7944 19612
rect 7944 19556 7948 19612
rect 7884 19552 7948 19556
rect 14336 19612 14400 19616
rect 14336 19556 14340 19612
rect 14340 19556 14396 19612
rect 14396 19556 14400 19612
rect 14336 19552 14400 19556
rect 14416 19612 14480 19616
rect 14416 19556 14420 19612
rect 14420 19556 14476 19612
rect 14476 19556 14480 19612
rect 14416 19552 14480 19556
rect 14496 19612 14560 19616
rect 14496 19556 14500 19612
rect 14500 19556 14556 19612
rect 14556 19556 14560 19612
rect 14496 19552 14560 19556
rect 14576 19612 14640 19616
rect 14576 19556 14580 19612
rect 14580 19556 14636 19612
rect 14636 19556 14640 19612
rect 14576 19552 14640 19556
rect 21028 19612 21092 19616
rect 21028 19556 21032 19612
rect 21032 19556 21088 19612
rect 21088 19556 21092 19612
rect 21028 19552 21092 19556
rect 21108 19612 21172 19616
rect 21108 19556 21112 19612
rect 21112 19556 21168 19612
rect 21168 19556 21172 19612
rect 21108 19552 21172 19556
rect 21188 19612 21252 19616
rect 21188 19556 21192 19612
rect 21192 19556 21248 19612
rect 21248 19556 21252 19612
rect 21188 19552 21252 19556
rect 21268 19612 21332 19616
rect 21268 19556 21272 19612
rect 21272 19556 21328 19612
rect 21328 19556 21332 19612
rect 21268 19552 21332 19556
rect 27720 19612 27784 19616
rect 27720 19556 27724 19612
rect 27724 19556 27780 19612
rect 27780 19556 27784 19612
rect 27720 19552 27784 19556
rect 27800 19612 27864 19616
rect 27800 19556 27804 19612
rect 27804 19556 27860 19612
rect 27860 19556 27864 19612
rect 27800 19552 27864 19556
rect 27880 19612 27944 19616
rect 27880 19556 27884 19612
rect 27884 19556 27940 19612
rect 27940 19556 27944 19612
rect 27880 19552 27944 19556
rect 27960 19612 28024 19616
rect 27960 19556 27964 19612
rect 27964 19556 28020 19612
rect 28020 19556 28024 19612
rect 27960 19552 28024 19556
rect 4298 19068 4362 19072
rect 4298 19012 4302 19068
rect 4302 19012 4358 19068
rect 4358 19012 4362 19068
rect 4298 19008 4362 19012
rect 4378 19068 4442 19072
rect 4378 19012 4382 19068
rect 4382 19012 4438 19068
rect 4438 19012 4442 19068
rect 4378 19008 4442 19012
rect 4458 19068 4522 19072
rect 4458 19012 4462 19068
rect 4462 19012 4518 19068
rect 4518 19012 4522 19068
rect 4458 19008 4522 19012
rect 4538 19068 4602 19072
rect 4538 19012 4542 19068
rect 4542 19012 4598 19068
rect 4598 19012 4602 19068
rect 4538 19008 4602 19012
rect 10990 19068 11054 19072
rect 10990 19012 10994 19068
rect 10994 19012 11050 19068
rect 11050 19012 11054 19068
rect 10990 19008 11054 19012
rect 11070 19068 11134 19072
rect 11070 19012 11074 19068
rect 11074 19012 11130 19068
rect 11130 19012 11134 19068
rect 11070 19008 11134 19012
rect 11150 19068 11214 19072
rect 11150 19012 11154 19068
rect 11154 19012 11210 19068
rect 11210 19012 11214 19068
rect 11150 19008 11214 19012
rect 11230 19068 11294 19072
rect 11230 19012 11234 19068
rect 11234 19012 11290 19068
rect 11290 19012 11294 19068
rect 11230 19008 11294 19012
rect 17682 19068 17746 19072
rect 17682 19012 17686 19068
rect 17686 19012 17742 19068
rect 17742 19012 17746 19068
rect 17682 19008 17746 19012
rect 17762 19068 17826 19072
rect 17762 19012 17766 19068
rect 17766 19012 17822 19068
rect 17822 19012 17826 19068
rect 17762 19008 17826 19012
rect 17842 19068 17906 19072
rect 17842 19012 17846 19068
rect 17846 19012 17902 19068
rect 17902 19012 17906 19068
rect 17842 19008 17906 19012
rect 17922 19068 17986 19072
rect 17922 19012 17926 19068
rect 17926 19012 17982 19068
rect 17982 19012 17986 19068
rect 17922 19008 17986 19012
rect 24374 19068 24438 19072
rect 24374 19012 24378 19068
rect 24378 19012 24434 19068
rect 24434 19012 24438 19068
rect 24374 19008 24438 19012
rect 24454 19068 24518 19072
rect 24454 19012 24458 19068
rect 24458 19012 24514 19068
rect 24514 19012 24518 19068
rect 24454 19008 24518 19012
rect 24534 19068 24598 19072
rect 24534 19012 24538 19068
rect 24538 19012 24594 19068
rect 24594 19012 24598 19068
rect 24534 19008 24598 19012
rect 24614 19068 24678 19072
rect 24614 19012 24618 19068
rect 24618 19012 24674 19068
rect 24674 19012 24678 19068
rect 24614 19008 24678 19012
rect 7644 18524 7708 18528
rect 7644 18468 7648 18524
rect 7648 18468 7704 18524
rect 7704 18468 7708 18524
rect 7644 18464 7708 18468
rect 7724 18524 7788 18528
rect 7724 18468 7728 18524
rect 7728 18468 7784 18524
rect 7784 18468 7788 18524
rect 7724 18464 7788 18468
rect 7804 18524 7868 18528
rect 7804 18468 7808 18524
rect 7808 18468 7864 18524
rect 7864 18468 7868 18524
rect 7804 18464 7868 18468
rect 7884 18524 7948 18528
rect 7884 18468 7888 18524
rect 7888 18468 7944 18524
rect 7944 18468 7948 18524
rect 7884 18464 7948 18468
rect 14336 18524 14400 18528
rect 14336 18468 14340 18524
rect 14340 18468 14396 18524
rect 14396 18468 14400 18524
rect 14336 18464 14400 18468
rect 14416 18524 14480 18528
rect 14416 18468 14420 18524
rect 14420 18468 14476 18524
rect 14476 18468 14480 18524
rect 14416 18464 14480 18468
rect 14496 18524 14560 18528
rect 14496 18468 14500 18524
rect 14500 18468 14556 18524
rect 14556 18468 14560 18524
rect 14496 18464 14560 18468
rect 14576 18524 14640 18528
rect 14576 18468 14580 18524
rect 14580 18468 14636 18524
rect 14636 18468 14640 18524
rect 14576 18464 14640 18468
rect 21028 18524 21092 18528
rect 21028 18468 21032 18524
rect 21032 18468 21088 18524
rect 21088 18468 21092 18524
rect 21028 18464 21092 18468
rect 21108 18524 21172 18528
rect 21108 18468 21112 18524
rect 21112 18468 21168 18524
rect 21168 18468 21172 18524
rect 21108 18464 21172 18468
rect 21188 18524 21252 18528
rect 21188 18468 21192 18524
rect 21192 18468 21248 18524
rect 21248 18468 21252 18524
rect 21188 18464 21252 18468
rect 21268 18524 21332 18528
rect 21268 18468 21272 18524
rect 21272 18468 21328 18524
rect 21328 18468 21332 18524
rect 21268 18464 21332 18468
rect 27720 18524 27784 18528
rect 27720 18468 27724 18524
rect 27724 18468 27780 18524
rect 27780 18468 27784 18524
rect 27720 18464 27784 18468
rect 27800 18524 27864 18528
rect 27800 18468 27804 18524
rect 27804 18468 27860 18524
rect 27860 18468 27864 18524
rect 27800 18464 27864 18468
rect 27880 18524 27944 18528
rect 27880 18468 27884 18524
rect 27884 18468 27940 18524
rect 27940 18468 27944 18524
rect 27880 18464 27944 18468
rect 27960 18524 28024 18528
rect 27960 18468 27964 18524
rect 27964 18468 28020 18524
rect 28020 18468 28024 18524
rect 27960 18464 28024 18468
rect 4298 17980 4362 17984
rect 4298 17924 4302 17980
rect 4302 17924 4358 17980
rect 4358 17924 4362 17980
rect 4298 17920 4362 17924
rect 4378 17980 4442 17984
rect 4378 17924 4382 17980
rect 4382 17924 4438 17980
rect 4438 17924 4442 17980
rect 4378 17920 4442 17924
rect 4458 17980 4522 17984
rect 4458 17924 4462 17980
rect 4462 17924 4518 17980
rect 4518 17924 4522 17980
rect 4458 17920 4522 17924
rect 4538 17980 4602 17984
rect 4538 17924 4542 17980
rect 4542 17924 4598 17980
rect 4598 17924 4602 17980
rect 4538 17920 4602 17924
rect 10990 17980 11054 17984
rect 10990 17924 10994 17980
rect 10994 17924 11050 17980
rect 11050 17924 11054 17980
rect 10990 17920 11054 17924
rect 11070 17980 11134 17984
rect 11070 17924 11074 17980
rect 11074 17924 11130 17980
rect 11130 17924 11134 17980
rect 11070 17920 11134 17924
rect 11150 17980 11214 17984
rect 11150 17924 11154 17980
rect 11154 17924 11210 17980
rect 11210 17924 11214 17980
rect 11150 17920 11214 17924
rect 11230 17980 11294 17984
rect 11230 17924 11234 17980
rect 11234 17924 11290 17980
rect 11290 17924 11294 17980
rect 11230 17920 11294 17924
rect 17682 17980 17746 17984
rect 17682 17924 17686 17980
rect 17686 17924 17742 17980
rect 17742 17924 17746 17980
rect 17682 17920 17746 17924
rect 17762 17980 17826 17984
rect 17762 17924 17766 17980
rect 17766 17924 17822 17980
rect 17822 17924 17826 17980
rect 17762 17920 17826 17924
rect 17842 17980 17906 17984
rect 17842 17924 17846 17980
rect 17846 17924 17902 17980
rect 17902 17924 17906 17980
rect 17842 17920 17906 17924
rect 17922 17980 17986 17984
rect 17922 17924 17926 17980
rect 17926 17924 17982 17980
rect 17982 17924 17986 17980
rect 17922 17920 17986 17924
rect 24374 17980 24438 17984
rect 24374 17924 24378 17980
rect 24378 17924 24434 17980
rect 24434 17924 24438 17980
rect 24374 17920 24438 17924
rect 24454 17980 24518 17984
rect 24454 17924 24458 17980
rect 24458 17924 24514 17980
rect 24514 17924 24518 17980
rect 24454 17920 24518 17924
rect 24534 17980 24598 17984
rect 24534 17924 24538 17980
rect 24538 17924 24594 17980
rect 24594 17924 24598 17980
rect 24534 17920 24598 17924
rect 24614 17980 24678 17984
rect 24614 17924 24618 17980
rect 24618 17924 24674 17980
rect 24674 17924 24678 17980
rect 24614 17920 24678 17924
rect 7644 17436 7708 17440
rect 7644 17380 7648 17436
rect 7648 17380 7704 17436
rect 7704 17380 7708 17436
rect 7644 17376 7708 17380
rect 7724 17436 7788 17440
rect 7724 17380 7728 17436
rect 7728 17380 7784 17436
rect 7784 17380 7788 17436
rect 7724 17376 7788 17380
rect 7804 17436 7868 17440
rect 7804 17380 7808 17436
rect 7808 17380 7864 17436
rect 7864 17380 7868 17436
rect 7804 17376 7868 17380
rect 7884 17436 7948 17440
rect 7884 17380 7888 17436
rect 7888 17380 7944 17436
rect 7944 17380 7948 17436
rect 7884 17376 7948 17380
rect 14336 17436 14400 17440
rect 14336 17380 14340 17436
rect 14340 17380 14396 17436
rect 14396 17380 14400 17436
rect 14336 17376 14400 17380
rect 14416 17436 14480 17440
rect 14416 17380 14420 17436
rect 14420 17380 14476 17436
rect 14476 17380 14480 17436
rect 14416 17376 14480 17380
rect 14496 17436 14560 17440
rect 14496 17380 14500 17436
rect 14500 17380 14556 17436
rect 14556 17380 14560 17436
rect 14496 17376 14560 17380
rect 14576 17436 14640 17440
rect 14576 17380 14580 17436
rect 14580 17380 14636 17436
rect 14636 17380 14640 17436
rect 14576 17376 14640 17380
rect 21028 17436 21092 17440
rect 21028 17380 21032 17436
rect 21032 17380 21088 17436
rect 21088 17380 21092 17436
rect 21028 17376 21092 17380
rect 21108 17436 21172 17440
rect 21108 17380 21112 17436
rect 21112 17380 21168 17436
rect 21168 17380 21172 17436
rect 21108 17376 21172 17380
rect 21188 17436 21252 17440
rect 21188 17380 21192 17436
rect 21192 17380 21248 17436
rect 21248 17380 21252 17436
rect 21188 17376 21252 17380
rect 21268 17436 21332 17440
rect 21268 17380 21272 17436
rect 21272 17380 21328 17436
rect 21328 17380 21332 17436
rect 21268 17376 21332 17380
rect 27720 17436 27784 17440
rect 27720 17380 27724 17436
rect 27724 17380 27780 17436
rect 27780 17380 27784 17436
rect 27720 17376 27784 17380
rect 27800 17436 27864 17440
rect 27800 17380 27804 17436
rect 27804 17380 27860 17436
rect 27860 17380 27864 17436
rect 27800 17376 27864 17380
rect 27880 17436 27944 17440
rect 27880 17380 27884 17436
rect 27884 17380 27940 17436
rect 27940 17380 27944 17436
rect 27880 17376 27944 17380
rect 27960 17436 28024 17440
rect 27960 17380 27964 17436
rect 27964 17380 28020 17436
rect 28020 17380 28024 17436
rect 27960 17376 28024 17380
rect 4298 16892 4362 16896
rect 4298 16836 4302 16892
rect 4302 16836 4358 16892
rect 4358 16836 4362 16892
rect 4298 16832 4362 16836
rect 4378 16892 4442 16896
rect 4378 16836 4382 16892
rect 4382 16836 4438 16892
rect 4438 16836 4442 16892
rect 4378 16832 4442 16836
rect 4458 16892 4522 16896
rect 4458 16836 4462 16892
rect 4462 16836 4518 16892
rect 4518 16836 4522 16892
rect 4458 16832 4522 16836
rect 4538 16892 4602 16896
rect 4538 16836 4542 16892
rect 4542 16836 4598 16892
rect 4598 16836 4602 16892
rect 4538 16832 4602 16836
rect 10990 16892 11054 16896
rect 10990 16836 10994 16892
rect 10994 16836 11050 16892
rect 11050 16836 11054 16892
rect 10990 16832 11054 16836
rect 11070 16892 11134 16896
rect 11070 16836 11074 16892
rect 11074 16836 11130 16892
rect 11130 16836 11134 16892
rect 11070 16832 11134 16836
rect 11150 16892 11214 16896
rect 11150 16836 11154 16892
rect 11154 16836 11210 16892
rect 11210 16836 11214 16892
rect 11150 16832 11214 16836
rect 11230 16892 11294 16896
rect 11230 16836 11234 16892
rect 11234 16836 11290 16892
rect 11290 16836 11294 16892
rect 11230 16832 11294 16836
rect 17682 16892 17746 16896
rect 17682 16836 17686 16892
rect 17686 16836 17742 16892
rect 17742 16836 17746 16892
rect 17682 16832 17746 16836
rect 17762 16892 17826 16896
rect 17762 16836 17766 16892
rect 17766 16836 17822 16892
rect 17822 16836 17826 16892
rect 17762 16832 17826 16836
rect 17842 16892 17906 16896
rect 17842 16836 17846 16892
rect 17846 16836 17902 16892
rect 17902 16836 17906 16892
rect 17842 16832 17906 16836
rect 17922 16892 17986 16896
rect 17922 16836 17926 16892
rect 17926 16836 17982 16892
rect 17982 16836 17986 16892
rect 17922 16832 17986 16836
rect 24374 16892 24438 16896
rect 24374 16836 24378 16892
rect 24378 16836 24434 16892
rect 24434 16836 24438 16892
rect 24374 16832 24438 16836
rect 24454 16892 24518 16896
rect 24454 16836 24458 16892
rect 24458 16836 24514 16892
rect 24514 16836 24518 16892
rect 24454 16832 24518 16836
rect 24534 16892 24598 16896
rect 24534 16836 24538 16892
rect 24538 16836 24594 16892
rect 24594 16836 24598 16892
rect 24534 16832 24598 16836
rect 24614 16892 24678 16896
rect 24614 16836 24618 16892
rect 24618 16836 24674 16892
rect 24674 16836 24678 16892
rect 24614 16832 24678 16836
rect 7644 16348 7708 16352
rect 7644 16292 7648 16348
rect 7648 16292 7704 16348
rect 7704 16292 7708 16348
rect 7644 16288 7708 16292
rect 7724 16348 7788 16352
rect 7724 16292 7728 16348
rect 7728 16292 7784 16348
rect 7784 16292 7788 16348
rect 7724 16288 7788 16292
rect 7804 16348 7868 16352
rect 7804 16292 7808 16348
rect 7808 16292 7864 16348
rect 7864 16292 7868 16348
rect 7804 16288 7868 16292
rect 7884 16348 7948 16352
rect 7884 16292 7888 16348
rect 7888 16292 7944 16348
rect 7944 16292 7948 16348
rect 7884 16288 7948 16292
rect 14336 16348 14400 16352
rect 14336 16292 14340 16348
rect 14340 16292 14396 16348
rect 14396 16292 14400 16348
rect 14336 16288 14400 16292
rect 14416 16348 14480 16352
rect 14416 16292 14420 16348
rect 14420 16292 14476 16348
rect 14476 16292 14480 16348
rect 14416 16288 14480 16292
rect 14496 16348 14560 16352
rect 14496 16292 14500 16348
rect 14500 16292 14556 16348
rect 14556 16292 14560 16348
rect 14496 16288 14560 16292
rect 14576 16348 14640 16352
rect 14576 16292 14580 16348
rect 14580 16292 14636 16348
rect 14636 16292 14640 16348
rect 14576 16288 14640 16292
rect 21028 16348 21092 16352
rect 21028 16292 21032 16348
rect 21032 16292 21088 16348
rect 21088 16292 21092 16348
rect 21028 16288 21092 16292
rect 21108 16348 21172 16352
rect 21108 16292 21112 16348
rect 21112 16292 21168 16348
rect 21168 16292 21172 16348
rect 21108 16288 21172 16292
rect 21188 16348 21252 16352
rect 21188 16292 21192 16348
rect 21192 16292 21248 16348
rect 21248 16292 21252 16348
rect 21188 16288 21252 16292
rect 21268 16348 21332 16352
rect 21268 16292 21272 16348
rect 21272 16292 21328 16348
rect 21328 16292 21332 16348
rect 21268 16288 21332 16292
rect 27720 16348 27784 16352
rect 27720 16292 27724 16348
rect 27724 16292 27780 16348
rect 27780 16292 27784 16348
rect 27720 16288 27784 16292
rect 27800 16348 27864 16352
rect 27800 16292 27804 16348
rect 27804 16292 27860 16348
rect 27860 16292 27864 16348
rect 27800 16288 27864 16292
rect 27880 16348 27944 16352
rect 27880 16292 27884 16348
rect 27884 16292 27940 16348
rect 27940 16292 27944 16348
rect 27880 16288 27944 16292
rect 27960 16348 28024 16352
rect 27960 16292 27964 16348
rect 27964 16292 28020 16348
rect 28020 16292 28024 16348
rect 27960 16288 28024 16292
rect 4298 15804 4362 15808
rect 4298 15748 4302 15804
rect 4302 15748 4358 15804
rect 4358 15748 4362 15804
rect 4298 15744 4362 15748
rect 4378 15804 4442 15808
rect 4378 15748 4382 15804
rect 4382 15748 4438 15804
rect 4438 15748 4442 15804
rect 4378 15744 4442 15748
rect 4458 15804 4522 15808
rect 4458 15748 4462 15804
rect 4462 15748 4518 15804
rect 4518 15748 4522 15804
rect 4458 15744 4522 15748
rect 4538 15804 4602 15808
rect 4538 15748 4542 15804
rect 4542 15748 4598 15804
rect 4598 15748 4602 15804
rect 4538 15744 4602 15748
rect 10990 15804 11054 15808
rect 10990 15748 10994 15804
rect 10994 15748 11050 15804
rect 11050 15748 11054 15804
rect 10990 15744 11054 15748
rect 11070 15804 11134 15808
rect 11070 15748 11074 15804
rect 11074 15748 11130 15804
rect 11130 15748 11134 15804
rect 11070 15744 11134 15748
rect 11150 15804 11214 15808
rect 11150 15748 11154 15804
rect 11154 15748 11210 15804
rect 11210 15748 11214 15804
rect 11150 15744 11214 15748
rect 11230 15804 11294 15808
rect 11230 15748 11234 15804
rect 11234 15748 11290 15804
rect 11290 15748 11294 15804
rect 11230 15744 11294 15748
rect 17682 15804 17746 15808
rect 17682 15748 17686 15804
rect 17686 15748 17742 15804
rect 17742 15748 17746 15804
rect 17682 15744 17746 15748
rect 17762 15804 17826 15808
rect 17762 15748 17766 15804
rect 17766 15748 17822 15804
rect 17822 15748 17826 15804
rect 17762 15744 17826 15748
rect 17842 15804 17906 15808
rect 17842 15748 17846 15804
rect 17846 15748 17902 15804
rect 17902 15748 17906 15804
rect 17842 15744 17906 15748
rect 17922 15804 17986 15808
rect 17922 15748 17926 15804
rect 17926 15748 17982 15804
rect 17982 15748 17986 15804
rect 17922 15744 17986 15748
rect 24374 15804 24438 15808
rect 24374 15748 24378 15804
rect 24378 15748 24434 15804
rect 24434 15748 24438 15804
rect 24374 15744 24438 15748
rect 24454 15804 24518 15808
rect 24454 15748 24458 15804
rect 24458 15748 24514 15804
rect 24514 15748 24518 15804
rect 24454 15744 24518 15748
rect 24534 15804 24598 15808
rect 24534 15748 24538 15804
rect 24538 15748 24594 15804
rect 24594 15748 24598 15804
rect 24534 15744 24598 15748
rect 24614 15804 24678 15808
rect 24614 15748 24618 15804
rect 24618 15748 24674 15804
rect 24674 15748 24678 15804
rect 24614 15744 24678 15748
rect 7644 15260 7708 15264
rect 7644 15204 7648 15260
rect 7648 15204 7704 15260
rect 7704 15204 7708 15260
rect 7644 15200 7708 15204
rect 7724 15260 7788 15264
rect 7724 15204 7728 15260
rect 7728 15204 7784 15260
rect 7784 15204 7788 15260
rect 7724 15200 7788 15204
rect 7804 15260 7868 15264
rect 7804 15204 7808 15260
rect 7808 15204 7864 15260
rect 7864 15204 7868 15260
rect 7804 15200 7868 15204
rect 7884 15260 7948 15264
rect 7884 15204 7888 15260
rect 7888 15204 7944 15260
rect 7944 15204 7948 15260
rect 7884 15200 7948 15204
rect 14336 15260 14400 15264
rect 14336 15204 14340 15260
rect 14340 15204 14396 15260
rect 14396 15204 14400 15260
rect 14336 15200 14400 15204
rect 14416 15260 14480 15264
rect 14416 15204 14420 15260
rect 14420 15204 14476 15260
rect 14476 15204 14480 15260
rect 14416 15200 14480 15204
rect 14496 15260 14560 15264
rect 14496 15204 14500 15260
rect 14500 15204 14556 15260
rect 14556 15204 14560 15260
rect 14496 15200 14560 15204
rect 14576 15260 14640 15264
rect 14576 15204 14580 15260
rect 14580 15204 14636 15260
rect 14636 15204 14640 15260
rect 14576 15200 14640 15204
rect 21028 15260 21092 15264
rect 21028 15204 21032 15260
rect 21032 15204 21088 15260
rect 21088 15204 21092 15260
rect 21028 15200 21092 15204
rect 21108 15260 21172 15264
rect 21108 15204 21112 15260
rect 21112 15204 21168 15260
rect 21168 15204 21172 15260
rect 21108 15200 21172 15204
rect 21188 15260 21252 15264
rect 21188 15204 21192 15260
rect 21192 15204 21248 15260
rect 21248 15204 21252 15260
rect 21188 15200 21252 15204
rect 21268 15260 21332 15264
rect 21268 15204 21272 15260
rect 21272 15204 21328 15260
rect 21328 15204 21332 15260
rect 21268 15200 21332 15204
rect 27720 15260 27784 15264
rect 27720 15204 27724 15260
rect 27724 15204 27780 15260
rect 27780 15204 27784 15260
rect 27720 15200 27784 15204
rect 27800 15260 27864 15264
rect 27800 15204 27804 15260
rect 27804 15204 27860 15260
rect 27860 15204 27864 15260
rect 27800 15200 27864 15204
rect 27880 15260 27944 15264
rect 27880 15204 27884 15260
rect 27884 15204 27940 15260
rect 27940 15204 27944 15260
rect 27880 15200 27944 15204
rect 27960 15260 28024 15264
rect 27960 15204 27964 15260
rect 27964 15204 28020 15260
rect 28020 15204 28024 15260
rect 27960 15200 28024 15204
rect 4298 14716 4362 14720
rect 4298 14660 4302 14716
rect 4302 14660 4358 14716
rect 4358 14660 4362 14716
rect 4298 14656 4362 14660
rect 4378 14716 4442 14720
rect 4378 14660 4382 14716
rect 4382 14660 4438 14716
rect 4438 14660 4442 14716
rect 4378 14656 4442 14660
rect 4458 14716 4522 14720
rect 4458 14660 4462 14716
rect 4462 14660 4518 14716
rect 4518 14660 4522 14716
rect 4458 14656 4522 14660
rect 4538 14716 4602 14720
rect 4538 14660 4542 14716
rect 4542 14660 4598 14716
rect 4598 14660 4602 14716
rect 4538 14656 4602 14660
rect 10990 14716 11054 14720
rect 10990 14660 10994 14716
rect 10994 14660 11050 14716
rect 11050 14660 11054 14716
rect 10990 14656 11054 14660
rect 11070 14716 11134 14720
rect 11070 14660 11074 14716
rect 11074 14660 11130 14716
rect 11130 14660 11134 14716
rect 11070 14656 11134 14660
rect 11150 14716 11214 14720
rect 11150 14660 11154 14716
rect 11154 14660 11210 14716
rect 11210 14660 11214 14716
rect 11150 14656 11214 14660
rect 11230 14716 11294 14720
rect 11230 14660 11234 14716
rect 11234 14660 11290 14716
rect 11290 14660 11294 14716
rect 11230 14656 11294 14660
rect 17682 14716 17746 14720
rect 17682 14660 17686 14716
rect 17686 14660 17742 14716
rect 17742 14660 17746 14716
rect 17682 14656 17746 14660
rect 17762 14716 17826 14720
rect 17762 14660 17766 14716
rect 17766 14660 17822 14716
rect 17822 14660 17826 14716
rect 17762 14656 17826 14660
rect 17842 14716 17906 14720
rect 17842 14660 17846 14716
rect 17846 14660 17902 14716
rect 17902 14660 17906 14716
rect 17842 14656 17906 14660
rect 17922 14716 17986 14720
rect 17922 14660 17926 14716
rect 17926 14660 17982 14716
rect 17982 14660 17986 14716
rect 17922 14656 17986 14660
rect 24374 14716 24438 14720
rect 24374 14660 24378 14716
rect 24378 14660 24434 14716
rect 24434 14660 24438 14716
rect 24374 14656 24438 14660
rect 24454 14716 24518 14720
rect 24454 14660 24458 14716
rect 24458 14660 24514 14716
rect 24514 14660 24518 14716
rect 24454 14656 24518 14660
rect 24534 14716 24598 14720
rect 24534 14660 24538 14716
rect 24538 14660 24594 14716
rect 24594 14660 24598 14716
rect 24534 14656 24598 14660
rect 24614 14716 24678 14720
rect 24614 14660 24618 14716
rect 24618 14660 24674 14716
rect 24674 14660 24678 14716
rect 24614 14656 24678 14660
rect 7644 14172 7708 14176
rect 7644 14116 7648 14172
rect 7648 14116 7704 14172
rect 7704 14116 7708 14172
rect 7644 14112 7708 14116
rect 7724 14172 7788 14176
rect 7724 14116 7728 14172
rect 7728 14116 7784 14172
rect 7784 14116 7788 14172
rect 7724 14112 7788 14116
rect 7804 14172 7868 14176
rect 7804 14116 7808 14172
rect 7808 14116 7864 14172
rect 7864 14116 7868 14172
rect 7804 14112 7868 14116
rect 7884 14172 7948 14176
rect 7884 14116 7888 14172
rect 7888 14116 7944 14172
rect 7944 14116 7948 14172
rect 7884 14112 7948 14116
rect 14336 14172 14400 14176
rect 14336 14116 14340 14172
rect 14340 14116 14396 14172
rect 14396 14116 14400 14172
rect 14336 14112 14400 14116
rect 14416 14172 14480 14176
rect 14416 14116 14420 14172
rect 14420 14116 14476 14172
rect 14476 14116 14480 14172
rect 14416 14112 14480 14116
rect 14496 14172 14560 14176
rect 14496 14116 14500 14172
rect 14500 14116 14556 14172
rect 14556 14116 14560 14172
rect 14496 14112 14560 14116
rect 14576 14172 14640 14176
rect 14576 14116 14580 14172
rect 14580 14116 14636 14172
rect 14636 14116 14640 14172
rect 14576 14112 14640 14116
rect 21028 14172 21092 14176
rect 21028 14116 21032 14172
rect 21032 14116 21088 14172
rect 21088 14116 21092 14172
rect 21028 14112 21092 14116
rect 21108 14172 21172 14176
rect 21108 14116 21112 14172
rect 21112 14116 21168 14172
rect 21168 14116 21172 14172
rect 21108 14112 21172 14116
rect 21188 14172 21252 14176
rect 21188 14116 21192 14172
rect 21192 14116 21248 14172
rect 21248 14116 21252 14172
rect 21188 14112 21252 14116
rect 21268 14172 21332 14176
rect 21268 14116 21272 14172
rect 21272 14116 21328 14172
rect 21328 14116 21332 14172
rect 21268 14112 21332 14116
rect 27720 14172 27784 14176
rect 27720 14116 27724 14172
rect 27724 14116 27780 14172
rect 27780 14116 27784 14172
rect 27720 14112 27784 14116
rect 27800 14172 27864 14176
rect 27800 14116 27804 14172
rect 27804 14116 27860 14172
rect 27860 14116 27864 14172
rect 27800 14112 27864 14116
rect 27880 14172 27944 14176
rect 27880 14116 27884 14172
rect 27884 14116 27940 14172
rect 27940 14116 27944 14172
rect 27880 14112 27944 14116
rect 27960 14172 28024 14176
rect 27960 14116 27964 14172
rect 27964 14116 28020 14172
rect 28020 14116 28024 14172
rect 27960 14112 28024 14116
rect 4298 13628 4362 13632
rect 4298 13572 4302 13628
rect 4302 13572 4358 13628
rect 4358 13572 4362 13628
rect 4298 13568 4362 13572
rect 4378 13628 4442 13632
rect 4378 13572 4382 13628
rect 4382 13572 4438 13628
rect 4438 13572 4442 13628
rect 4378 13568 4442 13572
rect 4458 13628 4522 13632
rect 4458 13572 4462 13628
rect 4462 13572 4518 13628
rect 4518 13572 4522 13628
rect 4458 13568 4522 13572
rect 4538 13628 4602 13632
rect 4538 13572 4542 13628
rect 4542 13572 4598 13628
rect 4598 13572 4602 13628
rect 4538 13568 4602 13572
rect 10990 13628 11054 13632
rect 10990 13572 10994 13628
rect 10994 13572 11050 13628
rect 11050 13572 11054 13628
rect 10990 13568 11054 13572
rect 11070 13628 11134 13632
rect 11070 13572 11074 13628
rect 11074 13572 11130 13628
rect 11130 13572 11134 13628
rect 11070 13568 11134 13572
rect 11150 13628 11214 13632
rect 11150 13572 11154 13628
rect 11154 13572 11210 13628
rect 11210 13572 11214 13628
rect 11150 13568 11214 13572
rect 11230 13628 11294 13632
rect 11230 13572 11234 13628
rect 11234 13572 11290 13628
rect 11290 13572 11294 13628
rect 11230 13568 11294 13572
rect 17682 13628 17746 13632
rect 17682 13572 17686 13628
rect 17686 13572 17742 13628
rect 17742 13572 17746 13628
rect 17682 13568 17746 13572
rect 17762 13628 17826 13632
rect 17762 13572 17766 13628
rect 17766 13572 17822 13628
rect 17822 13572 17826 13628
rect 17762 13568 17826 13572
rect 17842 13628 17906 13632
rect 17842 13572 17846 13628
rect 17846 13572 17902 13628
rect 17902 13572 17906 13628
rect 17842 13568 17906 13572
rect 17922 13628 17986 13632
rect 17922 13572 17926 13628
rect 17926 13572 17982 13628
rect 17982 13572 17986 13628
rect 17922 13568 17986 13572
rect 24374 13628 24438 13632
rect 24374 13572 24378 13628
rect 24378 13572 24434 13628
rect 24434 13572 24438 13628
rect 24374 13568 24438 13572
rect 24454 13628 24518 13632
rect 24454 13572 24458 13628
rect 24458 13572 24514 13628
rect 24514 13572 24518 13628
rect 24454 13568 24518 13572
rect 24534 13628 24598 13632
rect 24534 13572 24538 13628
rect 24538 13572 24594 13628
rect 24594 13572 24598 13628
rect 24534 13568 24598 13572
rect 24614 13628 24678 13632
rect 24614 13572 24618 13628
rect 24618 13572 24674 13628
rect 24674 13572 24678 13628
rect 24614 13568 24678 13572
rect 7644 13084 7708 13088
rect 7644 13028 7648 13084
rect 7648 13028 7704 13084
rect 7704 13028 7708 13084
rect 7644 13024 7708 13028
rect 7724 13084 7788 13088
rect 7724 13028 7728 13084
rect 7728 13028 7784 13084
rect 7784 13028 7788 13084
rect 7724 13024 7788 13028
rect 7804 13084 7868 13088
rect 7804 13028 7808 13084
rect 7808 13028 7864 13084
rect 7864 13028 7868 13084
rect 7804 13024 7868 13028
rect 7884 13084 7948 13088
rect 7884 13028 7888 13084
rect 7888 13028 7944 13084
rect 7944 13028 7948 13084
rect 7884 13024 7948 13028
rect 14336 13084 14400 13088
rect 14336 13028 14340 13084
rect 14340 13028 14396 13084
rect 14396 13028 14400 13084
rect 14336 13024 14400 13028
rect 14416 13084 14480 13088
rect 14416 13028 14420 13084
rect 14420 13028 14476 13084
rect 14476 13028 14480 13084
rect 14416 13024 14480 13028
rect 14496 13084 14560 13088
rect 14496 13028 14500 13084
rect 14500 13028 14556 13084
rect 14556 13028 14560 13084
rect 14496 13024 14560 13028
rect 14576 13084 14640 13088
rect 14576 13028 14580 13084
rect 14580 13028 14636 13084
rect 14636 13028 14640 13084
rect 14576 13024 14640 13028
rect 21028 13084 21092 13088
rect 21028 13028 21032 13084
rect 21032 13028 21088 13084
rect 21088 13028 21092 13084
rect 21028 13024 21092 13028
rect 21108 13084 21172 13088
rect 21108 13028 21112 13084
rect 21112 13028 21168 13084
rect 21168 13028 21172 13084
rect 21108 13024 21172 13028
rect 21188 13084 21252 13088
rect 21188 13028 21192 13084
rect 21192 13028 21248 13084
rect 21248 13028 21252 13084
rect 21188 13024 21252 13028
rect 21268 13084 21332 13088
rect 21268 13028 21272 13084
rect 21272 13028 21328 13084
rect 21328 13028 21332 13084
rect 21268 13024 21332 13028
rect 27720 13084 27784 13088
rect 27720 13028 27724 13084
rect 27724 13028 27780 13084
rect 27780 13028 27784 13084
rect 27720 13024 27784 13028
rect 27800 13084 27864 13088
rect 27800 13028 27804 13084
rect 27804 13028 27860 13084
rect 27860 13028 27864 13084
rect 27800 13024 27864 13028
rect 27880 13084 27944 13088
rect 27880 13028 27884 13084
rect 27884 13028 27940 13084
rect 27940 13028 27944 13084
rect 27880 13024 27944 13028
rect 27960 13084 28024 13088
rect 27960 13028 27964 13084
rect 27964 13028 28020 13084
rect 28020 13028 28024 13084
rect 27960 13024 28024 13028
rect 4298 12540 4362 12544
rect 4298 12484 4302 12540
rect 4302 12484 4358 12540
rect 4358 12484 4362 12540
rect 4298 12480 4362 12484
rect 4378 12540 4442 12544
rect 4378 12484 4382 12540
rect 4382 12484 4438 12540
rect 4438 12484 4442 12540
rect 4378 12480 4442 12484
rect 4458 12540 4522 12544
rect 4458 12484 4462 12540
rect 4462 12484 4518 12540
rect 4518 12484 4522 12540
rect 4458 12480 4522 12484
rect 4538 12540 4602 12544
rect 4538 12484 4542 12540
rect 4542 12484 4598 12540
rect 4598 12484 4602 12540
rect 4538 12480 4602 12484
rect 10990 12540 11054 12544
rect 10990 12484 10994 12540
rect 10994 12484 11050 12540
rect 11050 12484 11054 12540
rect 10990 12480 11054 12484
rect 11070 12540 11134 12544
rect 11070 12484 11074 12540
rect 11074 12484 11130 12540
rect 11130 12484 11134 12540
rect 11070 12480 11134 12484
rect 11150 12540 11214 12544
rect 11150 12484 11154 12540
rect 11154 12484 11210 12540
rect 11210 12484 11214 12540
rect 11150 12480 11214 12484
rect 11230 12540 11294 12544
rect 11230 12484 11234 12540
rect 11234 12484 11290 12540
rect 11290 12484 11294 12540
rect 11230 12480 11294 12484
rect 17682 12540 17746 12544
rect 17682 12484 17686 12540
rect 17686 12484 17742 12540
rect 17742 12484 17746 12540
rect 17682 12480 17746 12484
rect 17762 12540 17826 12544
rect 17762 12484 17766 12540
rect 17766 12484 17822 12540
rect 17822 12484 17826 12540
rect 17762 12480 17826 12484
rect 17842 12540 17906 12544
rect 17842 12484 17846 12540
rect 17846 12484 17902 12540
rect 17902 12484 17906 12540
rect 17842 12480 17906 12484
rect 17922 12540 17986 12544
rect 17922 12484 17926 12540
rect 17926 12484 17982 12540
rect 17982 12484 17986 12540
rect 17922 12480 17986 12484
rect 24374 12540 24438 12544
rect 24374 12484 24378 12540
rect 24378 12484 24434 12540
rect 24434 12484 24438 12540
rect 24374 12480 24438 12484
rect 24454 12540 24518 12544
rect 24454 12484 24458 12540
rect 24458 12484 24514 12540
rect 24514 12484 24518 12540
rect 24454 12480 24518 12484
rect 24534 12540 24598 12544
rect 24534 12484 24538 12540
rect 24538 12484 24594 12540
rect 24594 12484 24598 12540
rect 24534 12480 24598 12484
rect 24614 12540 24678 12544
rect 24614 12484 24618 12540
rect 24618 12484 24674 12540
rect 24674 12484 24678 12540
rect 24614 12480 24678 12484
rect 7644 11996 7708 12000
rect 7644 11940 7648 11996
rect 7648 11940 7704 11996
rect 7704 11940 7708 11996
rect 7644 11936 7708 11940
rect 7724 11996 7788 12000
rect 7724 11940 7728 11996
rect 7728 11940 7784 11996
rect 7784 11940 7788 11996
rect 7724 11936 7788 11940
rect 7804 11996 7868 12000
rect 7804 11940 7808 11996
rect 7808 11940 7864 11996
rect 7864 11940 7868 11996
rect 7804 11936 7868 11940
rect 7884 11996 7948 12000
rect 7884 11940 7888 11996
rect 7888 11940 7944 11996
rect 7944 11940 7948 11996
rect 7884 11936 7948 11940
rect 14336 11996 14400 12000
rect 14336 11940 14340 11996
rect 14340 11940 14396 11996
rect 14396 11940 14400 11996
rect 14336 11936 14400 11940
rect 14416 11996 14480 12000
rect 14416 11940 14420 11996
rect 14420 11940 14476 11996
rect 14476 11940 14480 11996
rect 14416 11936 14480 11940
rect 14496 11996 14560 12000
rect 14496 11940 14500 11996
rect 14500 11940 14556 11996
rect 14556 11940 14560 11996
rect 14496 11936 14560 11940
rect 14576 11996 14640 12000
rect 14576 11940 14580 11996
rect 14580 11940 14636 11996
rect 14636 11940 14640 11996
rect 14576 11936 14640 11940
rect 21028 11996 21092 12000
rect 21028 11940 21032 11996
rect 21032 11940 21088 11996
rect 21088 11940 21092 11996
rect 21028 11936 21092 11940
rect 21108 11996 21172 12000
rect 21108 11940 21112 11996
rect 21112 11940 21168 11996
rect 21168 11940 21172 11996
rect 21108 11936 21172 11940
rect 21188 11996 21252 12000
rect 21188 11940 21192 11996
rect 21192 11940 21248 11996
rect 21248 11940 21252 11996
rect 21188 11936 21252 11940
rect 21268 11996 21332 12000
rect 21268 11940 21272 11996
rect 21272 11940 21328 11996
rect 21328 11940 21332 11996
rect 21268 11936 21332 11940
rect 27720 11996 27784 12000
rect 27720 11940 27724 11996
rect 27724 11940 27780 11996
rect 27780 11940 27784 11996
rect 27720 11936 27784 11940
rect 27800 11996 27864 12000
rect 27800 11940 27804 11996
rect 27804 11940 27860 11996
rect 27860 11940 27864 11996
rect 27800 11936 27864 11940
rect 27880 11996 27944 12000
rect 27880 11940 27884 11996
rect 27884 11940 27940 11996
rect 27940 11940 27944 11996
rect 27880 11936 27944 11940
rect 27960 11996 28024 12000
rect 27960 11940 27964 11996
rect 27964 11940 28020 11996
rect 28020 11940 28024 11996
rect 27960 11936 28024 11940
rect 4298 11452 4362 11456
rect 4298 11396 4302 11452
rect 4302 11396 4358 11452
rect 4358 11396 4362 11452
rect 4298 11392 4362 11396
rect 4378 11452 4442 11456
rect 4378 11396 4382 11452
rect 4382 11396 4438 11452
rect 4438 11396 4442 11452
rect 4378 11392 4442 11396
rect 4458 11452 4522 11456
rect 4458 11396 4462 11452
rect 4462 11396 4518 11452
rect 4518 11396 4522 11452
rect 4458 11392 4522 11396
rect 4538 11452 4602 11456
rect 4538 11396 4542 11452
rect 4542 11396 4598 11452
rect 4598 11396 4602 11452
rect 4538 11392 4602 11396
rect 10990 11452 11054 11456
rect 10990 11396 10994 11452
rect 10994 11396 11050 11452
rect 11050 11396 11054 11452
rect 10990 11392 11054 11396
rect 11070 11452 11134 11456
rect 11070 11396 11074 11452
rect 11074 11396 11130 11452
rect 11130 11396 11134 11452
rect 11070 11392 11134 11396
rect 11150 11452 11214 11456
rect 11150 11396 11154 11452
rect 11154 11396 11210 11452
rect 11210 11396 11214 11452
rect 11150 11392 11214 11396
rect 11230 11452 11294 11456
rect 11230 11396 11234 11452
rect 11234 11396 11290 11452
rect 11290 11396 11294 11452
rect 11230 11392 11294 11396
rect 17682 11452 17746 11456
rect 17682 11396 17686 11452
rect 17686 11396 17742 11452
rect 17742 11396 17746 11452
rect 17682 11392 17746 11396
rect 17762 11452 17826 11456
rect 17762 11396 17766 11452
rect 17766 11396 17822 11452
rect 17822 11396 17826 11452
rect 17762 11392 17826 11396
rect 17842 11452 17906 11456
rect 17842 11396 17846 11452
rect 17846 11396 17902 11452
rect 17902 11396 17906 11452
rect 17842 11392 17906 11396
rect 17922 11452 17986 11456
rect 17922 11396 17926 11452
rect 17926 11396 17982 11452
rect 17982 11396 17986 11452
rect 17922 11392 17986 11396
rect 24374 11452 24438 11456
rect 24374 11396 24378 11452
rect 24378 11396 24434 11452
rect 24434 11396 24438 11452
rect 24374 11392 24438 11396
rect 24454 11452 24518 11456
rect 24454 11396 24458 11452
rect 24458 11396 24514 11452
rect 24514 11396 24518 11452
rect 24454 11392 24518 11396
rect 24534 11452 24598 11456
rect 24534 11396 24538 11452
rect 24538 11396 24594 11452
rect 24594 11396 24598 11452
rect 24534 11392 24598 11396
rect 24614 11452 24678 11456
rect 24614 11396 24618 11452
rect 24618 11396 24674 11452
rect 24674 11396 24678 11452
rect 24614 11392 24678 11396
rect 7644 10908 7708 10912
rect 7644 10852 7648 10908
rect 7648 10852 7704 10908
rect 7704 10852 7708 10908
rect 7644 10848 7708 10852
rect 7724 10908 7788 10912
rect 7724 10852 7728 10908
rect 7728 10852 7784 10908
rect 7784 10852 7788 10908
rect 7724 10848 7788 10852
rect 7804 10908 7868 10912
rect 7804 10852 7808 10908
rect 7808 10852 7864 10908
rect 7864 10852 7868 10908
rect 7804 10848 7868 10852
rect 7884 10908 7948 10912
rect 7884 10852 7888 10908
rect 7888 10852 7944 10908
rect 7944 10852 7948 10908
rect 7884 10848 7948 10852
rect 14336 10908 14400 10912
rect 14336 10852 14340 10908
rect 14340 10852 14396 10908
rect 14396 10852 14400 10908
rect 14336 10848 14400 10852
rect 14416 10908 14480 10912
rect 14416 10852 14420 10908
rect 14420 10852 14476 10908
rect 14476 10852 14480 10908
rect 14416 10848 14480 10852
rect 14496 10908 14560 10912
rect 14496 10852 14500 10908
rect 14500 10852 14556 10908
rect 14556 10852 14560 10908
rect 14496 10848 14560 10852
rect 14576 10908 14640 10912
rect 14576 10852 14580 10908
rect 14580 10852 14636 10908
rect 14636 10852 14640 10908
rect 14576 10848 14640 10852
rect 21028 10908 21092 10912
rect 21028 10852 21032 10908
rect 21032 10852 21088 10908
rect 21088 10852 21092 10908
rect 21028 10848 21092 10852
rect 21108 10908 21172 10912
rect 21108 10852 21112 10908
rect 21112 10852 21168 10908
rect 21168 10852 21172 10908
rect 21108 10848 21172 10852
rect 21188 10908 21252 10912
rect 21188 10852 21192 10908
rect 21192 10852 21248 10908
rect 21248 10852 21252 10908
rect 21188 10848 21252 10852
rect 21268 10908 21332 10912
rect 21268 10852 21272 10908
rect 21272 10852 21328 10908
rect 21328 10852 21332 10908
rect 21268 10848 21332 10852
rect 27720 10908 27784 10912
rect 27720 10852 27724 10908
rect 27724 10852 27780 10908
rect 27780 10852 27784 10908
rect 27720 10848 27784 10852
rect 27800 10908 27864 10912
rect 27800 10852 27804 10908
rect 27804 10852 27860 10908
rect 27860 10852 27864 10908
rect 27800 10848 27864 10852
rect 27880 10908 27944 10912
rect 27880 10852 27884 10908
rect 27884 10852 27940 10908
rect 27940 10852 27944 10908
rect 27880 10848 27944 10852
rect 27960 10908 28024 10912
rect 27960 10852 27964 10908
rect 27964 10852 28020 10908
rect 28020 10852 28024 10908
rect 27960 10848 28024 10852
rect 4298 10364 4362 10368
rect 4298 10308 4302 10364
rect 4302 10308 4358 10364
rect 4358 10308 4362 10364
rect 4298 10304 4362 10308
rect 4378 10364 4442 10368
rect 4378 10308 4382 10364
rect 4382 10308 4438 10364
rect 4438 10308 4442 10364
rect 4378 10304 4442 10308
rect 4458 10364 4522 10368
rect 4458 10308 4462 10364
rect 4462 10308 4518 10364
rect 4518 10308 4522 10364
rect 4458 10304 4522 10308
rect 4538 10364 4602 10368
rect 4538 10308 4542 10364
rect 4542 10308 4598 10364
rect 4598 10308 4602 10364
rect 4538 10304 4602 10308
rect 10990 10364 11054 10368
rect 10990 10308 10994 10364
rect 10994 10308 11050 10364
rect 11050 10308 11054 10364
rect 10990 10304 11054 10308
rect 11070 10364 11134 10368
rect 11070 10308 11074 10364
rect 11074 10308 11130 10364
rect 11130 10308 11134 10364
rect 11070 10304 11134 10308
rect 11150 10364 11214 10368
rect 11150 10308 11154 10364
rect 11154 10308 11210 10364
rect 11210 10308 11214 10364
rect 11150 10304 11214 10308
rect 11230 10364 11294 10368
rect 11230 10308 11234 10364
rect 11234 10308 11290 10364
rect 11290 10308 11294 10364
rect 11230 10304 11294 10308
rect 17682 10364 17746 10368
rect 17682 10308 17686 10364
rect 17686 10308 17742 10364
rect 17742 10308 17746 10364
rect 17682 10304 17746 10308
rect 17762 10364 17826 10368
rect 17762 10308 17766 10364
rect 17766 10308 17822 10364
rect 17822 10308 17826 10364
rect 17762 10304 17826 10308
rect 17842 10364 17906 10368
rect 17842 10308 17846 10364
rect 17846 10308 17902 10364
rect 17902 10308 17906 10364
rect 17842 10304 17906 10308
rect 17922 10364 17986 10368
rect 17922 10308 17926 10364
rect 17926 10308 17982 10364
rect 17982 10308 17986 10364
rect 17922 10304 17986 10308
rect 24374 10364 24438 10368
rect 24374 10308 24378 10364
rect 24378 10308 24434 10364
rect 24434 10308 24438 10364
rect 24374 10304 24438 10308
rect 24454 10364 24518 10368
rect 24454 10308 24458 10364
rect 24458 10308 24514 10364
rect 24514 10308 24518 10364
rect 24454 10304 24518 10308
rect 24534 10364 24598 10368
rect 24534 10308 24538 10364
rect 24538 10308 24594 10364
rect 24594 10308 24598 10364
rect 24534 10304 24598 10308
rect 24614 10364 24678 10368
rect 24614 10308 24618 10364
rect 24618 10308 24674 10364
rect 24674 10308 24678 10364
rect 24614 10304 24678 10308
rect 7644 9820 7708 9824
rect 7644 9764 7648 9820
rect 7648 9764 7704 9820
rect 7704 9764 7708 9820
rect 7644 9760 7708 9764
rect 7724 9820 7788 9824
rect 7724 9764 7728 9820
rect 7728 9764 7784 9820
rect 7784 9764 7788 9820
rect 7724 9760 7788 9764
rect 7804 9820 7868 9824
rect 7804 9764 7808 9820
rect 7808 9764 7864 9820
rect 7864 9764 7868 9820
rect 7804 9760 7868 9764
rect 7884 9820 7948 9824
rect 7884 9764 7888 9820
rect 7888 9764 7944 9820
rect 7944 9764 7948 9820
rect 7884 9760 7948 9764
rect 14336 9820 14400 9824
rect 14336 9764 14340 9820
rect 14340 9764 14396 9820
rect 14396 9764 14400 9820
rect 14336 9760 14400 9764
rect 14416 9820 14480 9824
rect 14416 9764 14420 9820
rect 14420 9764 14476 9820
rect 14476 9764 14480 9820
rect 14416 9760 14480 9764
rect 14496 9820 14560 9824
rect 14496 9764 14500 9820
rect 14500 9764 14556 9820
rect 14556 9764 14560 9820
rect 14496 9760 14560 9764
rect 14576 9820 14640 9824
rect 14576 9764 14580 9820
rect 14580 9764 14636 9820
rect 14636 9764 14640 9820
rect 14576 9760 14640 9764
rect 21028 9820 21092 9824
rect 21028 9764 21032 9820
rect 21032 9764 21088 9820
rect 21088 9764 21092 9820
rect 21028 9760 21092 9764
rect 21108 9820 21172 9824
rect 21108 9764 21112 9820
rect 21112 9764 21168 9820
rect 21168 9764 21172 9820
rect 21108 9760 21172 9764
rect 21188 9820 21252 9824
rect 21188 9764 21192 9820
rect 21192 9764 21248 9820
rect 21248 9764 21252 9820
rect 21188 9760 21252 9764
rect 21268 9820 21332 9824
rect 21268 9764 21272 9820
rect 21272 9764 21328 9820
rect 21328 9764 21332 9820
rect 21268 9760 21332 9764
rect 27720 9820 27784 9824
rect 27720 9764 27724 9820
rect 27724 9764 27780 9820
rect 27780 9764 27784 9820
rect 27720 9760 27784 9764
rect 27800 9820 27864 9824
rect 27800 9764 27804 9820
rect 27804 9764 27860 9820
rect 27860 9764 27864 9820
rect 27800 9760 27864 9764
rect 27880 9820 27944 9824
rect 27880 9764 27884 9820
rect 27884 9764 27940 9820
rect 27940 9764 27944 9820
rect 27880 9760 27944 9764
rect 27960 9820 28024 9824
rect 27960 9764 27964 9820
rect 27964 9764 28020 9820
rect 28020 9764 28024 9820
rect 27960 9760 28024 9764
rect 4298 9276 4362 9280
rect 4298 9220 4302 9276
rect 4302 9220 4358 9276
rect 4358 9220 4362 9276
rect 4298 9216 4362 9220
rect 4378 9276 4442 9280
rect 4378 9220 4382 9276
rect 4382 9220 4438 9276
rect 4438 9220 4442 9276
rect 4378 9216 4442 9220
rect 4458 9276 4522 9280
rect 4458 9220 4462 9276
rect 4462 9220 4518 9276
rect 4518 9220 4522 9276
rect 4458 9216 4522 9220
rect 4538 9276 4602 9280
rect 4538 9220 4542 9276
rect 4542 9220 4598 9276
rect 4598 9220 4602 9276
rect 4538 9216 4602 9220
rect 10990 9276 11054 9280
rect 10990 9220 10994 9276
rect 10994 9220 11050 9276
rect 11050 9220 11054 9276
rect 10990 9216 11054 9220
rect 11070 9276 11134 9280
rect 11070 9220 11074 9276
rect 11074 9220 11130 9276
rect 11130 9220 11134 9276
rect 11070 9216 11134 9220
rect 11150 9276 11214 9280
rect 11150 9220 11154 9276
rect 11154 9220 11210 9276
rect 11210 9220 11214 9276
rect 11150 9216 11214 9220
rect 11230 9276 11294 9280
rect 11230 9220 11234 9276
rect 11234 9220 11290 9276
rect 11290 9220 11294 9276
rect 11230 9216 11294 9220
rect 17682 9276 17746 9280
rect 17682 9220 17686 9276
rect 17686 9220 17742 9276
rect 17742 9220 17746 9276
rect 17682 9216 17746 9220
rect 17762 9276 17826 9280
rect 17762 9220 17766 9276
rect 17766 9220 17822 9276
rect 17822 9220 17826 9276
rect 17762 9216 17826 9220
rect 17842 9276 17906 9280
rect 17842 9220 17846 9276
rect 17846 9220 17902 9276
rect 17902 9220 17906 9276
rect 17842 9216 17906 9220
rect 17922 9276 17986 9280
rect 17922 9220 17926 9276
rect 17926 9220 17982 9276
rect 17982 9220 17986 9276
rect 17922 9216 17986 9220
rect 24374 9276 24438 9280
rect 24374 9220 24378 9276
rect 24378 9220 24434 9276
rect 24434 9220 24438 9276
rect 24374 9216 24438 9220
rect 24454 9276 24518 9280
rect 24454 9220 24458 9276
rect 24458 9220 24514 9276
rect 24514 9220 24518 9276
rect 24454 9216 24518 9220
rect 24534 9276 24598 9280
rect 24534 9220 24538 9276
rect 24538 9220 24594 9276
rect 24594 9220 24598 9276
rect 24534 9216 24598 9220
rect 24614 9276 24678 9280
rect 24614 9220 24618 9276
rect 24618 9220 24674 9276
rect 24674 9220 24678 9276
rect 24614 9216 24678 9220
rect 7644 8732 7708 8736
rect 7644 8676 7648 8732
rect 7648 8676 7704 8732
rect 7704 8676 7708 8732
rect 7644 8672 7708 8676
rect 7724 8732 7788 8736
rect 7724 8676 7728 8732
rect 7728 8676 7784 8732
rect 7784 8676 7788 8732
rect 7724 8672 7788 8676
rect 7804 8732 7868 8736
rect 7804 8676 7808 8732
rect 7808 8676 7864 8732
rect 7864 8676 7868 8732
rect 7804 8672 7868 8676
rect 7884 8732 7948 8736
rect 7884 8676 7888 8732
rect 7888 8676 7944 8732
rect 7944 8676 7948 8732
rect 7884 8672 7948 8676
rect 14336 8732 14400 8736
rect 14336 8676 14340 8732
rect 14340 8676 14396 8732
rect 14396 8676 14400 8732
rect 14336 8672 14400 8676
rect 14416 8732 14480 8736
rect 14416 8676 14420 8732
rect 14420 8676 14476 8732
rect 14476 8676 14480 8732
rect 14416 8672 14480 8676
rect 14496 8732 14560 8736
rect 14496 8676 14500 8732
rect 14500 8676 14556 8732
rect 14556 8676 14560 8732
rect 14496 8672 14560 8676
rect 14576 8732 14640 8736
rect 14576 8676 14580 8732
rect 14580 8676 14636 8732
rect 14636 8676 14640 8732
rect 14576 8672 14640 8676
rect 21028 8732 21092 8736
rect 21028 8676 21032 8732
rect 21032 8676 21088 8732
rect 21088 8676 21092 8732
rect 21028 8672 21092 8676
rect 21108 8732 21172 8736
rect 21108 8676 21112 8732
rect 21112 8676 21168 8732
rect 21168 8676 21172 8732
rect 21108 8672 21172 8676
rect 21188 8732 21252 8736
rect 21188 8676 21192 8732
rect 21192 8676 21248 8732
rect 21248 8676 21252 8732
rect 21188 8672 21252 8676
rect 21268 8732 21332 8736
rect 21268 8676 21272 8732
rect 21272 8676 21328 8732
rect 21328 8676 21332 8732
rect 21268 8672 21332 8676
rect 27720 8732 27784 8736
rect 27720 8676 27724 8732
rect 27724 8676 27780 8732
rect 27780 8676 27784 8732
rect 27720 8672 27784 8676
rect 27800 8732 27864 8736
rect 27800 8676 27804 8732
rect 27804 8676 27860 8732
rect 27860 8676 27864 8732
rect 27800 8672 27864 8676
rect 27880 8732 27944 8736
rect 27880 8676 27884 8732
rect 27884 8676 27940 8732
rect 27940 8676 27944 8732
rect 27880 8672 27944 8676
rect 27960 8732 28024 8736
rect 27960 8676 27964 8732
rect 27964 8676 28020 8732
rect 28020 8676 28024 8732
rect 27960 8672 28024 8676
rect 4298 8188 4362 8192
rect 4298 8132 4302 8188
rect 4302 8132 4358 8188
rect 4358 8132 4362 8188
rect 4298 8128 4362 8132
rect 4378 8188 4442 8192
rect 4378 8132 4382 8188
rect 4382 8132 4438 8188
rect 4438 8132 4442 8188
rect 4378 8128 4442 8132
rect 4458 8188 4522 8192
rect 4458 8132 4462 8188
rect 4462 8132 4518 8188
rect 4518 8132 4522 8188
rect 4458 8128 4522 8132
rect 4538 8188 4602 8192
rect 4538 8132 4542 8188
rect 4542 8132 4598 8188
rect 4598 8132 4602 8188
rect 4538 8128 4602 8132
rect 10990 8188 11054 8192
rect 10990 8132 10994 8188
rect 10994 8132 11050 8188
rect 11050 8132 11054 8188
rect 10990 8128 11054 8132
rect 11070 8188 11134 8192
rect 11070 8132 11074 8188
rect 11074 8132 11130 8188
rect 11130 8132 11134 8188
rect 11070 8128 11134 8132
rect 11150 8188 11214 8192
rect 11150 8132 11154 8188
rect 11154 8132 11210 8188
rect 11210 8132 11214 8188
rect 11150 8128 11214 8132
rect 11230 8188 11294 8192
rect 11230 8132 11234 8188
rect 11234 8132 11290 8188
rect 11290 8132 11294 8188
rect 11230 8128 11294 8132
rect 17682 8188 17746 8192
rect 17682 8132 17686 8188
rect 17686 8132 17742 8188
rect 17742 8132 17746 8188
rect 17682 8128 17746 8132
rect 17762 8188 17826 8192
rect 17762 8132 17766 8188
rect 17766 8132 17822 8188
rect 17822 8132 17826 8188
rect 17762 8128 17826 8132
rect 17842 8188 17906 8192
rect 17842 8132 17846 8188
rect 17846 8132 17902 8188
rect 17902 8132 17906 8188
rect 17842 8128 17906 8132
rect 17922 8188 17986 8192
rect 17922 8132 17926 8188
rect 17926 8132 17982 8188
rect 17982 8132 17986 8188
rect 17922 8128 17986 8132
rect 24374 8188 24438 8192
rect 24374 8132 24378 8188
rect 24378 8132 24434 8188
rect 24434 8132 24438 8188
rect 24374 8128 24438 8132
rect 24454 8188 24518 8192
rect 24454 8132 24458 8188
rect 24458 8132 24514 8188
rect 24514 8132 24518 8188
rect 24454 8128 24518 8132
rect 24534 8188 24598 8192
rect 24534 8132 24538 8188
rect 24538 8132 24594 8188
rect 24594 8132 24598 8188
rect 24534 8128 24598 8132
rect 24614 8188 24678 8192
rect 24614 8132 24618 8188
rect 24618 8132 24674 8188
rect 24674 8132 24678 8188
rect 24614 8128 24678 8132
rect 7644 7644 7708 7648
rect 7644 7588 7648 7644
rect 7648 7588 7704 7644
rect 7704 7588 7708 7644
rect 7644 7584 7708 7588
rect 7724 7644 7788 7648
rect 7724 7588 7728 7644
rect 7728 7588 7784 7644
rect 7784 7588 7788 7644
rect 7724 7584 7788 7588
rect 7804 7644 7868 7648
rect 7804 7588 7808 7644
rect 7808 7588 7864 7644
rect 7864 7588 7868 7644
rect 7804 7584 7868 7588
rect 7884 7644 7948 7648
rect 7884 7588 7888 7644
rect 7888 7588 7944 7644
rect 7944 7588 7948 7644
rect 7884 7584 7948 7588
rect 14336 7644 14400 7648
rect 14336 7588 14340 7644
rect 14340 7588 14396 7644
rect 14396 7588 14400 7644
rect 14336 7584 14400 7588
rect 14416 7644 14480 7648
rect 14416 7588 14420 7644
rect 14420 7588 14476 7644
rect 14476 7588 14480 7644
rect 14416 7584 14480 7588
rect 14496 7644 14560 7648
rect 14496 7588 14500 7644
rect 14500 7588 14556 7644
rect 14556 7588 14560 7644
rect 14496 7584 14560 7588
rect 14576 7644 14640 7648
rect 14576 7588 14580 7644
rect 14580 7588 14636 7644
rect 14636 7588 14640 7644
rect 14576 7584 14640 7588
rect 21028 7644 21092 7648
rect 21028 7588 21032 7644
rect 21032 7588 21088 7644
rect 21088 7588 21092 7644
rect 21028 7584 21092 7588
rect 21108 7644 21172 7648
rect 21108 7588 21112 7644
rect 21112 7588 21168 7644
rect 21168 7588 21172 7644
rect 21108 7584 21172 7588
rect 21188 7644 21252 7648
rect 21188 7588 21192 7644
rect 21192 7588 21248 7644
rect 21248 7588 21252 7644
rect 21188 7584 21252 7588
rect 21268 7644 21332 7648
rect 21268 7588 21272 7644
rect 21272 7588 21328 7644
rect 21328 7588 21332 7644
rect 21268 7584 21332 7588
rect 27720 7644 27784 7648
rect 27720 7588 27724 7644
rect 27724 7588 27780 7644
rect 27780 7588 27784 7644
rect 27720 7584 27784 7588
rect 27800 7644 27864 7648
rect 27800 7588 27804 7644
rect 27804 7588 27860 7644
rect 27860 7588 27864 7644
rect 27800 7584 27864 7588
rect 27880 7644 27944 7648
rect 27880 7588 27884 7644
rect 27884 7588 27940 7644
rect 27940 7588 27944 7644
rect 27880 7584 27944 7588
rect 27960 7644 28024 7648
rect 27960 7588 27964 7644
rect 27964 7588 28020 7644
rect 28020 7588 28024 7644
rect 27960 7584 28024 7588
rect 4298 7100 4362 7104
rect 4298 7044 4302 7100
rect 4302 7044 4358 7100
rect 4358 7044 4362 7100
rect 4298 7040 4362 7044
rect 4378 7100 4442 7104
rect 4378 7044 4382 7100
rect 4382 7044 4438 7100
rect 4438 7044 4442 7100
rect 4378 7040 4442 7044
rect 4458 7100 4522 7104
rect 4458 7044 4462 7100
rect 4462 7044 4518 7100
rect 4518 7044 4522 7100
rect 4458 7040 4522 7044
rect 4538 7100 4602 7104
rect 4538 7044 4542 7100
rect 4542 7044 4598 7100
rect 4598 7044 4602 7100
rect 4538 7040 4602 7044
rect 10990 7100 11054 7104
rect 10990 7044 10994 7100
rect 10994 7044 11050 7100
rect 11050 7044 11054 7100
rect 10990 7040 11054 7044
rect 11070 7100 11134 7104
rect 11070 7044 11074 7100
rect 11074 7044 11130 7100
rect 11130 7044 11134 7100
rect 11070 7040 11134 7044
rect 11150 7100 11214 7104
rect 11150 7044 11154 7100
rect 11154 7044 11210 7100
rect 11210 7044 11214 7100
rect 11150 7040 11214 7044
rect 11230 7100 11294 7104
rect 11230 7044 11234 7100
rect 11234 7044 11290 7100
rect 11290 7044 11294 7100
rect 11230 7040 11294 7044
rect 17682 7100 17746 7104
rect 17682 7044 17686 7100
rect 17686 7044 17742 7100
rect 17742 7044 17746 7100
rect 17682 7040 17746 7044
rect 17762 7100 17826 7104
rect 17762 7044 17766 7100
rect 17766 7044 17822 7100
rect 17822 7044 17826 7100
rect 17762 7040 17826 7044
rect 17842 7100 17906 7104
rect 17842 7044 17846 7100
rect 17846 7044 17902 7100
rect 17902 7044 17906 7100
rect 17842 7040 17906 7044
rect 17922 7100 17986 7104
rect 17922 7044 17926 7100
rect 17926 7044 17982 7100
rect 17982 7044 17986 7100
rect 17922 7040 17986 7044
rect 24374 7100 24438 7104
rect 24374 7044 24378 7100
rect 24378 7044 24434 7100
rect 24434 7044 24438 7100
rect 24374 7040 24438 7044
rect 24454 7100 24518 7104
rect 24454 7044 24458 7100
rect 24458 7044 24514 7100
rect 24514 7044 24518 7100
rect 24454 7040 24518 7044
rect 24534 7100 24598 7104
rect 24534 7044 24538 7100
rect 24538 7044 24594 7100
rect 24594 7044 24598 7100
rect 24534 7040 24598 7044
rect 24614 7100 24678 7104
rect 24614 7044 24618 7100
rect 24618 7044 24674 7100
rect 24674 7044 24678 7100
rect 24614 7040 24678 7044
rect 7644 6556 7708 6560
rect 7644 6500 7648 6556
rect 7648 6500 7704 6556
rect 7704 6500 7708 6556
rect 7644 6496 7708 6500
rect 7724 6556 7788 6560
rect 7724 6500 7728 6556
rect 7728 6500 7784 6556
rect 7784 6500 7788 6556
rect 7724 6496 7788 6500
rect 7804 6556 7868 6560
rect 7804 6500 7808 6556
rect 7808 6500 7864 6556
rect 7864 6500 7868 6556
rect 7804 6496 7868 6500
rect 7884 6556 7948 6560
rect 7884 6500 7888 6556
rect 7888 6500 7944 6556
rect 7944 6500 7948 6556
rect 7884 6496 7948 6500
rect 14336 6556 14400 6560
rect 14336 6500 14340 6556
rect 14340 6500 14396 6556
rect 14396 6500 14400 6556
rect 14336 6496 14400 6500
rect 14416 6556 14480 6560
rect 14416 6500 14420 6556
rect 14420 6500 14476 6556
rect 14476 6500 14480 6556
rect 14416 6496 14480 6500
rect 14496 6556 14560 6560
rect 14496 6500 14500 6556
rect 14500 6500 14556 6556
rect 14556 6500 14560 6556
rect 14496 6496 14560 6500
rect 14576 6556 14640 6560
rect 14576 6500 14580 6556
rect 14580 6500 14636 6556
rect 14636 6500 14640 6556
rect 14576 6496 14640 6500
rect 21028 6556 21092 6560
rect 21028 6500 21032 6556
rect 21032 6500 21088 6556
rect 21088 6500 21092 6556
rect 21028 6496 21092 6500
rect 21108 6556 21172 6560
rect 21108 6500 21112 6556
rect 21112 6500 21168 6556
rect 21168 6500 21172 6556
rect 21108 6496 21172 6500
rect 21188 6556 21252 6560
rect 21188 6500 21192 6556
rect 21192 6500 21248 6556
rect 21248 6500 21252 6556
rect 21188 6496 21252 6500
rect 21268 6556 21332 6560
rect 21268 6500 21272 6556
rect 21272 6500 21328 6556
rect 21328 6500 21332 6556
rect 21268 6496 21332 6500
rect 27720 6556 27784 6560
rect 27720 6500 27724 6556
rect 27724 6500 27780 6556
rect 27780 6500 27784 6556
rect 27720 6496 27784 6500
rect 27800 6556 27864 6560
rect 27800 6500 27804 6556
rect 27804 6500 27860 6556
rect 27860 6500 27864 6556
rect 27800 6496 27864 6500
rect 27880 6556 27944 6560
rect 27880 6500 27884 6556
rect 27884 6500 27940 6556
rect 27940 6500 27944 6556
rect 27880 6496 27944 6500
rect 27960 6556 28024 6560
rect 27960 6500 27964 6556
rect 27964 6500 28020 6556
rect 28020 6500 28024 6556
rect 27960 6496 28024 6500
rect 4298 6012 4362 6016
rect 4298 5956 4302 6012
rect 4302 5956 4358 6012
rect 4358 5956 4362 6012
rect 4298 5952 4362 5956
rect 4378 6012 4442 6016
rect 4378 5956 4382 6012
rect 4382 5956 4438 6012
rect 4438 5956 4442 6012
rect 4378 5952 4442 5956
rect 4458 6012 4522 6016
rect 4458 5956 4462 6012
rect 4462 5956 4518 6012
rect 4518 5956 4522 6012
rect 4458 5952 4522 5956
rect 4538 6012 4602 6016
rect 4538 5956 4542 6012
rect 4542 5956 4598 6012
rect 4598 5956 4602 6012
rect 4538 5952 4602 5956
rect 10990 6012 11054 6016
rect 10990 5956 10994 6012
rect 10994 5956 11050 6012
rect 11050 5956 11054 6012
rect 10990 5952 11054 5956
rect 11070 6012 11134 6016
rect 11070 5956 11074 6012
rect 11074 5956 11130 6012
rect 11130 5956 11134 6012
rect 11070 5952 11134 5956
rect 11150 6012 11214 6016
rect 11150 5956 11154 6012
rect 11154 5956 11210 6012
rect 11210 5956 11214 6012
rect 11150 5952 11214 5956
rect 11230 6012 11294 6016
rect 11230 5956 11234 6012
rect 11234 5956 11290 6012
rect 11290 5956 11294 6012
rect 11230 5952 11294 5956
rect 17682 6012 17746 6016
rect 17682 5956 17686 6012
rect 17686 5956 17742 6012
rect 17742 5956 17746 6012
rect 17682 5952 17746 5956
rect 17762 6012 17826 6016
rect 17762 5956 17766 6012
rect 17766 5956 17822 6012
rect 17822 5956 17826 6012
rect 17762 5952 17826 5956
rect 17842 6012 17906 6016
rect 17842 5956 17846 6012
rect 17846 5956 17902 6012
rect 17902 5956 17906 6012
rect 17842 5952 17906 5956
rect 17922 6012 17986 6016
rect 17922 5956 17926 6012
rect 17926 5956 17982 6012
rect 17982 5956 17986 6012
rect 17922 5952 17986 5956
rect 24374 6012 24438 6016
rect 24374 5956 24378 6012
rect 24378 5956 24434 6012
rect 24434 5956 24438 6012
rect 24374 5952 24438 5956
rect 24454 6012 24518 6016
rect 24454 5956 24458 6012
rect 24458 5956 24514 6012
rect 24514 5956 24518 6012
rect 24454 5952 24518 5956
rect 24534 6012 24598 6016
rect 24534 5956 24538 6012
rect 24538 5956 24594 6012
rect 24594 5956 24598 6012
rect 24534 5952 24598 5956
rect 24614 6012 24678 6016
rect 24614 5956 24618 6012
rect 24618 5956 24674 6012
rect 24674 5956 24678 6012
rect 24614 5952 24678 5956
rect 7644 5468 7708 5472
rect 7644 5412 7648 5468
rect 7648 5412 7704 5468
rect 7704 5412 7708 5468
rect 7644 5408 7708 5412
rect 7724 5468 7788 5472
rect 7724 5412 7728 5468
rect 7728 5412 7784 5468
rect 7784 5412 7788 5468
rect 7724 5408 7788 5412
rect 7804 5468 7868 5472
rect 7804 5412 7808 5468
rect 7808 5412 7864 5468
rect 7864 5412 7868 5468
rect 7804 5408 7868 5412
rect 7884 5468 7948 5472
rect 7884 5412 7888 5468
rect 7888 5412 7944 5468
rect 7944 5412 7948 5468
rect 7884 5408 7948 5412
rect 14336 5468 14400 5472
rect 14336 5412 14340 5468
rect 14340 5412 14396 5468
rect 14396 5412 14400 5468
rect 14336 5408 14400 5412
rect 14416 5468 14480 5472
rect 14416 5412 14420 5468
rect 14420 5412 14476 5468
rect 14476 5412 14480 5468
rect 14416 5408 14480 5412
rect 14496 5468 14560 5472
rect 14496 5412 14500 5468
rect 14500 5412 14556 5468
rect 14556 5412 14560 5468
rect 14496 5408 14560 5412
rect 14576 5468 14640 5472
rect 14576 5412 14580 5468
rect 14580 5412 14636 5468
rect 14636 5412 14640 5468
rect 14576 5408 14640 5412
rect 21028 5468 21092 5472
rect 21028 5412 21032 5468
rect 21032 5412 21088 5468
rect 21088 5412 21092 5468
rect 21028 5408 21092 5412
rect 21108 5468 21172 5472
rect 21108 5412 21112 5468
rect 21112 5412 21168 5468
rect 21168 5412 21172 5468
rect 21108 5408 21172 5412
rect 21188 5468 21252 5472
rect 21188 5412 21192 5468
rect 21192 5412 21248 5468
rect 21248 5412 21252 5468
rect 21188 5408 21252 5412
rect 21268 5468 21332 5472
rect 21268 5412 21272 5468
rect 21272 5412 21328 5468
rect 21328 5412 21332 5468
rect 21268 5408 21332 5412
rect 27720 5468 27784 5472
rect 27720 5412 27724 5468
rect 27724 5412 27780 5468
rect 27780 5412 27784 5468
rect 27720 5408 27784 5412
rect 27800 5468 27864 5472
rect 27800 5412 27804 5468
rect 27804 5412 27860 5468
rect 27860 5412 27864 5468
rect 27800 5408 27864 5412
rect 27880 5468 27944 5472
rect 27880 5412 27884 5468
rect 27884 5412 27940 5468
rect 27940 5412 27944 5468
rect 27880 5408 27944 5412
rect 27960 5468 28024 5472
rect 27960 5412 27964 5468
rect 27964 5412 28020 5468
rect 28020 5412 28024 5468
rect 27960 5408 28024 5412
rect 4298 4924 4362 4928
rect 4298 4868 4302 4924
rect 4302 4868 4358 4924
rect 4358 4868 4362 4924
rect 4298 4864 4362 4868
rect 4378 4924 4442 4928
rect 4378 4868 4382 4924
rect 4382 4868 4438 4924
rect 4438 4868 4442 4924
rect 4378 4864 4442 4868
rect 4458 4924 4522 4928
rect 4458 4868 4462 4924
rect 4462 4868 4518 4924
rect 4518 4868 4522 4924
rect 4458 4864 4522 4868
rect 4538 4924 4602 4928
rect 4538 4868 4542 4924
rect 4542 4868 4598 4924
rect 4598 4868 4602 4924
rect 4538 4864 4602 4868
rect 10990 4924 11054 4928
rect 10990 4868 10994 4924
rect 10994 4868 11050 4924
rect 11050 4868 11054 4924
rect 10990 4864 11054 4868
rect 11070 4924 11134 4928
rect 11070 4868 11074 4924
rect 11074 4868 11130 4924
rect 11130 4868 11134 4924
rect 11070 4864 11134 4868
rect 11150 4924 11214 4928
rect 11150 4868 11154 4924
rect 11154 4868 11210 4924
rect 11210 4868 11214 4924
rect 11150 4864 11214 4868
rect 11230 4924 11294 4928
rect 11230 4868 11234 4924
rect 11234 4868 11290 4924
rect 11290 4868 11294 4924
rect 11230 4864 11294 4868
rect 17682 4924 17746 4928
rect 17682 4868 17686 4924
rect 17686 4868 17742 4924
rect 17742 4868 17746 4924
rect 17682 4864 17746 4868
rect 17762 4924 17826 4928
rect 17762 4868 17766 4924
rect 17766 4868 17822 4924
rect 17822 4868 17826 4924
rect 17762 4864 17826 4868
rect 17842 4924 17906 4928
rect 17842 4868 17846 4924
rect 17846 4868 17902 4924
rect 17902 4868 17906 4924
rect 17842 4864 17906 4868
rect 17922 4924 17986 4928
rect 17922 4868 17926 4924
rect 17926 4868 17982 4924
rect 17982 4868 17986 4924
rect 17922 4864 17986 4868
rect 24374 4924 24438 4928
rect 24374 4868 24378 4924
rect 24378 4868 24434 4924
rect 24434 4868 24438 4924
rect 24374 4864 24438 4868
rect 24454 4924 24518 4928
rect 24454 4868 24458 4924
rect 24458 4868 24514 4924
rect 24514 4868 24518 4924
rect 24454 4864 24518 4868
rect 24534 4924 24598 4928
rect 24534 4868 24538 4924
rect 24538 4868 24594 4924
rect 24594 4868 24598 4924
rect 24534 4864 24598 4868
rect 24614 4924 24678 4928
rect 24614 4868 24618 4924
rect 24618 4868 24674 4924
rect 24674 4868 24678 4924
rect 24614 4864 24678 4868
rect 7644 4380 7708 4384
rect 7644 4324 7648 4380
rect 7648 4324 7704 4380
rect 7704 4324 7708 4380
rect 7644 4320 7708 4324
rect 7724 4380 7788 4384
rect 7724 4324 7728 4380
rect 7728 4324 7784 4380
rect 7784 4324 7788 4380
rect 7724 4320 7788 4324
rect 7804 4380 7868 4384
rect 7804 4324 7808 4380
rect 7808 4324 7864 4380
rect 7864 4324 7868 4380
rect 7804 4320 7868 4324
rect 7884 4380 7948 4384
rect 7884 4324 7888 4380
rect 7888 4324 7944 4380
rect 7944 4324 7948 4380
rect 7884 4320 7948 4324
rect 14336 4380 14400 4384
rect 14336 4324 14340 4380
rect 14340 4324 14396 4380
rect 14396 4324 14400 4380
rect 14336 4320 14400 4324
rect 14416 4380 14480 4384
rect 14416 4324 14420 4380
rect 14420 4324 14476 4380
rect 14476 4324 14480 4380
rect 14416 4320 14480 4324
rect 14496 4380 14560 4384
rect 14496 4324 14500 4380
rect 14500 4324 14556 4380
rect 14556 4324 14560 4380
rect 14496 4320 14560 4324
rect 14576 4380 14640 4384
rect 14576 4324 14580 4380
rect 14580 4324 14636 4380
rect 14636 4324 14640 4380
rect 14576 4320 14640 4324
rect 21028 4380 21092 4384
rect 21028 4324 21032 4380
rect 21032 4324 21088 4380
rect 21088 4324 21092 4380
rect 21028 4320 21092 4324
rect 21108 4380 21172 4384
rect 21108 4324 21112 4380
rect 21112 4324 21168 4380
rect 21168 4324 21172 4380
rect 21108 4320 21172 4324
rect 21188 4380 21252 4384
rect 21188 4324 21192 4380
rect 21192 4324 21248 4380
rect 21248 4324 21252 4380
rect 21188 4320 21252 4324
rect 21268 4380 21332 4384
rect 21268 4324 21272 4380
rect 21272 4324 21328 4380
rect 21328 4324 21332 4380
rect 21268 4320 21332 4324
rect 27720 4380 27784 4384
rect 27720 4324 27724 4380
rect 27724 4324 27780 4380
rect 27780 4324 27784 4380
rect 27720 4320 27784 4324
rect 27800 4380 27864 4384
rect 27800 4324 27804 4380
rect 27804 4324 27860 4380
rect 27860 4324 27864 4380
rect 27800 4320 27864 4324
rect 27880 4380 27944 4384
rect 27880 4324 27884 4380
rect 27884 4324 27940 4380
rect 27940 4324 27944 4380
rect 27880 4320 27944 4324
rect 27960 4380 28024 4384
rect 27960 4324 27964 4380
rect 27964 4324 28020 4380
rect 28020 4324 28024 4380
rect 27960 4320 28024 4324
rect 4298 3836 4362 3840
rect 4298 3780 4302 3836
rect 4302 3780 4358 3836
rect 4358 3780 4362 3836
rect 4298 3776 4362 3780
rect 4378 3836 4442 3840
rect 4378 3780 4382 3836
rect 4382 3780 4438 3836
rect 4438 3780 4442 3836
rect 4378 3776 4442 3780
rect 4458 3836 4522 3840
rect 4458 3780 4462 3836
rect 4462 3780 4518 3836
rect 4518 3780 4522 3836
rect 4458 3776 4522 3780
rect 4538 3836 4602 3840
rect 4538 3780 4542 3836
rect 4542 3780 4598 3836
rect 4598 3780 4602 3836
rect 4538 3776 4602 3780
rect 10990 3836 11054 3840
rect 10990 3780 10994 3836
rect 10994 3780 11050 3836
rect 11050 3780 11054 3836
rect 10990 3776 11054 3780
rect 11070 3836 11134 3840
rect 11070 3780 11074 3836
rect 11074 3780 11130 3836
rect 11130 3780 11134 3836
rect 11070 3776 11134 3780
rect 11150 3836 11214 3840
rect 11150 3780 11154 3836
rect 11154 3780 11210 3836
rect 11210 3780 11214 3836
rect 11150 3776 11214 3780
rect 11230 3836 11294 3840
rect 11230 3780 11234 3836
rect 11234 3780 11290 3836
rect 11290 3780 11294 3836
rect 11230 3776 11294 3780
rect 17682 3836 17746 3840
rect 17682 3780 17686 3836
rect 17686 3780 17742 3836
rect 17742 3780 17746 3836
rect 17682 3776 17746 3780
rect 17762 3836 17826 3840
rect 17762 3780 17766 3836
rect 17766 3780 17822 3836
rect 17822 3780 17826 3836
rect 17762 3776 17826 3780
rect 17842 3836 17906 3840
rect 17842 3780 17846 3836
rect 17846 3780 17902 3836
rect 17902 3780 17906 3836
rect 17842 3776 17906 3780
rect 17922 3836 17986 3840
rect 17922 3780 17926 3836
rect 17926 3780 17982 3836
rect 17982 3780 17986 3836
rect 17922 3776 17986 3780
rect 24374 3836 24438 3840
rect 24374 3780 24378 3836
rect 24378 3780 24434 3836
rect 24434 3780 24438 3836
rect 24374 3776 24438 3780
rect 24454 3836 24518 3840
rect 24454 3780 24458 3836
rect 24458 3780 24514 3836
rect 24514 3780 24518 3836
rect 24454 3776 24518 3780
rect 24534 3836 24598 3840
rect 24534 3780 24538 3836
rect 24538 3780 24594 3836
rect 24594 3780 24598 3836
rect 24534 3776 24598 3780
rect 24614 3836 24678 3840
rect 24614 3780 24618 3836
rect 24618 3780 24674 3836
rect 24674 3780 24678 3836
rect 24614 3776 24678 3780
rect 7644 3292 7708 3296
rect 7644 3236 7648 3292
rect 7648 3236 7704 3292
rect 7704 3236 7708 3292
rect 7644 3232 7708 3236
rect 7724 3292 7788 3296
rect 7724 3236 7728 3292
rect 7728 3236 7784 3292
rect 7784 3236 7788 3292
rect 7724 3232 7788 3236
rect 7804 3292 7868 3296
rect 7804 3236 7808 3292
rect 7808 3236 7864 3292
rect 7864 3236 7868 3292
rect 7804 3232 7868 3236
rect 7884 3292 7948 3296
rect 7884 3236 7888 3292
rect 7888 3236 7944 3292
rect 7944 3236 7948 3292
rect 7884 3232 7948 3236
rect 14336 3292 14400 3296
rect 14336 3236 14340 3292
rect 14340 3236 14396 3292
rect 14396 3236 14400 3292
rect 14336 3232 14400 3236
rect 14416 3292 14480 3296
rect 14416 3236 14420 3292
rect 14420 3236 14476 3292
rect 14476 3236 14480 3292
rect 14416 3232 14480 3236
rect 14496 3292 14560 3296
rect 14496 3236 14500 3292
rect 14500 3236 14556 3292
rect 14556 3236 14560 3292
rect 14496 3232 14560 3236
rect 14576 3292 14640 3296
rect 14576 3236 14580 3292
rect 14580 3236 14636 3292
rect 14636 3236 14640 3292
rect 14576 3232 14640 3236
rect 21028 3292 21092 3296
rect 21028 3236 21032 3292
rect 21032 3236 21088 3292
rect 21088 3236 21092 3292
rect 21028 3232 21092 3236
rect 21108 3292 21172 3296
rect 21108 3236 21112 3292
rect 21112 3236 21168 3292
rect 21168 3236 21172 3292
rect 21108 3232 21172 3236
rect 21188 3292 21252 3296
rect 21188 3236 21192 3292
rect 21192 3236 21248 3292
rect 21248 3236 21252 3292
rect 21188 3232 21252 3236
rect 21268 3292 21332 3296
rect 21268 3236 21272 3292
rect 21272 3236 21328 3292
rect 21328 3236 21332 3292
rect 21268 3232 21332 3236
rect 27720 3292 27784 3296
rect 27720 3236 27724 3292
rect 27724 3236 27780 3292
rect 27780 3236 27784 3292
rect 27720 3232 27784 3236
rect 27800 3292 27864 3296
rect 27800 3236 27804 3292
rect 27804 3236 27860 3292
rect 27860 3236 27864 3292
rect 27800 3232 27864 3236
rect 27880 3292 27944 3296
rect 27880 3236 27884 3292
rect 27884 3236 27940 3292
rect 27940 3236 27944 3292
rect 27880 3232 27944 3236
rect 27960 3292 28024 3296
rect 27960 3236 27964 3292
rect 27964 3236 28020 3292
rect 28020 3236 28024 3292
rect 27960 3232 28024 3236
rect 4298 2748 4362 2752
rect 4298 2692 4302 2748
rect 4302 2692 4358 2748
rect 4358 2692 4362 2748
rect 4298 2688 4362 2692
rect 4378 2748 4442 2752
rect 4378 2692 4382 2748
rect 4382 2692 4438 2748
rect 4438 2692 4442 2748
rect 4378 2688 4442 2692
rect 4458 2748 4522 2752
rect 4458 2692 4462 2748
rect 4462 2692 4518 2748
rect 4518 2692 4522 2748
rect 4458 2688 4522 2692
rect 4538 2748 4602 2752
rect 4538 2692 4542 2748
rect 4542 2692 4598 2748
rect 4598 2692 4602 2748
rect 4538 2688 4602 2692
rect 10990 2748 11054 2752
rect 10990 2692 10994 2748
rect 10994 2692 11050 2748
rect 11050 2692 11054 2748
rect 10990 2688 11054 2692
rect 11070 2748 11134 2752
rect 11070 2692 11074 2748
rect 11074 2692 11130 2748
rect 11130 2692 11134 2748
rect 11070 2688 11134 2692
rect 11150 2748 11214 2752
rect 11150 2692 11154 2748
rect 11154 2692 11210 2748
rect 11210 2692 11214 2748
rect 11150 2688 11214 2692
rect 11230 2748 11294 2752
rect 11230 2692 11234 2748
rect 11234 2692 11290 2748
rect 11290 2692 11294 2748
rect 11230 2688 11294 2692
rect 17682 2748 17746 2752
rect 17682 2692 17686 2748
rect 17686 2692 17742 2748
rect 17742 2692 17746 2748
rect 17682 2688 17746 2692
rect 17762 2748 17826 2752
rect 17762 2692 17766 2748
rect 17766 2692 17822 2748
rect 17822 2692 17826 2748
rect 17762 2688 17826 2692
rect 17842 2748 17906 2752
rect 17842 2692 17846 2748
rect 17846 2692 17902 2748
rect 17902 2692 17906 2748
rect 17842 2688 17906 2692
rect 17922 2748 17986 2752
rect 17922 2692 17926 2748
rect 17926 2692 17982 2748
rect 17982 2692 17986 2748
rect 17922 2688 17986 2692
rect 24374 2748 24438 2752
rect 24374 2692 24378 2748
rect 24378 2692 24434 2748
rect 24434 2692 24438 2748
rect 24374 2688 24438 2692
rect 24454 2748 24518 2752
rect 24454 2692 24458 2748
rect 24458 2692 24514 2748
rect 24514 2692 24518 2748
rect 24454 2688 24518 2692
rect 24534 2748 24598 2752
rect 24534 2692 24538 2748
rect 24538 2692 24594 2748
rect 24594 2692 24598 2748
rect 24534 2688 24598 2692
rect 24614 2748 24678 2752
rect 24614 2692 24618 2748
rect 24618 2692 24674 2748
rect 24674 2692 24678 2748
rect 24614 2688 24678 2692
rect 7644 2204 7708 2208
rect 7644 2148 7648 2204
rect 7648 2148 7704 2204
rect 7704 2148 7708 2204
rect 7644 2144 7708 2148
rect 7724 2204 7788 2208
rect 7724 2148 7728 2204
rect 7728 2148 7784 2204
rect 7784 2148 7788 2204
rect 7724 2144 7788 2148
rect 7804 2204 7868 2208
rect 7804 2148 7808 2204
rect 7808 2148 7864 2204
rect 7864 2148 7868 2204
rect 7804 2144 7868 2148
rect 7884 2204 7948 2208
rect 7884 2148 7888 2204
rect 7888 2148 7944 2204
rect 7944 2148 7948 2204
rect 7884 2144 7948 2148
rect 14336 2204 14400 2208
rect 14336 2148 14340 2204
rect 14340 2148 14396 2204
rect 14396 2148 14400 2204
rect 14336 2144 14400 2148
rect 14416 2204 14480 2208
rect 14416 2148 14420 2204
rect 14420 2148 14476 2204
rect 14476 2148 14480 2204
rect 14416 2144 14480 2148
rect 14496 2204 14560 2208
rect 14496 2148 14500 2204
rect 14500 2148 14556 2204
rect 14556 2148 14560 2204
rect 14496 2144 14560 2148
rect 14576 2204 14640 2208
rect 14576 2148 14580 2204
rect 14580 2148 14636 2204
rect 14636 2148 14640 2204
rect 14576 2144 14640 2148
rect 21028 2204 21092 2208
rect 21028 2148 21032 2204
rect 21032 2148 21088 2204
rect 21088 2148 21092 2204
rect 21028 2144 21092 2148
rect 21108 2204 21172 2208
rect 21108 2148 21112 2204
rect 21112 2148 21168 2204
rect 21168 2148 21172 2204
rect 21108 2144 21172 2148
rect 21188 2204 21252 2208
rect 21188 2148 21192 2204
rect 21192 2148 21248 2204
rect 21248 2148 21252 2204
rect 21188 2144 21252 2148
rect 21268 2204 21332 2208
rect 21268 2148 21272 2204
rect 21272 2148 21328 2204
rect 21328 2148 21332 2204
rect 21268 2144 21332 2148
rect 27720 2204 27784 2208
rect 27720 2148 27724 2204
rect 27724 2148 27780 2204
rect 27780 2148 27784 2204
rect 27720 2144 27784 2148
rect 27800 2204 27864 2208
rect 27800 2148 27804 2204
rect 27804 2148 27860 2204
rect 27860 2148 27864 2204
rect 27800 2144 27864 2148
rect 27880 2204 27944 2208
rect 27880 2148 27884 2204
rect 27884 2148 27940 2204
rect 27940 2148 27944 2204
rect 27880 2144 27944 2148
rect 27960 2204 28024 2208
rect 27960 2148 27964 2204
rect 27964 2148 28020 2204
rect 28020 2148 28024 2204
rect 27960 2144 28024 2148
<< metal4 >>
rect 4290 26688 4610 26704
rect 4290 26624 4298 26688
rect 4362 26624 4378 26688
rect 4442 26624 4458 26688
rect 4522 26624 4538 26688
rect 4602 26624 4610 26688
rect 4290 25600 4610 26624
rect 4290 25536 4298 25600
rect 4362 25536 4378 25600
rect 4442 25536 4458 25600
rect 4522 25536 4538 25600
rect 4602 25536 4610 25600
rect 4290 24512 4610 25536
rect 4290 24448 4298 24512
rect 4362 24448 4378 24512
rect 4442 24448 4458 24512
rect 4522 24448 4538 24512
rect 4602 24448 4610 24512
rect 4290 23424 4610 24448
rect 4290 23360 4298 23424
rect 4362 23360 4378 23424
rect 4442 23360 4458 23424
rect 4522 23360 4538 23424
rect 4602 23360 4610 23424
rect 4290 22336 4610 23360
rect 4290 22272 4298 22336
rect 4362 22272 4378 22336
rect 4442 22272 4458 22336
rect 4522 22272 4538 22336
rect 4602 22272 4610 22336
rect 4290 21248 4610 22272
rect 4290 21184 4298 21248
rect 4362 21184 4378 21248
rect 4442 21184 4458 21248
rect 4522 21184 4538 21248
rect 4602 21184 4610 21248
rect 4290 20160 4610 21184
rect 4290 20096 4298 20160
rect 4362 20096 4378 20160
rect 4442 20096 4458 20160
rect 4522 20096 4538 20160
rect 4602 20096 4610 20160
rect 4290 19072 4610 20096
rect 4290 19008 4298 19072
rect 4362 19008 4378 19072
rect 4442 19008 4458 19072
rect 4522 19008 4538 19072
rect 4602 19008 4610 19072
rect 4290 17984 4610 19008
rect 4290 17920 4298 17984
rect 4362 17920 4378 17984
rect 4442 17920 4458 17984
rect 4522 17920 4538 17984
rect 4602 17920 4610 17984
rect 4290 16896 4610 17920
rect 4290 16832 4298 16896
rect 4362 16832 4378 16896
rect 4442 16832 4458 16896
rect 4522 16832 4538 16896
rect 4602 16832 4610 16896
rect 4290 15808 4610 16832
rect 4290 15744 4298 15808
rect 4362 15744 4378 15808
rect 4442 15744 4458 15808
rect 4522 15744 4538 15808
rect 4602 15744 4610 15808
rect 4290 14720 4610 15744
rect 4290 14656 4298 14720
rect 4362 14656 4378 14720
rect 4442 14656 4458 14720
rect 4522 14656 4538 14720
rect 4602 14656 4610 14720
rect 4290 13632 4610 14656
rect 4290 13568 4298 13632
rect 4362 13568 4378 13632
rect 4442 13568 4458 13632
rect 4522 13568 4538 13632
rect 4602 13568 4610 13632
rect 4290 12544 4610 13568
rect 4290 12480 4298 12544
rect 4362 12480 4378 12544
rect 4442 12480 4458 12544
rect 4522 12480 4538 12544
rect 4602 12480 4610 12544
rect 4290 11456 4610 12480
rect 4290 11392 4298 11456
rect 4362 11392 4378 11456
rect 4442 11392 4458 11456
rect 4522 11392 4538 11456
rect 4602 11392 4610 11456
rect 4290 10368 4610 11392
rect 4290 10304 4298 10368
rect 4362 10304 4378 10368
rect 4442 10304 4458 10368
rect 4522 10304 4538 10368
rect 4602 10304 4610 10368
rect 4290 9280 4610 10304
rect 4290 9216 4298 9280
rect 4362 9216 4378 9280
rect 4442 9216 4458 9280
rect 4522 9216 4538 9280
rect 4602 9216 4610 9280
rect 4290 8192 4610 9216
rect 4290 8128 4298 8192
rect 4362 8128 4378 8192
rect 4442 8128 4458 8192
rect 4522 8128 4538 8192
rect 4602 8128 4610 8192
rect 4290 7104 4610 8128
rect 4290 7040 4298 7104
rect 4362 7040 4378 7104
rect 4442 7040 4458 7104
rect 4522 7040 4538 7104
rect 4602 7040 4610 7104
rect 4290 6016 4610 7040
rect 4290 5952 4298 6016
rect 4362 5952 4378 6016
rect 4442 5952 4458 6016
rect 4522 5952 4538 6016
rect 4602 5952 4610 6016
rect 4290 4928 4610 5952
rect 4290 4864 4298 4928
rect 4362 4864 4378 4928
rect 4442 4864 4458 4928
rect 4522 4864 4538 4928
rect 4602 4864 4610 4928
rect 4290 3840 4610 4864
rect 4290 3776 4298 3840
rect 4362 3776 4378 3840
rect 4442 3776 4458 3840
rect 4522 3776 4538 3840
rect 4602 3776 4610 3840
rect 4290 2752 4610 3776
rect 4290 2688 4298 2752
rect 4362 2688 4378 2752
rect 4442 2688 4458 2752
rect 4522 2688 4538 2752
rect 4602 2688 4610 2752
rect 4290 2128 4610 2688
rect 7636 26144 7956 26704
rect 7636 26080 7644 26144
rect 7708 26080 7724 26144
rect 7788 26080 7804 26144
rect 7868 26080 7884 26144
rect 7948 26080 7956 26144
rect 7636 25056 7956 26080
rect 7636 24992 7644 25056
rect 7708 24992 7724 25056
rect 7788 24992 7804 25056
rect 7868 24992 7884 25056
rect 7948 24992 7956 25056
rect 7636 23968 7956 24992
rect 7636 23904 7644 23968
rect 7708 23904 7724 23968
rect 7788 23904 7804 23968
rect 7868 23904 7884 23968
rect 7948 23904 7956 23968
rect 7636 22880 7956 23904
rect 7636 22816 7644 22880
rect 7708 22816 7724 22880
rect 7788 22816 7804 22880
rect 7868 22816 7884 22880
rect 7948 22816 7956 22880
rect 7636 21792 7956 22816
rect 7636 21728 7644 21792
rect 7708 21728 7724 21792
rect 7788 21728 7804 21792
rect 7868 21728 7884 21792
rect 7948 21728 7956 21792
rect 7636 20704 7956 21728
rect 7636 20640 7644 20704
rect 7708 20640 7724 20704
rect 7788 20640 7804 20704
rect 7868 20640 7884 20704
rect 7948 20640 7956 20704
rect 7636 19616 7956 20640
rect 7636 19552 7644 19616
rect 7708 19552 7724 19616
rect 7788 19552 7804 19616
rect 7868 19552 7884 19616
rect 7948 19552 7956 19616
rect 7636 18528 7956 19552
rect 7636 18464 7644 18528
rect 7708 18464 7724 18528
rect 7788 18464 7804 18528
rect 7868 18464 7884 18528
rect 7948 18464 7956 18528
rect 7636 17440 7956 18464
rect 7636 17376 7644 17440
rect 7708 17376 7724 17440
rect 7788 17376 7804 17440
rect 7868 17376 7884 17440
rect 7948 17376 7956 17440
rect 7636 16352 7956 17376
rect 7636 16288 7644 16352
rect 7708 16288 7724 16352
rect 7788 16288 7804 16352
rect 7868 16288 7884 16352
rect 7948 16288 7956 16352
rect 7636 15264 7956 16288
rect 7636 15200 7644 15264
rect 7708 15200 7724 15264
rect 7788 15200 7804 15264
rect 7868 15200 7884 15264
rect 7948 15200 7956 15264
rect 7636 14176 7956 15200
rect 7636 14112 7644 14176
rect 7708 14112 7724 14176
rect 7788 14112 7804 14176
rect 7868 14112 7884 14176
rect 7948 14112 7956 14176
rect 7636 13088 7956 14112
rect 7636 13024 7644 13088
rect 7708 13024 7724 13088
rect 7788 13024 7804 13088
rect 7868 13024 7884 13088
rect 7948 13024 7956 13088
rect 7636 12000 7956 13024
rect 7636 11936 7644 12000
rect 7708 11936 7724 12000
rect 7788 11936 7804 12000
rect 7868 11936 7884 12000
rect 7948 11936 7956 12000
rect 7636 10912 7956 11936
rect 7636 10848 7644 10912
rect 7708 10848 7724 10912
rect 7788 10848 7804 10912
rect 7868 10848 7884 10912
rect 7948 10848 7956 10912
rect 7636 9824 7956 10848
rect 7636 9760 7644 9824
rect 7708 9760 7724 9824
rect 7788 9760 7804 9824
rect 7868 9760 7884 9824
rect 7948 9760 7956 9824
rect 7636 8736 7956 9760
rect 7636 8672 7644 8736
rect 7708 8672 7724 8736
rect 7788 8672 7804 8736
rect 7868 8672 7884 8736
rect 7948 8672 7956 8736
rect 7636 7648 7956 8672
rect 7636 7584 7644 7648
rect 7708 7584 7724 7648
rect 7788 7584 7804 7648
rect 7868 7584 7884 7648
rect 7948 7584 7956 7648
rect 7636 6560 7956 7584
rect 7636 6496 7644 6560
rect 7708 6496 7724 6560
rect 7788 6496 7804 6560
rect 7868 6496 7884 6560
rect 7948 6496 7956 6560
rect 7636 5472 7956 6496
rect 7636 5408 7644 5472
rect 7708 5408 7724 5472
rect 7788 5408 7804 5472
rect 7868 5408 7884 5472
rect 7948 5408 7956 5472
rect 7636 4384 7956 5408
rect 7636 4320 7644 4384
rect 7708 4320 7724 4384
rect 7788 4320 7804 4384
rect 7868 4320 7884 4384
rect 7948 4320 7956 4384
rect 7636 3296 7956 4320
rect 7636 3232 7644 3296
rect 7708 3232 7724 3296
rect 7788 3232 7804 3296
rect 7868 3232 7884 3296
rect 7948 3232 7956 3296
rect 7636 2208 7956 3232
rect 7636 2144 7644 2208
rect 7708 2144 7724 2208
rect 7788 2144 7804 2208
rect 7868 2144 7884 2208
rect 7948 2144 7956 2208
rect 7636 2128 7956 2144
rect 10982 26688 11302 26704
rect 10982 26624 10990 26688
rect 11054 26624 11070 26688
rect 11134 26624 11150 26688
rect 11214 26624 11230 26688
rect 11294 26624 11302 26688
rect 10982 25600 11302 26624
rect 10982 25536 10990 25600
rect 11054 25536 11070 25600
rect 11134 25536 11150 25600
rect 11214 25536 11230 25600
rect 11294 25536 11302 25600
rect 10982 24512 11302 25536
rect 10982 24448 10990 24512
rect 11054 24448 11070 24512
rect 11134 24448 11150 24512
rect 11214 24448 11230 24512
rect 11294 24448 11302 24512
rect 10982 23424 11302 24448
rect 10982 23360 10990 23424
rect 11054 23360 11070 23424
rect 11134 23360 11150 23424
rect 11214 23360 11230 23424
rect 11294 23360 11302 23424
rect 10982 22336 11302 23360
rect 10982 22272 10990 22336
rect 11054 22272 11070 22336
rect 11134 22272 11150 22336
rect 11214 22272 11230 22336
rect 11294 22272 11302 22336
rect 10982 21248 11302 22272
rect 10982 21184 10990 21248
rect 11054 21184 11070 21248
rect 11134 21184 11150 21248
rect 11214 21184 11230 21248
rect 11294 21184 11302 21248
rect 10982 20160 11302 21184
rect 10982 20096 10990 20160
rect 11054 20096 11070 20160
rect 11134 20096 11150 20160
rect 11214 20096 11230 20160
rect 11294 20096 11302 20160
rect 10982 19072 11302 20096
rect 10982 19008 10990 19072
rect 11054 19008 11070 19072
rect 11134 19008 11150 19072
rect 11214 19008 11230 19072
rect 11294 19008 11302 19072
rect 10982 17984 11302 19008
rect 10982 17920 10990 17984
rect 11054 17920 11070 17984
rect 11134 17920 11150 17984
rect 11214 17920 11230 17984
rect 11294 17920 11302 17984
rect 10982 16896 11302 17920
rect 10982 16832 10990 16896
rect 11054 16832 11070 16896
rect 11134 16832 11150 16896
rect 11214 16832 11230 16896
rect 11294 16832 11302 16896
rect 10982 15808 11302 16832
rect 10982 15744 10990 15808
rect 11054 15744 11070 15808
rect 11134 15744 11150 15808
rect 11214 15744 11230 15808
rect 11294 15744 11302 15808
rect 10982 14720 11302 15744
rect 10982 14656 10990 14720
rect 11054 14656 11070 14720
rect 11134 14656 11150 14720
rect 11214 14656 11230 14720
rect 11294 14656 11302 14720
rect 10982 13632 11302 14656
rect 10982 13568 10990 13632
rect 11054 13568 11070 13632
rect 11134 13568 11150 13632
rect 11214 13568 11230 13632
rect 11294 13568 11302 13632
rect 10982 12544 11302 13568
rect 10982 12480 10990 12544
rect 11054 12480 11070 12544
rect 11134 12480 11150 12544
rect 11214 12480 11230 12544
rect 11294 12480 11302 12544
rect 10982 11456 11302 12480
rect 10982 11392 10990 11456
rect 11054 11392 11070 11456
rect 11134 11392 11150 11456
rect 11214 11392 11230 11456
rect 11294 11392 11302 11456
rect 10982 10368 11302 11392
rect 10982 10304 10990 10368
rect 11054 10304 11070 10368
rect 11134 10304 11150 10368
rect 11214 10304 11230 10368
rect 11294 10304 11302 10368
rect 10982 9280 11302 10304
rect 10982 9216 10990 9280
rect 11054 9216 11070 9280
rect 11134 9216 11150 9280
rect 11214 9216 11230 9280
rect 11294 9216 11302 9280
rect 10982 8192 11302 9216
rect 10982 8128 10990 8192
rect 11054 8128 11070 8192
rect 11134 8128 11150 8192
rect 11214 8128 11230 8192
rect 11294 8128 11302 8192
rect 10982 7104 11302 8128
rect 10982 7040 10990 7104
rect 11054 7040 11070 7104
rect 11134 7040 11150 7104
rect 11214 7040 11230 7104
rect 11294 7040 11302 7104
rect 10982 6016 11302 7040
rect 10982 5952 10990 6016
rect 11054 5952 11070 6016
rect 11134 5952 11150 6016
rect 11214 5952 11230 6016
rect 11294 5952 11302 6016
rect 10982 4928 11302 5952
rect 10982 4864 10990 4928
rect 11054 4864 11070 4928
rect 11134 4864 11150 4928
rect 11214 4864 11230 4928
rect 11294 4864 11302 4928
rect 10982 3840 11302 4864
rect 10982 3776 10990 3840
rect 11054 3776 11070 3840
rect 11134 3776 11150 3840
rect 11214 3776 11230 3840
rect 11294 3776 11302 3840
rect 10982 2752 11302 3776
rect 10982 2688 10990 2752
rect 11054 2688 11070 2752
rect 11134 2688 11150 2752
rect 11214 2688 11230 2752
rect 11294 2688 11302 2752
rect 10982 2128 11302 2688
rect 14328 26144 14648 26704
rect 14328 26080 14336 26144
rect 14400 26080 14416 26144
rect 14480 26080 14496 26144
rect 14560 26080 14576 26144
rect 14640 26080 14648 26144
rect 14328 25056 14648 26080
rect 14328 24992 14336 25056
rect 14400 24992 14416 25056
rect 14480 24992 14496 25056
rect 14560 24992 14576 25056
rect 14640 24992 14648 25056
rect 14328 23968 14648 24992
rect 14328 23904 14336 23968
rect 14400 23904 14416 23968
rect 14480 23904 14496 23968
rect 14560 23904 14576 23968
rect 14640 23904 14648 23968
rect 14328 22880 14648 23904
rect 14328 22816 14336 22880
rect 14400 22816 14416 22880
rect 14480 22816 14496 22880
rect 14560 22816 14576 22880
rect 14640 22816 14648 22880
rect 14328 21792 14648 22816
rect 14328 21728 14336 21792
rect 14400 21728 14416 21792
rect 14480 21728 14496 21792
rect 14560 21728 14576 21792
rect 14640 21728 14648 21792
rect 14328 20704 14648 21728
rect 14328 20640 14336 20704
rect 14400 20640 14416 20704
rect 14480 20640 14496 20704
rect 14560 20640 14576 20704
rect 14640 20640 14648 20704
rect 14328 19616 14648 20640
rect 14328 19552 14336 19616
rect 14400 19552 14416 19616
rect 14480 19552 14496 19616
rect 14560 19552 14576 19616
rect 14640 19552 14648 19616
rect 14328 18528 14648 19552
rect 14328 18464 14336 18528
rect 14400 18464 14416 18528
rect 14480 18464 14496 18528
rect 14560 18464 14576 18528
rect 14640 18464 14648 18528
rect 14328 17440 14648 18464
rect 14328 17376 14336 17440
rect 14400 17376 14416 17440
rect 14480 17376 14496 17440
rect 14560 17376 14576 17440
rect 14640 17376 14648 17440
rect 14328 16352 14648 17376
rect 14328 16288 14336 16352
rect 14400 16288 14416 16352
rect 14480 16288 14496 16352
rect 14560 16288 14576 16352
rect 14640 16288 14648 16352
rect 14328 15264 14648 16288
rect 14328 15200 14336 15264
rect 14400 15200 14416 15264
rect 14480 15200 14496 15264
rect 14560 15200 14576 15264
rect 14640 15200 14648 15264
rect 14328 14176 14648 15200
rect 14328 14112 14336 14176
rect 14400 14112 14416 14176
rect 14480 14112 14496 14176
rect 14560 14112 14576 14176
rect 14640 14112 14648 14176
rect 14328 13088 14648 14112
rect 14328 13024 14336 13088
rect 14400 13024 14416 13088
rect 14480 13024 14496 13088
rect 14560 13024 14576 13088
rect 14640 13024 14648 13088
rect 14328 12000 14648 13024
rect 14328 11936 14336 12000
rect 14400 11936 14416 12000
rect 14480 11936 14496 12000
rect 14560 11936 14576 12000
rect 14640 11936 14648 12000
rect 14328 10912 14648 11936
rect 14328 10848 14336 10912
rect 14400 10848 14416 10912
rect 14480 10848 14496 10912
rect 14560 10848 14576 10912
rect 14640 10848 14648 10912
rect 14328 9824 14648 10848
rect 14328 9760 14336 9824
rect 14400 9760 14416 9824
rect 14480 9760 14496 9824
rect 14560 9760 14576 9824
rect 14640 9760 14648 9824
rect 14328 8736 14648 9760
rect 14328 8672 14336 8736
rect 14400 8672 14416 8736
rect 14480 8672 14496 8736
rect 14560 8672 14576 8736
rect 14640 8672 14648 8736
rect 14328 7648 14648 8672
rect 14328 7584 14336 7648
rect 14400 7584 14416 7648
rect 14480 7584 14496 7648
rect 14560 7584 14576 7648
rect 14640 7584 14648 7648
rect 14328 6560 14648 7584
rect 14328 6496 14336 6560
rect 14400 6496 14416 6560
rect 14480 6496 14496 6560
rect 14560 6496 14576 6560
rect 14640 6496 14648 6560
rect 14328 5472 14648 6496
rect 14328 5408 14336 5472
rect 14400 5408 14416 5472
rect 14480 5408 14496 5472
rect 14560 5408 14576 5472
rect 14640 5408 14648 5472
rect 14328 4384 14648 5408
rect 14328 4320 14336 4384
rect 14400 4320 14416 4384
rect 14480 4320 14496 4384
rect 14560 4320 14576 4384
rect 14640 4320 14648 4384
rect 14328 3296 14648 4320
rect 14328 3232 14336 3296
rect 14400 3232 14416 3296
rect 14480 3232 14496 3296
rect 14560 3232 14576 3296
rect 14640 3232 14648 3296
rect 14328 2208 14648 3232
rect 14328 2144 14336 2208
rect 14400 2144 14416 2208
rect 14480 2144 14496 2208
rect 14560 2144 14576 2208
rect 14640 2144 14648 2208
rect 14328 2128 14648 2144
rect 17674 26688 17994 26704
rect 17674 26624 17682 26688
rect 17746 26624 17762 26688
rect 17826 26624 17842 26688
rect 17906 26624 17922 26688
rect 17986 26624 17994 26688
rect 17674 25600 17994 26624
rect 17674 25536 17682 25600
rect 17746 25536 17762 25600
rect 17826 25536 17842 25600
rect 17906 25536 17922 25600
rect 17986 25536 17994 25600
rect 17674 24512 17994 25536
rect 17674 24448 17682 24512
rect 17746 24448 17762 24512
rect 17826 24448 17842 24512
rect 17906 24448 17922 24512
rect 17986 24448 17994 24512
rect 17674 23424 17994 24448
rect 17674 23360 17682 23424
rect 17746 23360 17762 23424
rect 17826 23360 17842 23424
rect 17906 23360 17922 23424
rect 17986 23360 17994 23424
rect 17674 22336 17994 23360
rect 17674 22272 17682 22336
rect 17746 22272 17762 22336
rect 17826 22272 17842 22336
rect 17906 22272 17922 22336
rect 17986 22272 17994 22336
rect 17674 21248 17994 22272
rect 17674 21184 17682 21248
rect 17746 21184 17762 21248
rect 17826 21184 17842 21248
rect 17906 21184 17922 21248
rect 17986 21184 17994 21248
rect 17674 20160 17994 21184
rect 17674 20096 17682 20160
rect 17746 20096 17762 20160
rect 17826 20096 17842 20160
rect 17906 20096 17922 20160
rect 17986 20096 17994 20160
rect 17674 19072 17994 20096
rect 17674 19008 17682 19072
rect 17746 19008 17762 19072
rect 17826 19008 17842 19072
rect 17906 19008 17922 19072
rect 17986 19008 17994 19072
rect 17674 17984 17994 19008
rect 17674 17920 17682 17984
rect 17746 17920 17762 17984
rect 17826 17920 17842 17984
rect 17906 17920 17922 17984
rect 17986 17920 17994 17984
rect 17674 16896 17994 17920
rect 17674 16832 17682 16896
rect 17746 16832 17762 16896
rect 17826 16832 17842 16896
rect 17906 16832 17922 16896
rect 17986 16832 17994 16896
rect 17674 15808 17994 16832
rect 17674 15744 17682 15808
rect 17746 15744 17762 15808
rect 17826 15744 17842 15808
rect 17906 15744 17922 15808
rect 17986 15744 17994 15808
rect 17674 14720 17994 15744
rect 17674 14656 17682 14720
rect 17746 14656 17762 14720
rect 17826 14656 17842 14720
rect 17906 14656 17922 14720
rect 17986 14656 17994 14720
rect 17674 13632 17994 14656
rect 17674 13568 17682 13632
rect 17746 13568 17762 13632
rect 17826 13568 17842 13632
rect 17906 13568 17922 13632
rect 17986 13568 17994 13632
rect 17674 12544 17994 13568
rect 17674 12480 17682 12544
rect 17746 12480 17762 12544
rect 17826 12480 17842 12544
rect 17906 12480 17922 12544
rect 17986 12480 17994 12544
rect 17674 11456 17994 12480
rect 17674 11392 17682 11456
rect 17746 11392 17762 11456
rect 17826 11392 17842 11456
rect 17906 11392 17922 11456
rect 17986 11392 17994 11456
rect 17674 10368 17994 11392
rect 17674 10304 17682 10368
rect 17746 10304 17762 10368
rect 17826 10304 17842 10368
rect 17906 10304 17922 10368
rect 17986 10304 17994 10368
rect 17674 9280 17994 10304
rect 17674 9216 17682 9280
rect 17746 9216 17762 9280
rect 17826 9216 17842 9280
rect 17906 9216 17922 9280
rect 17986 9216 17994 9280
rect 17674 8192 17994 9216
rect 17674 8128 17682 8192
rect 17746 8128 17762 8192
rect 17826 8128 17842 8192
rect 17906 8128 17922 8192
rect 17986 8128 17994 8192
rect 17674 7104 17994 8128
rect 17674 7040 17682 7104
rect 17746 7040 17762 7104
rect 17826 7040 17842 7104
rect 17906 7040 17922 7104
rect 17986 7040 17994 7104
rect 17674 6016 17994 7040
rect 17674 5952 17682 6016
rect 17746 5952 17762 6016
rect 17826 5952 17842 6016
rect 17906 5952 17922 6016
rect 17986 5952 17994 6016
rect 17674 4928 17994 5952
rect 17674 4864 17682 4928
rect 17746 4864 17762 4928
rect 17826 4864 17842 4928
rect 17906 4864 17922 4928
rect 17986 4864 17994 4928
rect 17674 3840 17994 4864
rect 17674 3776 17682 3840
rect 17746 3776 17762 3840
rect 17826 3776 17842 3840
rect 17906 3776 17922 3840
rect 17986 3776 17994 3840
rect 17674 2752 17994 3776
rect 17674 2688 17682 2752
rect 17746 2688 17762 2752
rect 17826 2688 17842 2752
rect 17906 2688 17922 2752
rect 17986 2688 17994 2752
rect 17674 2128 17994 2688
rect 21020 26144 21340 26704
rect 21020 26080 21028 26144
rect 21092 26080 21108 26144
rect 21172 26080 21188 26144
rect 21252 26080 21268 26144
rect 21332 26080 21340 26144
rect 21020 25056 21340 26080
rect 21020 24992 21028 25056
rect 21092 24992 21108 25056
rect 21172 24992 21188 25056
rect 21252 24992 21268 25056
rect 21332 24992 21340 25056
rect 21020 23968 21340 24992
rect 21020 23904 21028 23968
rect 21092 23904 21108 23968
rect 21172 23904 21188 23968
rect 21252 23904 21268 23968
rect 21332 23904 21340 23968
rect 21020 22880 21340 23904
rect 21020 22816 21028 22880
rect 21092 22816 21108 22880
rect 21172 22816 21188 22880
rect 21252 22816 21268 22880
rect 21332 22816 21340 22880
rect 21020 21792 21340 22816
rect 21020 21728 21028 21792
rect 21092 21728 21108 21792
rect 21172 21728 21188 21792
rect 21252 21728 21268 21792
rect 21332 21728 21340 21792
rect 21020 20704 21340 21728
rect 21020 20640 21028 20704
rect 21092 20640 21108 20704
rect 21172 20640 21188 20704
rect 21252 20640 21268 20704
rect 21332 20640 21340 20704
rect 21020 19616 21340 20640
rect 21020 19552 21028 19616
rect 21092 19552 21108 19616
rect 21172 19552 21188 19616
rect 21252 19552 21268 19616
rect 21332 19552 21340 19616
rect 21020 18528 21340 19552
rect 21020 18464 21028 18528
rect 21092 18464 21108 18528
rect 21172 18464 21188 18528
rect 21252 18464 21268 18528
rect 21332 18464 21340 18528
rect 21020 17440 21340 18464
rect 21020 17376 21028 17440
rect 21092 17376 21108 17440
rect 21172 17376 21188 17440
rect 21252 17376 21268 17440
rect 21332 17376 21340 17440
rect 21020 16352 21340 17376
rect 21020 16288 21028 16352
rect 21092 16288 21108 16352
rect 21172 16288 21188 16352
rect 21252 16288 21268 16352
rect 21332 16288 21340 16352
rect 21020 15264 21340 16288
rect 21020 15200 21028 15264
rect 21092 15200 21108 15264
rect 21172 15200 21188 15264
rect 21252 15200 21268 15264
rect 21332 15200 21340 15264
rect 21020 14176 21340 15200
rect 21020 14112 21028 14176
rect 21092 14112 21108 14176
rect 21172 14112 21188 14176
rect 21252 14112 21268 14176
rect 21332 14112 21340 14176
rect 21020 13088 21340 14112
rect 21020 13024 21028 13088
rect 21092 13024 21108 13088
rect 21172 13024 21188 13088
rect 21252 13024 21268 13088
rect 21332 13024 21340 13088
rect 21020 12000 21340 13024
rect 21020 11936 21028 12000
rect 21092 11936 21108 12000
rect 21172 11936 21188 12000
rect 21252 11936 21268 12000
rect 21332 11936 21340 12000
rect 21020 10912 21340 11936
rect 21020 10848 21028 10912
rect 21092 10848 21108 10912
rect 21172 10848 21188 10912
rect 21252 10848 21268 10912
rect 21332 10848 21340 10912
rect 21020 9824 21340 10848
rect 21020 9760 21028 9824
rect 21092 9760 21108 9824
rect 21172 9760 21188 9824
rect 21252 9760 21268 9824
rect 21332 9760 21340 9824
rect 21020 8736 21340 9760
rect 21020 8672 21028 8736
rect 21092 8672 21108 8736
rect 21172 8672 21188 8736
rect 21252 8672 21268 8736
rect 21332 8672 21340 8736
rect 21020 7648 21340 8672
rect 21020 7584 21028 7648
rect 21092 7584 21108 7648
rect 21172 7584 21188 7648
rect 21252 7584 21268 7648
rect 21332 7584 21340 7648
rect 21020 6560 21340 7584
rect 21020 6496 21028 6560
rect 21092 6496 21108 6560
rect 21172 6496 21188 6560
rect 21252 6496 21268 6560
rect 21332 6496 21340 6560
rect 21020 5472 21340 6496
rect 21020 5408 21028 5472
rect 21092 5408 21108 5472
rect 21172 5408 21188 5472
rect 21252 5408 21268 5472
rect 21332 5408 21340 5472
rect 21020 4384 21340 5408
rect 21020 4320 21028 4384
rect 21092 4320 21108 4384
rect 21172 4320 21188 4384
rect 21252 4320 21268 4384
rect 21332 4320 21340 4384
rect 21020 3296 21340 4320
rect 21020 3232 21028 3296
rect 21092 3232 21108 3296
rect 21172 3232 21188 3296
rect 21252 3232 21268 3296
rect 21332 3232 21340 3296
rect 21020 2208 21340 3232
rect 21020 2144 21028 2208
rect 21092 2144 21108 2208
rect 21172 2144 21188 2208
rect 21252 2144 21268 2208
rect 21332 2144 21340 2208
rect 21020 2128 21340 2144
rect 24366 26688 24686 26704
rect 24366 26624 24374 26688
rect 24438 26624 24454 26688
rect 24518 26624 24534 26688
rect 24598 26624 24614 26688
rect 24678 26624 24686 26688
rect 24366 25600 24686 26624
rect 24366 25536 24374 25600
rect 24438 25536 24454 25600
rect 24518 25536 24534 25600
rect 24598 25536 24614 25600
rect 24678 25536 24686 25600
rect 24366 24512 24686 25536
rect 24366 24448 24374 24512
rect 24438 24448 24454 24512
rect 24518 24448 24534 24512
rect 24598 24448 24614 24512
rect 24678 24448 24686 24512
rect 24366 23424 24686 24448
rect 24366 23360 24374 23424
rect 24438 23360 24454 23424
rect 24518 23360 24534 23424
rect 24598 23360 24614 23424
rect 24678 23360 24686 23424
rect 24366 22336 24686 23360
rect 24366 22272 24374 22336
rect 24438 22272 24454 22336
rect 24518 22272 24534 22336
rect 24598 22272 24614 22336
rect 24678 22272 24686 22336
rect 24366 21248 24686 22272
rect 24366 21184 24374 21248
rect 24438 21184 24454 21248
rect 24518 21184 24534 21248
rect 24598 21184 24614 21248
rect 24678 21184 24686 21248
rect 24366 20160 24686 21184
rect 24366 20096 24374 20160
rect 24438 20096 24454 20160
rect 24518 20096 24534 20160
rect 24598 20096 24614 20160
rect 24678 20096 24686 20160
rect 24366 19072 24686 20096
rect 24366 19008 24374 19072
rect 24438 19008 24454 19072
rect 24518 19008 24534 19072
rect 24598 19008 24614 19072
rect 24678 19008 24686 19072
rect 24366 17984 24686 19008
rect 24366 17920 24374 17984
rect 24438 17920 24454 17984
rect 24518 17920 24534 17984
rect 24598 17920 24614 17984
rect 24678 17920 24686 17984
rect 24366 16896 24686 17920
rect 24366 16832 24374 16896
rect 24438 16832 24454 16896
rect 24518 16832 24534 16896
rect 24598 16832 24614 16896
rect 24678 16832 24686 16896
rect 24366 15808 24686 16832
rect 24366 15744 24374 15808
rect 24438 15744 24454 15808
rect 24518 15744 24534 15808
rect 24598 15744 24614 15808
rect 24678 15744 24686 15808
rect 24366 14720 24686 15744
rect 24366 14656 24374 14720
rect 24438 14656 24454 14720
rect 24518 14656 24534 14720
rect 24598 14656 24614 14720
rect 24678 14656 24686 14720
rect 24366 13632 24686 14656
rect 24366 13568 24374 13632
rect 24438 13568 24454 13632
rect 24518 13568 24534 13632
rect 24598 13568 24614 13632
rect 24678 13568 24686 13632
rect 24366 12544 24686 13568
rect 24366 12480 24374 12544
rect 24438 12480 24454 12544
rect 24518 12480 24534 12544
rect 24598 12480 24614 12544
rect 24678 12480 24686 12544
rect 24366 11456 24686 12480
rect 24366 11392 24374 11456
rect 24438 11392 24454 11456
rect 24518 11392 24534 11456
rect 24598 11392 24614 11456
rect 24678 11392 24686 11456
rect 24366 10368 24686 11392
rect 24366 10304 24374 10368
rect 24438 10304 24454 10368
rect 24518 10304 24534 10368
rect 24598 10304 24614 10368
rect 24678 10304 24686 10368
rect 24366 9280 24686 10304
rect 24366 9216 24374 9280
rect 24438 9216 24454 9280
rect 24518 9216 24534 9280
rect 24598 9216 24614 9280
rect 24678 9216 24686 9280
rect 24366 8192 24686 9216
rect 24366 8128 24374 8192
rect 24438 8128 24454 8192
rect 24518 8128 24534 8192
rect 24598 8128 24614 8192
rect 24678 8128 24686 8192
rect 24366 7104 24686 8128
rect 24366 7040 24374 7104
rect 24438 7040 24454 7104
rect 24518 7040 24534 7104
rect 24598 7040 24614 7104
rect 24678 7040 24686 7104
rect 24366 6016 24686 7040
rect 24366 5952 24374 6016
rect 24438 5952 24454 6016
rect 24518 5952 24534 6016
rect 24598 5952 24614 6016
rect 24678 5952 24686 6016
rect 24366 4928 24686 5952
rect 24366 4864 24374 4928
rect 24438 4864 24454 4928
rect 24518 4864 24534 4928
rect 24598 4864 24614 4928
rect 24678 4864 24686 4928
rect 24366 3840 24686 4864
rect 24366 3776 24374 3840
rect 24438 3776 24454 3840
rect 24518 3776 24534 3840
rect 24598 3776 24614 3840
rect 24678 3776 24686 3840
rect 24366 2752 24686 3776
rect 24366 2688 24374 2752
rect 24438 2688 24454 2752
rect 24518 2688 24534 2752
rect 24598 2688 24614 2752
rect 24678 2688 24686 2752
rect 24366 2128 24686 2688
rect 27712 26144 28032 26704
rect 27712 26080 27720 26144
rect 27784 26080 27800 26144
rect 27864 26080 27880 26144
rect 27944 26080 27960 26144
rect 28024 26080 28032 26144
rect 27712 25056 28032 26080
rect 27712 24992 27720 25056
rect 27784 24992 27800 25056
rect 27864 24992 27880 25056
rect 27944 24992 27960 25056
rect 28024 24992 28032 25056
rect 27712 23968 28032 24992
rect 27712 23904 27720 23968
rect 27784 23904 27800 23968
rect 27864 23904 27880 23968
rect 27944 23904 27960 23968
rect 28024 23904 28032 23968
rect 27712 22880 28032 23904
rect 27712 22816 27720 22880
rect 27784 22816 27800 22880
rect 27864 22816 27880 22880
rect 27944 22816 27960 22880
rect 28024 22816 28032 22880
rect 27712 21792 28032 22816
rect 27712 21728 27720 21792
rect 27784 21728 27800 21792
rect 27864 21728 27880 21792
rect 27944 21728 27960 21792
rect 28024 21728 28032 21792
rect 27712 20704 28032 21728
rect 27712 20640 27720 20704
rect 27784 20640 27800 20704
rect 27864 20640 27880 20704
rect 27944 20640 27960 20704
rect 28024 20640 28032 20704
rect 27712 19616 28032 20640
rect 27712 19552 27720 19616
rect 27784 19552 27800 19616
rect 27864 19552 27880 19616
rect 27944 19552 27960 19616
rect 28024 19552 28032 19616
rect 27712 18528 28032 19552
rect 27712 18464 27720 18528
rect 27784 18464 27800 18528
rect 27864 18464 27880 18528
rect 27944 18464 27960 18528
rect 28024 18464 28032 18528
rect 27712 17440 28032 18464
rect 27712 17376 27720 17440
rect 27784 17376 27800 17440
rect 27864 17376 27880 17440
rect 27944 17376 27960 17440
rect 28024 17376 28032 17440
rect 27712 16352 28032 17376
rect 27712 16288 27720 16352
rect 27784 16288 27800 16352
rect 27864 16288 27880 16352
rect 27944 16288 27960 16352
rect 28024 16288 28032 16352
rect 27712 15264 28032 16288
rect 27712 15200 27720 15264
rect 27784 15200 27800 15264
rect 27864 15200 27880 15264
rect 27944 15200 27960 15264
rect 28024 15200 28032 15264
rect 27712 14176 28032 15200
rect 27712 14112 27720 14176
rect 27784 14112 27800 14176
rect 27864 14112 27880 14176
rect 27944 14112 27960 14176
rect 28024 14112 28032 14176
rect 27712 13088 28032 14112
rect 27712 13024 27720 13088
rect 27784 13024 27800 13088
rect 27864 13024 27880 13088
rect 27944 13024 27960 13088
rect 28024 13024 28032 13088
rect 27712 12000 28032 13024
rect 27712 11936 27720 12000
rect 27784 11936 27800 12000
rect 27864 11936 27880 12000
rect 27944 11936 27960 12000
rect 28024 11936 28032 12000
rect 27712 10912 28032 11936
rect 27712 10848 27720 10912
rect 27784 10848 27800 10912
rect 27864 10848 27880 10912
rect 27944 10848 27960 10912
rect 28024 10848 28032 10912
rect 27712 9824 28032 10848
rect 27712 9760 27720 9824
rect 27784 9760 27800 9824
rect 27864 9760 27880 9824
rect 27944 9760 27960 9824
rect 28024 9760 28032 9824
rect 27712 8736 28032 9760
rect 27712 8672 27720 8736
rect 27784 8672 27800 8736
rect 27864 8672 27880 8736
rect 27944 8672 27960 8736
rect 28024 8672 28032 8736
rect 27712 7648 28032 8672
rect 27712 7584 27720 7648
rect 27784 7584 27800 7648
rect 27864 7584 27880 7648
rect 27944 7584 27960 7648
rect 28024 7584 28032 7648
rect 27712 6560 28032 7584
rect 27712 6496 27720 6560
rect 27784 6496 27800 6560
rect 27864 6496 27880 6560
rect 27944 6496 27960 6560
rect 28024 6496 28032 6560
rect 27712 5472 28032 6496
rect 27712 5408 27720 5472
rect 27784 5408 27800 5472
rect 27864 5408 27880 5472
rect 27944 5408 27960 5472
rect 28024 5408 28032 5472
rect 27712 4384 28032 5408
rect 27712 4320 27720 4384
rect 27784 4320 27800 4384
rect 27864 4320 27880 4384
rect 27944 4320 27960 4384
rect 28024 4320 28032 4384
rect 27712 3296 28032 4320
rect 27712 3232 27720 3296
rect 27784 3232 27800 3296
rect 27864 3232 27880 3296
rect 27944 3232 27960 3296
rect 28024 3232 28032 3296
rect 27712 2208 28032 3232
rect 27712 2144 27720 2208
rect 27784 2144 27800 2208
rect 27864 2144 27880 2208
rect 27944 2144 27960 2208
rect 28024 2144 28032 2208
rect 27712 2128 28032 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__389__B $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6992 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__B
timestamp 1666464484
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A0
timestamp 1666464484
transform 1 0 4968 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A0
timestamp 1666464484
transform -1 0 8188 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1666464484
transform -1 0 13156 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A0
timestamp 1666464484
transform -1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1666464484
transform -1 0 24012 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A0
timestamp 1666464484
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1666464484
transform -1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__C1
timestamp 1666464484
transform -1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__C1
timestamp 1666464484
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1666464484
transform 1 0 14996 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1666464484
transform 1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1666464484
transform 1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1666464484
transform -1 0 11868 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1666464484
transform 1 0 10488 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1666464484
transform 1 0 20976 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__C
timestamp 1666464484
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__A
timestamp 1666464484
transform -1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A
timestamp 1666464484
transform -1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1666464484
transform -1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__D
timestamp 1666464484
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__A
timestamp 1666464484
transform 1 0 23828 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A
timestamp 1666464484
transform -1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__A
timestamp 1666464484
transform 1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__A
timestamp 1666464484
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__A
timestamp 1666464484
transform -1 0 26312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__A
timestamp 1666464484
transform -1 0 26312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__A
timestamp 1666464484
transform 1 0 22264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__A
timestamp 1666464484
transform -1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__A
timestamp 1666464484
transform -1 0 27324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A
timestamp 1666464484
transform -1 0 27324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A
timestamp 1666464484
transform -1 0 27324 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1666464484
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__B
timestamp 1666464484
transform -1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A0
timestamp 1666464484
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__A0
timestamp 1666464484
transform -1 0 25484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__A0
timestamp 1666464484
transform 1 0 23460 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__B
timestamp 1666464484
transform 1 0 6900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__B1
timestamp 1666464484
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__A
timestamp 1666464484
transform -1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__A
timestamp 1666464484
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__A
timestamp 1666464484
transform -1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__651__A
timestamp 1666464484
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__A
timestamp 1666464484
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__656__B1
timestamp 1666464484
transform -1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__B
timestamp 1666464484
transform 1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__B
timestamp 1666464484
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__B
timestamp 1666464484
transform -1 0 4416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__B
timestamp 1666464484
transform 1 0 4416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__B
timestamp 1666464484
transform 1 0 6624 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__B
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__B
timestamp 1666464484
transform 1 0 3128 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__B
timestamp 1666464484
transform -1 0 5336 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__A0
timestamp 1666464484
transform -1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__A0
timestamp 1666464484
transform 1 0 23552 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__673__A0
timestamp 1666464484
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__A0
timestamp 1666464484
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__D
timestamp 1666464484
transform 1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__A0
timestamp 1666464484
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__A0
timestamp 1666464484
transform 1 0 23736 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__A0
timestamp 1666464484
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__685__A0
timestamp 1666464484
transform -1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__A
timestamp 1666464484
transform -1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__A0
timestamp 1666464484
transform -1 0 8096 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__690__A0
timestamp 1666464484
transform -1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__692__A0
timestamp 1666464484
transform -1 0 6992 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__694__A0
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__A
timestamp 1666464484
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__711__A
timestamp 1666464484
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__722__A0
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__724__A0
timestamp 1666464484
transform -1 0 19688 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__726__A0
timestamp 1666464484
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__728__A0
timestamp 1666464484
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__730__A0
timestamp 1666464484
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__732__A0
timestamp 1666464484
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__734__A0
timestamp 1666464484
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__737__A0
timestamp 1666464484
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__739__A0
timestamp 1666464484
transform 1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__741__A0
timestamp 1666464484
transform -1 0 19596 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__743__A0
timestamp 1666464484
transform 1 0 19964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__749__A
timestamp 1666464484
transform -1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__757__A0
timestamp 1666464484
transform -1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__759__A0
timestamp 1666464484
transform 1 0 24104 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__761__A0
timestamp 1666464484
transform -1 0 24840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__764__A0
timestamp 1666464484
transform -1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__766__A0
timestamp 1666464484
transform -1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__768__A0
timestamp 1666464484
transform -1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__770__A0
timestamp 1666464484
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__773__A0
timestamp 1666464484
transform -1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__775__A0
timestamp 1666464484
transform -1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__777__A0
timestamp 1666464484
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__779__A0
timestamp 1666464484
transform -1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__785__A
timestamp 1666464484
transform -1 0 13156 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__793__A0
timestamp 1666464484
transform -1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__795__A0
timestamp 1666464484
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__797__A0
timestamp 1666464484
transform -1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__800__A0
timestamp 1666464484
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__802__A0
timestamp 1666464484
transform 1 0 9568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__804__A0
timestamp 1666464484
transform 1 0 9476 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__806__A0
timestamp 1666464484
transform 1 0 11040 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__809__A0
timestamp 1666464484
transform -1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__811__A0
timestamp 1666464484
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__813__A0
timestamp 1666464484
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__815__A0
timestamp 1666464484
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__821__B
timestamp 1666464484
transform 1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__822__B
timestamp 1666464484
transform 1 0 5520 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__823__B
timestamp 1666464484
transform -1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__824__B
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__856__SET_B
timestamp 1666464484
transform -1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__953__CLK
timestamp 1666464484
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__955__CLK
timestamp 1666464484
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__956__CLK
timestamp 1666464484
transform 1 0 9200 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__961__D
timestamp 1666464484
transform 1 0 21988 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__962__D
timestamp 1666464484
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1666464484
transform -1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout18_A
timestamp 1666464484
transform -1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout19_A
timestamp 1666464484
transform 1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout20_A
timestamp 1666464484
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout23_A
timestamp 1666464484
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout24_A
timestamp 1666464484
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout25_A
timestamp 1666464484
transform -1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold1_A
timestamp 1666464484
transform -1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 1748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 1748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 3496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 1748 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 6716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1666464484
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19
timestamp 1666464484
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1666464484
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1666464484
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1666464484
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1666464484
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_287
timestamp 1666464484
transform 1 0 27508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1666464484
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1666464484
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_61
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_73
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_85
timestamp 1666464484
transform 1 0 8924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_97
timestamp 1666464484
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1666464484
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_287
timestamp 1666464484
transform 1 0 27508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1666464484
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1666464484
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1666464484
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1666464484
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1666464484
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1666464484
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1666464484
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_285
timestamp 1666464484
transform 1 0 27324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1666464484
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_35
timestamp 1666464484
transform 1 0 4324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_41
timestamp 1666464484
transform 1 0 4876 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_47
timestamp 1666464484
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1666464484
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 1666464484
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp 1666464484
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_72
timestamp 1666464484
transform 1 0 7728 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_78
timestamp 1666464484
transform 1 0 8280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_84
timestamp 1666464484
transform 1 0 8832 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1666464484
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_99
timestamp 1666464484
transform 1 0 10212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_202
timestamp 1666464484
transform 1 0 19688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1666464484
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_287
timestamp 1666464484
transform 1 0 27508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1666464484
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1666464484
transform 1 0 2576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1666464484
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_38
timestamp 1666464484
transform 1 0 4600 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_44
timestamp 1666464484
transform 1 0 5152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_89
timestamp 1666464484
transform 1 0 9292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_277
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_285
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1666464484
transform 1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_32
timestamp 1666464484
transform 1 0 4048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_40
timestamp 1666464484
transform 1 0 4784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1666464484
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1666464484
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1666464484
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1666464484
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_83
timestamp 1666464484
transform 1 0 8740 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_88
timestamp 1666464484
transform 1 0 9200 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1666464484
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1666464484
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_119
timestamp 1666464484
transform 1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_126
timestamp 1666464484
transform 1 0 12696 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1666464484
transform 1 0 13800 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_146
timestamp 1666464484
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_151
timestamp 1666464484
transform 1 0 14996 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1666464484
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1666464484
transform 1 0 17204 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_183
timestamp 1666464484
transform 1 0 17940 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1666464484
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_218
timestamp 1666464484
transform 1 0 21160 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1666464484
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_287
timestamp 1666464484
transform 1 0 27508 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_8
timestamp 1666464484
transform 1 0 1840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_16
timestamp 1666464484
transform 1 0 2576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1666464484
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_35
timestamp 1666464484
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_39
timestamp 1666464484
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_43
timestamp 1666464484
transform 1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1666464484
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1666464484
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1666464484
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_128
timestamp 1666464484
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1666464484
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_147
timestamp 1666464484
transform 1 0 14628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1666464484
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1666464484
transform 1 0 16560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1666464484
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1666464484
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_219
timestamp 1666464484
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_231
timestamp 1666464484
transform 1 0 22356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_243
timestamp 1666464484
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_285
timestamp 1666464484
transform 1 0 27324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1666464484
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1666464484
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_35
timestamp 1666464484
transform 1 0 4324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1666464484
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp 1666464484
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1666464484
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_102
timestamp 1666464484
transform 1 0 10488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1666464484
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1666464484
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1666464484
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_148
timestamp 1666464484
transform 1 0 14720 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1666464484
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1666464484
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1666464484
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1666464484
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_232
timestamp 1666464484
transform 1 0 22448 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1666464484
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1666464484
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_287
timestamp 1666464484
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1666464484
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1666464484
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 1666464484
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_42
timestamp 1666464484
transform 1 0 4968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_66
timestamp 1666464484
transform 1 0 7176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1666464484
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1666464484
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1666464484
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1666464484
transform 1 0 14444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1666464484
transform 1 0 16652 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_185
timestamp 1666464484
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1666464484
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_203
timestamp 1666464484
transform 1 0 19780 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_211
timestamp 1666464484
transform 1 0 20516 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_235
timestamp 1666464484
transform 1 0 22724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1666464484
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1666464484
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_277
timestamp 1666464484
transform 1 0 26588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_285
timestamp 1666464484
transform 1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1666464484
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1666464484
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_36
timestamp 1666464484
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1666464484
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1666464484
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_72
timestamp 1666464484
transform 1 0 7728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1666464484
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_101
timestamp 1666464484
transform 1 0 10396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1666464484
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1666464484
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1666464484
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_142
timestamp 1666464484
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1666464484
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_175
timestamp 1666464484
transform 1 0 17204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1666464484
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_197
timestamp 1666464484
transform 1 0 19228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1666464484
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1666464484
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_254
timestamp 1666464484
transform 1 0 24472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1666464484
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1666464484
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1666464484
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_287
timestamp 1666464484
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1666464484
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1666464484
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1666464484
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1666464484
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_60
timestamp 1666464484
transform 1 0 6624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1666464484
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_89
timestamp 1666464484
transform 1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1666464484
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_150
timestamp 1666464484
transform 1 0 14904 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1666464484
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_168
timestamp 1666464484
transform 1 0 16560 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1666464484
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_201
timestamp 1666464484
transform 1 0 19596 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_205
timestamp 1666464484
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1666464484
transform 1 0 20424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_234
timestamp 1666464484
transform 1 0 22632 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_268
timestamp 1666464484
transform 1 0 25760 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_274
timestamp 1666464484
transform 1 0 26312 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_286
timestamp 1666464484
transform 1 0 27416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1666464484
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_23
timestamp 1666464484
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_31
timestamp 1666464484
transform 1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_44
timestamp 1666464484
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1666464484
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_72
timestamp 1666464484
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1666464484
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1666464484
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1666464484
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_119
timestamp 1666464484
transform 1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_157
timestamp 1666464484
transform 1 0 15548 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1666464484
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_173
timestamp 1666464484
transform 1 0 17020 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_185
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1666464484
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1666464484
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_234
timestamp 1666464484
transform 1 0 22632 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_240
timestamp 1666464484
transform 1 0 23184 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_261
timestamp 1666464484
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1666464484
transform 1 0 25852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1666464484
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_287
timestamp 1666464484
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1666464484
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1666464484
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_36
timestamp 1666464484
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1666464484
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_68
timestamp 1666464484
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_74
timestamp 1666464484
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1666464484
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1666464484
transform 1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1666464484
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1666464484
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1666464484
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1666464484
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1666464484
transform 1 0 14812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_169
timestamp 1666464484
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_180
timestamp 1666464484
transform 1 0 17664 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1666464484
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1666464484
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_232
timestamp 1666464484
transform 1 0 22448 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_243
timestamp 1666464484
transform 1 0 23460 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1666464484
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_268
timestamp 1666464484
transform 1 0 25760 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_274
timestamp 1666464484
transform 1 0 26312 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_286
timestamp 1666464484
transform 1 0 27416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 1666464484
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_26
timestamp 1666464484
transform 1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_30
timestamp 1666464484
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_35
timestamp 1666464484
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1666464484
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1666464484
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_80
timestamp 1666464484
transform 1 0 8464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1666464484
transform 1 0 11960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1666464484
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_138
timestamp 1666464484
transform 1 0 13800 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1666464484
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_180
timestamp 1666464484
transform 1 0 17664 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1666464484
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_212
timestamp 1666464484
transform 1 0 20608 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1666464484
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1666464484
transform 1 0 22632 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_242
timestamp 1666464484
transform 1 0 23368 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_266
timestamp 1666464484
transform 1 0 25576 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1666464484
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_287
timestamp 1666464484
transform 1 0 27508 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1666464484
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1666464484
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_39
timestamp 1666464484
transform 1 0 4692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_43
timestamp 1666464484
transform 1 0 5060 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1666464484
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1666464484
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1666464484
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1666464484
transform 1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_108
timestamp 1666464484
transform 1 0 11040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_114
timestamp 1666464484
transform 1 0 11592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1666464484
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_132
timestamp 1666464484
transform 1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1666464484
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1666464484
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1666464484
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_173
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1666464484
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_208
timestamp 1666464484
transform 1 0 20240 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_212
timestamp 1666464484
transform 1 0 20608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_229
timestamp 1666464484
transform 1 0 22172 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_242
timestamp 1666464484
transform 1 0 23368 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1666464484
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_259
timestamp 1666464484
transform 1 0 24932 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1666464484
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_285
timestamp 1666464484
transform 1 0 27324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1666464484
transform 1 0 2208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_32
timestamp 1666464484
transform 1 0 4048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_38
timestamp 1666464484
transform 1 0 4600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1666464484
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_66
timestamp 1666464484
transform 1 0 7176 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_72
timestamp 1666464484
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1666464484
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1666464484
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_132
timestamp 1666464484
transform 1 0 13248 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1666464484
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1666464484
transform 1 0 14720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1666464484
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_192
timestamp 1666464484
transform 1 0 18768 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_201
timestamp 1666464484
transform 1 0 19596 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_207
timestamp 1666464484
transform 1 0 20148 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_211
timestamp 1666464484
transform 1 0 20516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1666464484
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1666464484
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1666464484
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_266
timestamp 1666464484
transform 1 0 25576 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1666464484
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1666464484
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1666464484
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1666464484
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_40
timestamp 1666464484
transform 1 0 4784 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_52
timestamp 1666464484
transform 1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 1666464484
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1666464484
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1666464484
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1666464484
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_91
timestamp 1666464484
transform 1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1666464484
transform 1 0 11868 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1666464484
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1666464484
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1666464484
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_176
timestamp 1666464484
transform 1 0 17296 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1666464484
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1666464484
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_201
timestamp 1666464484
transform 1 0 19596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1666464484
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1666464484
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_239
timestamp 1666464484
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_275
timestamp 1666464484
transform 1 0 26404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_287
timestamp 1666464484
transform 1 0 27508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1666464484
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_33
timestamp 1666464484
transform 1 0 4140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_46
timestamp 1666464484
transform 1 0 5336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_50
timestamp 1666464484
transform 1 0 5704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1666464484
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_66
timestamp 1666464484
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_70
timestamp 1666464484
transform 1 0 7544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1666464484
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_85
timestamp 1666464484
transform 1 0 8924 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1666464484
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_106
timestamp 1666464484
transform 1 0 10856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1666464484
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1666464484
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1666464484
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1666464484
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_156
timestamp 1666464484
transform 1 0 15456 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1666464484
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1666464484
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_178
timestamp 1666464484
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1666464484
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1666464484
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1666464484
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1666464484
transform 1 0 20976 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1666464484
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_243
timestamp 1666464484
transform 1 0 23460 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_255
timestamp 1666464484
transform 1 0 24564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1666464484
transform 1 0 25668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_287
timestamp 1666464484
transform 1 0 27508 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1666464484
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_17
timestamp 1666464484
transform 1 0 2668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1666464484
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1666464484
transform 1 0 4784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_60
timestamp 1666464484
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1666464484
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1666464484
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_108
timestamp 1666464484
transform 1 0 11040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1666464484
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1666464484
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_156
timestamp 1666464484
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_176
timestamp 1666464484
transform 1 0 17296 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1666464484
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_204
timestamp 1666464484
transform 1 0 19872 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_216
timestamp 1666464484
transform 1 0 20976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_227
timestamp 1666464484
transform 1 0 21988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_235
timestamp 1666464484
transform 1 0 22724 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_243
timestamp 1666464484
transform 1 0 23460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1666464484
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1666464484
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_285
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_8
timestamp 1666464484
transform 1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_32
timestamp 1666464484
transform 1 0 4048 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1666464484
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1666464484
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_72
timestamp 1666464484
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_97
timestamp 1666464484
transform 1 0 10028 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1666464484
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_126
timestamp 1666464484
transform 1 0 12696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1666464484
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1666464484
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_180
timestamp 1666464484
transform 1 0 17664 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_194
timestamp 1666464484
transform 1 0 18952 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1666464484
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1666464484
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1666464484
transform 1 0 20884 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1666464484
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1666464484
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_242
timestamp 1666464484
transform 1 0 23368 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_248
timestamp 1666464484
transform 1 0 23920 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_260
timestamp 1666464484
transform 1 0 25024 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_267
timestamp 1666464484
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_287
timestamp 1666464484
transform 1 0 27508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_10
timestamp 1666464484
transform 1 0 2024 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1666464484
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_22
timestamp 1666464484
transform 1 0 3128 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1666464484
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1666464484
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_42
timestamp 1666464484
transform 1 0 4968 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_49
timestamp 1666464484
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1666464484
transform 1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1666464484
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1666464484
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1666464484
transform 1 0 12052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1666464484
transform 1 0 13248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1666464484
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1666464484
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1666464484
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1666464484
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1666464484
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1666464484
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_219
timestamp 1666464484
transform 1 0 21252 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_259
timestamp 1666464484
transform 1 0 24932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_283
timestamp 1666464484
transform 1 0 27140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_287
timestamp 1666464484
transform 1 0 27508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1666464484
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_23
timestamp 1666464484
transform 1 0 3220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_30
timestamp 1666464484
transform 1 0 3864 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_37
timestamp 1666464484
transform 1 0 4508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_43
timestamp 1666464484
transform 1 0 5060 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_47
timestamp 1666464484
transform 1 0 5428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1666464484
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_63
timestamp 1666464484
transform 1 0 6900 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_90
timestamp 1666464484
transform 1 0 9384 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_101
timestamp 1666464484
transform 1 0 10396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1666464484
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1666464484
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1666464484
transform 1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1666464484
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_214
timestamp 1666464484
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_218
timestamp 1666464484
transform 1 0 21160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1666464484
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_243
timestamp 1666464484
transform 1 0 23460 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1666464484
transform 1 0 24380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1666464484
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_285
timestamp 1666464484
transform 1 0 27324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1666464484
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_37
timestamp 1666464484
transform 1 0 4508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_44
timestamp 1666464484
transform 1 0 5152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1666464484
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1666464484
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_66
timestamp 1666464484
transform 1 0 7176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1666464484
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1666464484
transform 1 0 8280 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1666464484
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_91
timestamp 1666464484
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1666464484
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_132
timestamp 1666464484
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1666464484
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1666464484
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_180
timestamp 1666464484
transform 1 0 17664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_184
timestamp 1666464484
transform 1 0 18032 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1666464484
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_202
timestamp 1666464484
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_233
timestamp 1666464484
transform 1 0 22540 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1666464484
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_257
timestamp 1666464484
transform 1 0 24748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_261
timestamp 1666464484
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_275
timestamp 1666464484
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_283
timestamp 1666464484
transform 1 0 27140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_287
timestamp 1666464484
transform 1 0 27508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_7
timestamp 1666464484
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1666464484
transform 1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1666464484
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1666464484
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1666464484
transform 1 0 6808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1666464484
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_76
timestamp 1666464484
transform 1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1666464484
transform 1 0 8740 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1666464484
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1666464484
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1666464484
transform 1 0 12512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_128
timestamp 1666464484
transform 1 0 12880 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_174
timestamp 1666464484
transform 1 0 17112 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1666464484
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_203
timestamp 1666464484
transform 1 0 19780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1666464484
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_247
timestamp 1666464484
transform 1 0 23828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_258
timestamp 1666464484
transform 1 0 24840 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1666464484
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_285
timestamp 1666464484
transform 1 0 27324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1666464484
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_37
timestamp 1666464484
transform 1 0 4508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1666464484
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1666464484
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_76
timestamp 1666464484
transform 1 0 8096 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1666464484
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1666464484
transform 1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1666464484
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1666464484
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_151
timestamp 1666464484
transform 1 0 14996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_157
timestamp 1666464484
transform 1 0 15548 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_178
timestamp 1666464484
transform 1 0 17480 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_186
timestamp 1666464484
transform 1 0 18216 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_202
timestamp 1666464484
transform 1 0 19688 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1666464484
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_233
timestamp 1666464484
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1666464484
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_261
timestamp 1666464484
transform 1 0 25116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_286
timestamp 1666464484
transform 1 0 27416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1666464484
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_28
timestamp 1666464484
transform 1 0 3680 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1666464484
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_63
timestamp 1666464484
transform 1 0 6900 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_67
timestamp 1666464484
transform 1 0 7268 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1666464484
transform 1 0 7636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_78
timestamp 1666464484
transform 1 0 8280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1666464484
transform 1 0 10120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1666464484
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1666464484
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1666464484
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1666464484
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_182
timestamp 1666464484
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1666464484
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_210
timestamp 1666464484
transform 1 0 20424 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1666464484
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1666464484
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_271
timestamp 1666464484
transform 1 0 26036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1666464484
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_285
timestamp 1666464484
transform 1 0 27324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1666464484
transform 1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1666464484
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_35
timestamp 1666464484
transform 1 0 4324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_43
timestamp 1666464484
transform 1 0 5060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1666464484
transform 1 0 5796 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_63
timestamp 1666464484
transform 1 0 6900 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1666464484
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1666464484
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_103
timestamp 1666464484
transform 1 0 10580 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1666464484
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1666464484
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1666464484
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1666464484
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1666464484
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1666464484
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_211
timestamp 1666464484
transform 1 0 20516 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_217
timestamp 1666464484
transform 1 0 21068 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1666464484
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1666464484
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_268
timestamp 1666464484
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_285
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_9
timestamp 1666464484
transform 1 0 1932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1666464484
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_24
timestamp 1666464484
transform 1 0 3312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1666464484
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_40
timestamp 1666464484
transform 1 0 4784 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_48
timestamp 1666464484
transform 1 0 5520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1666464484
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_75
timestamp 1666464484
transform 1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1666464484
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_86
timestamp 1666464484
transform 1 0 9016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1666464484
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1666464484
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1666464484
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1666464484
transform 1 0 14352 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1666464484
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1666464484
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1666464484
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1666464484
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1666464484
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_242
timestamp 1666464484
transform 1 0 23368 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp 1666464484
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1666464484
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_287
timestamp 1666464484
transform 1 0 27508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1666464484
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_52
timestamp 1666464484
transform 1 0 5888 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1666464484
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_64
timestamp 1666464484
transform 1 0 6992 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_71
timestamp 1666464484
transform 1 0 7636 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_79
timestamp 1666464484
transform 1 0 8372 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1666464484
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_96
timestamp 1666464484
transform 1 0 9936 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 1666464484
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_118
timestamp 1666464484
transform 1 0 11960 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_124
timestamp 1666464484
transform 1 0 12512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1666464484
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_150
timestamp 1666464484
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1666464484
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1666464484
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_187
timestamp 1666464484
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1666464484
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_213
timestamp 1666464484
transform 1 0 20700 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_217
timestamp 1666464484
transform 1 0 21068 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_225
timestamp 1666464484
transform 1 0 21804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_240
timestamp 1666464484
transform 1 0 23184 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_244
timestamp 1666464484
transform 1 0 23552 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_259
timestamp 1666464484
transform 1 0 24932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_286
timestamp 1666464484
transform 1 0 27416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1666464484
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_29
timestamp 1666464484
transform 1 0 3772 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1666464484
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_62
timestamp 1666464484
transform 1 0 6808 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1666464484
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1666464484
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1666464484
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_127
timestamp 1666464484
transform 1 0 12788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_151
timestamp 1666464484
transform 1 0 14996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1666464484
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1666464484
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_175
timestamp 1666464484
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_183
timestamp 1666464484
transform 1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_187
timestamp 1666464484
transform 1 0 18308 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1666464484
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_216
timestamp 1666464484
transform 1 0 20976 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1666464484
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1666464484
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_246
timestamp 1666464484
transform 1 0 23736 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_252
timestamp 1666464484
transform 1 0 24288 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_258
timestamp 1666464484
transform 1 0 24840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1666464484
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 1666464484
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_8
timestamp 1666464484
transform 1 0 1840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_14
timestamp 1666464484
transform 1 0 2392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_20
timestamp 1666464484
transform 1 0 2944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1666464484
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1666464484
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_37
timestamp 1666464484
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1666464484
transform 1 0 6808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1666464484
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1666464484
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1666464484
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1666464484
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_131
timestamp 1666464484
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1666464484
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_148
timestamp 1666464484
transform 1 0 14720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_156
timestamp 1666464484
transform 1 0 15456 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_173
timestamp 1666464484
transform 1 0 17020 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_181
timestamp 1666464484
transform 1 0 17756 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_186
timestamp 1666464484
transform 1 0 18216 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_190
timestamp 1666464484
transform 1 0 18584 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_215
timestamp 1666464484
transform 1 0 20884 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1666464484
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1666464484
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1666464484
transform 1 0 26496 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1666464484
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_21
timestamp 1666464484
transform 1 0 3036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_29
timestamp 1666464484
transform 1 0 3772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_34
timestamp 1666464484
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1666464484
transform 1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_44
timestamp 1666464484
transform 1 0 5152 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_48
timestamp 1666464484
transform 1 0 5520 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1666464484
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1666464484
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1666464484
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1666464484
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1666464484
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_180
timestamp 1666464484
transform 1 0 17664 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1666464484
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_204
timestamp 1666464484
transform 1 0 19872 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1666464484
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1666464484
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_236
timestamp 1666464484
transform 1 0 22816 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_246
timestamp 1666464484
transform 1 0 23736 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1666464484
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_287
timestamp 1666464484
transform 1 0 27508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1666464484
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1666464484
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_38
timestamp 1666464484
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_44
timestamp 1666464484
transform 1 0 5152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_50
timestamp 1666464484
transform 1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1666464484
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_67
timestamp 1666464484
transform 1 0 7268 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_71
timestamp 1666464484
transform 1 0 7636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_79
timestamp 1666464484
transform 1 0 8372 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1666464484
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_90
timestamp 1666464484
transform 1 0 9384 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_96
timestamp 1666464484
transform 1 0 9936 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_104
timestamp 1666464484
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1666464484
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1666464484
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_131
timestamp 1666464484
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1666464484
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1666464484
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1666464484
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1666464484
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1666464484
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1666464484
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_218
timestamp 1666464484
transform 1 0 21160 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_238
timestamp 1666464484
transform 1 0 23000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_262
timestamp 1666464484
transform 1 0 25208 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_278
timestamp 1666464484
transform 1 0 26680 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_286
timestamp 1666464484
transform 1 0 27416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_9
timestamp 1666464484
transform 1 0 1932 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_20
timestamp 1666464484
transform 1 0 2944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_62
timestamp 1666464484
transform 1 0 6808 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_68
timestamp 1666464484
transform 1 0 7360 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_71
timestamp 1666464484
transform 1 0 7636 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1666464484
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_85
timestamp 1666464484
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1666464484
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_101
timestamp 1666464484
transform 1 0 10396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_107
timestamp 1666464484
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1666464484
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_121
timestamp 1666464484
transform 1 0 12236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1666464484
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1666464484
transform 1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_152
timestamp 1666464484
transform 1 0 15088 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1666464484
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1666464484
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_189
timestamp 1666464484
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_195
timestamp 1666464484
transform 1 0 19044 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_212
timestamp 1666464484
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1666464484
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1666464484
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_239
timestamp 1666464484
transform 1 0 23092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_246
timestamp 1666464484
transform 1 0 23736 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_252
timestamp 1666464484
transform 1 0 24288 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_258
timestamp 1666464484
transform 1 0 24840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1666464484
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1666464484
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_287
timestamp 1666464484
transform 1 0 27508 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1666464484
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_35
timestamp 1666464484
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_39
timestamp 1666464484
transform 1 0 4692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1666464484
transform 1 0 6992 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_71
timestamp 1666464484
transform 1 0 7636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1666464484
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_94
timestamp 1666464484
transform 1 0 9752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_101
timestamp 1666464484
transform 1 0 10396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_114
timestamp 1666464484
transform 1 0 11592 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_124
timestamp 1666464484
transform 1 0 12512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1666464484
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1666464484
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_152
timestamp 1666464484
transform 1 0 15088 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_164
timestamp 1666464484
transform 1 0 16192 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1666464484
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_216
timestamp 1666464484
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_223
timestamp 1666464484
transform 1 0 21620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1666464484
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_285
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_7
timestamp 1666464484
transform 1 0 1748 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1666464484
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_42
timestamp 1666464484
transform 1 0 4968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_49
timestamp 1666464484
transform 1 0 5612 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_79
timestamp 1666464484
transform 1 0 8372 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1666464484
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_90
timestamp 1666464484
transform 1 0 9384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1666464484
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1666464484
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_131
timestamp 1666464484
transform 1 0 13156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_151
timestamp 1666464484
transform 1 0 14996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_189
timestamp 1666464484
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1666464484
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_216
timestamp 1666464484
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_243
timestamp 1666464484
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_255
timestamp 1666464484
transform 1 0 24564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_267
timestamp 1666464484
transform 1 0 25668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1666464484
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_7
timestamp 1666464484
transform 1 0 1748 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_17
timestamp 1666464484
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_21
timestamp 1666464484
transform 1 0 3036 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1666464484
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_52
timestamp 1666464484
transform 1 0 5888 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1666464484
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1666464484
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1666464484
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1666464484
transform 1 0 9660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1666464484
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_126
timestamp 1666464484
transform 1 0 12696 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_134
timestamp 1666464484
transform 1 0 13432 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1666464484
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1666464484
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_163
timestamp 1666464484
transform 1 0 16100 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_167
timestamp 1666464484
transform 1 0 16468 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_187
timestamp 1666464484
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1666464484
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1666464484
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_213
timestamp 1666464484
transform 1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_220
timestamp 1666464484
transform 1 0 21344 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1666464484
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1666464484
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_285
timestamp 1666464484
transform 1 0 27324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_14
timestamp 1666464484
transform 1 0 2392 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_22
timestamp 1666464484
transform 1 0 3128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_26
timestamp 1666464484
transform 1 0 3496 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_36
timestamp 1666464484
transform 1 0 4416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_46
timestamp 1666464484
transform 1 0 5336 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1666464484
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_79
timestamp 1666464484
transform 1 0 8372 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_87
timestamp 1666464484
transform 1 0 9108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1666464484
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1666464484
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1666464484
transform 1 0 11960 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1666464484
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_145
timestamp 1666464484
transform 1 0 14444 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1666464484
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1666464484
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_182
timestamp 1666464484
transform 1 0 17848 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_190
timestamp 1666464484
transform 1 0 18584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1666464484
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_215
timestamp 1666464484
transform 1 0 20884 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_219
timestamp 1666464484
transform 1 0 21252 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_229
timestamp 1666464484
transform 1 0 22172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_241
timestamp 1666464484
transform 1 0 23276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_253
timestamp 1666464484
transform 1 0 24380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_265
timestamp 1666464484
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1666464484
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1666464484
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1666464484
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 1666464484
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_50
timestamp 1666464484
transform 1 0 5704 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_56
timestamp 1666464484
transform 1 0 6256 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_73
timestamp 1666464484
transform 1 0 7820 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_81
timestamp 1666464484
transform 1 0 8556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1666464484
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1666464484
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_113
timestamp 1666464484
transform 1 0 11500 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_132
timestamp 1666464484
transform 1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1666464484
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_152
timestamp 1666464484
transform 1 0 15088 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_164
timestamp 1666464484
transform 1 0 16192 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1666464484
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1666464484
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_201
timestamp 1666464484
transform 1 0 19596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_222
timestamp 1666464484
transform 1 0 21528 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_230
timestamp 1666464484
transform 1 0 22264 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_242
timestamp 1666464484
transform 1 0 23368 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_277
timestamp 1666464484
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_285
timestamp 1666464484
transform 1 0 27324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_22
timestamp 1666464484
transform 1 0 3128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_30
timestamp 1666464484
transform 1 0 3864 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1666464484
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1666464484
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1666464484
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_74
timestamp 1666464484
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1666464484
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_101
timestamp 1666464484
transform 1 0 10396 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_104
timestamp 1666464484
transform 1 0 10672 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1666464484
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_124
timestamp 1666464484
transform 1 0 12512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_128
timestamp 1666464484
transform 1 0 12880 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1666464484
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1666464484
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1666464484
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_287
timestamp 1666464484
transform 1 0 27508 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1666464484
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_38
timestamp 1666464484
transform 1 0 4600 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1666464484
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_71
timestamp 1666464484
transform 1 0 7636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1666464484
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_103
timestamp 1666464484
transform 1 0 10580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1666464484
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1666464484
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_147
timestamp 1666464484
transform 1 0 14628 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_170
timestamp 1666464484
transform 1 0 16744 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1666464484
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_212
timestamp 1666464484
transform 1 0 20608 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_220
timestamp 1666464484
transform 1 0 21344 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_232
timestamp 1666464484
transform 1 0 22448 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_244
timestamp 1666464484
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_285
timestamp 1666464484
transform 1 0 27324 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_11
timestamp 1666464484
transform 1 0 2116 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_28
timestamp 1666464484
transform 1 0 3680 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_43
timestamp 1666464484
transform 1 0 5060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1666464484
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_63
timestamp 1666464484
transform 1 0 6900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1666464484
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_91
timestamp 1666464484
transform 1 0 9476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_101
timestamp 1666464484
transform 1 0 10396 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1666464484
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_117
timestamp 1666464484
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_122
timestamp 1666464484
transform 1 0 12328 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1666464484
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_142
timestamp 1666464484
transform 1 0 14168 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1666464484
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_175
timestamp 1666464484
transform 1 0 17204 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_183
timestamp 1666464484
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_208
timestamp 1666464484
transform 1 0 20240 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1666464484
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1666464484
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_9
timestamp 1666464484
transform 1 0 1932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1666464484
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_36
timestamp 1666464484
transform 1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_46
timestamp 1666464484
transform 1 0 5336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_58
timestamp 1666464484
transform 1 0 6440 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_70
timestamp 1666464484
transform 1 0 7544 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1666464484
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_94
timestamp 1666464484
transform 1 0 9752 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_102
timestamp 1666464484
transform 1 0 10488 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1666464484
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_145
timestamp 1666464484
transform 1 0 14444 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_149
timestamp 1666464484
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_154
timestamp 1666464484
transform 1 0 15272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_178
timestamp 1666464484
transform 1 0 17480 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_186
timestamp 1666464484
transform 1 0 18216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1666464484
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_219
timestamp 1666464484
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_231
timestamp 1666464484
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1666464484
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_285
timestamp 1666464484
transform 1 0 27324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1666464484
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_11
timestamp 1666464484
transform 1 0 2116 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_19
timestamp 1666464484
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_31
timestamp 1666464484
transform 1 0 3956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_35
timestamp 1666464484
transform 1 0 4324 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1666464484
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_63
timestamp 1666464484
transform 1 0 6900 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_75
timestamp 1666464484
transform 1 0 8004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_83
timestamp 1666464484
transform 1 0 8740 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_91
timestamp 1666464484
transform 1 0 9476 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1666464484
transform 1 0 10212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1666464484
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_120
timestamp 1666464484
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_128
timestamp 1666464484
transform 1 0 12880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_152
timestamp 1666464484
transform 1 0 15088 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_160
timestamp 1666464484
transform 1 0 15824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1666464484
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_176
timestamp 1666464484
transform 1 0 17296 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_188
timestamp 1666464484
transform 1 0 18400 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_199
timestamp 1666464484
transform 1 0 19412 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1666464484
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1666464484
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_287
timestamp 1666464484
transform 1 0 27508 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1666464484
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1666464484
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_46
timestamp 1666464484
transform 1 0 5336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_54
timestamp 1666464484
transform 1 0 6072 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_57
timestamp 1666464484
transform 1 0 6348 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_62
timestamp 1666464484
transform 1 0 6808 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_74
timestamp 1666464484
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1666464484
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_91
timestamp 1666464484
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_98
timestamp 1666464484
transform 1 0 10120 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_110
timestamp 1666464484
transform 1 0 11224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_113
timestamp 1666464484
transform 1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_117
timestamp 1666464484
transform 1 0 11868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1666464484
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_147
timestamp 1666464484
transform 1 0 14628 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1666464484
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_169
timestamp 1666464484
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_175
timestamp 1666464484
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1666464484
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_203
timestamp 1666464484
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_211
timestamp 1666464484
transform 1 0 20516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_223
timestamp 1666464484
transform 1 0 21620 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_225
timestamp 1666464484
transform 1 0 21804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_237
timestamp 1666464484
transform 1 0 22908 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_247
timestamp 1666464484
transform 1 0 23828 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_273
timestamp 1666464484
transform 1 0 26220 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_278
timestamp 1666464484
transform 1 0 26680 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_281
timestamp 1666464484
transform 1 0 26956 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_287
timestamp 1666464484
transform 1 0 27508 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 27876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 27876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 27876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 27876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 27876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 27876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 27876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 27876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 27876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 27876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 27876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 27876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 27876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 27876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 27876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 27876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 27876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 27876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 27876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 27876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 27876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 27876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 27876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 27876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 27876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 27876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 27876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 27876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 27876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 27876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 27876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 27876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 27876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 27876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 27876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 6256 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 11408 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 16560 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 21712 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 26864 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _380_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _381_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1666464484
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1666464484
transform -1 0 3864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1666464484
transform -1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1666464484
transform -1 0 1840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1666464484
transform -1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _389_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _390_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10580 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12144 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _392_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6072 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _393_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _394_
timestamp 1666464484
transform 1 0 7636 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1666464484
transform 1 0 6624 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _396_
timestamp 1666464484
transform 1 0 6532 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _397_
timestamp 1666464484
transform 1 0 11684 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1666464484
transform 1 0 10028 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1666464484
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1666464484
transform 1 0 7820 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1666464484
transform -1 0 7452 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _403_
timestamp 1666464484
transform 1 0 3956 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _404_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7544 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _405_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_4  _406_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__o211ai_4  _407_
timestamp 1666464484
transform -1 0 15824 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1666464484
transform -1 0 13800 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1666464484
transform -1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _410_
timestamp 1666464484
transform 1 0 3036 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _411_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11960 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _412_
timestamp 1666464484
transform 1 0 11868 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _413_
timestamp 1666464484
transform 1 0 14444 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _414_
timestamp 1666464484
transform -1 0 20700 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _415_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15364 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _416_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16560 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _418_
timestamp 1666464484
transform -1 0 17388 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _419_
timestamp 1666464484
transform 1 0 18400 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _420_
timestamp 1666464484
transform 1 0 13248 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _421_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _422_
timestamp 1666464484
transform -1 0 17848 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _423_
timestamp 1666464484
transform -1 0 19320 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _424_
timestamp 1666464484
transform 1 0 12328 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _425_
timestamp 1666464484
transform 1 0 15732 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _426_
timestamp 1666464484
transform 1 0 16560 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_2  _428_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11960 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _430_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15548 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _431_
timestamp 1666464484
transform 1 0 14996 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _432_
timestamp 1666464484
transform 1 0 12972 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _433_
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _434_
timestamp 1666464484
transform 1 0 12052 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_8  _435_
timestamp 1666464484
transform -1 0 20516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_2  _436_
timestamp 1666464484
transform -1 0 18492 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _437_
timestamp 1666464484
transform 1 0 19688 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _438_
timestamp 1666464484
transform 1 0 19504 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _439_
timestamp 1666464484
transform -1 0 20608 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _440_
timestamp 1666464484
transform 1 0 17480 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_16  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 6716 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__xor2_1  _442_
timestamp 1666464484
transform -1 0 13708 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _443_
timestamp 1666464484
transform 1 0 11040 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _444_
timestamp 1666464484
transform 1 0 11684 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _445_
timestamp 1666464484
transform -1 0 14904 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _446_
timestamp 1666464484
transform -1 0 13248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _447_
timestamp 1666464484
transform 1 0 6900 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _448_
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1666464484
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _450_
timestamp 1666464484
transform -1 0 8648 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _451_
timestamp 1666464484
transform 1 0 6532 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _452_
timestamp 1666464484
transform 1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _453_
timestamp 1666464484
transform 1 0 6532 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _454_
timestamp 1666464484
transform 1 0 4968 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _455_
timestamp 1666464484
transform 1 0 5060 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _456_
timestamp 1666464484
transform -1 0 8648 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _457_
timestamp 1666464484
transform 1 0 7360 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _458_
timestamp 1666464484
transform 1 0 9108 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11224 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 12328 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10120 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _463_
timestamp 1666464484
transform -1 0 13248 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 7728 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _465_
timestamp 1666464484
transform -1 0 7728 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _466_
timestamp 1666464484
transform 1 0 9108 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_8  _467_
timestamp 1666464484
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_2  _468_
timestamp 1666464484
transform -1 0 10488 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _469_
timestamp 1666464484
transform 1 0 11500 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _470_
timestamp 1666464484
transform 1 0 10028 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _471_
timestamp 1666464484
transform 1 0 9476 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _472_
timestamp 1666464484
transform 1 0 7176 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _473_
timestamp 1666464484
transform 1 0 4876 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _474_
timestamp 1666464484
transform -1 0 7728 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _475__1
timestamp 1666464484
transform -1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _475__2
timestamp 1666464484
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _476_
timestamp 1666464484
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _477_
timestamp 1666464484
transform 1 0 19412 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _478_
timestamp 1666464484
transform 1 0 19412 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _479_
timestamp 1666464484
transform 1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _480_
timestamp 1666464484
transform -1 0 23460 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _481_
timestamp 1666464484
transform -1 0 18952 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _482_
timestamp 1666464484
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _483_
timestamp 1666464484
transform -1 0 18860 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _484_
timestamp 1666464484
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _485_
timestamp 1666464484
transform 1 0 16928 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17940 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _487_
timestamp 1666464484
transform -1 0 22632 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _488_
timestamp 1666464484
transform -1 0 22632 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _489_
timestamp 1666464484
transform -1 0 23644 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _490_
timestamp 1666464484
transform -1 0 23460 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _491_
timestamp 1666464484
transform 1 0 14536 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _492_
timestamp 1666464484
transform 1 0 17020 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _493_
timestamp 1666464484
transform 1 0 18216 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _494_
timestamp 1666464484
transform -1 0 18952 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _495_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _496_
timestamp 1666464484
transform 1 0 14260 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _497_
timestamp 1666464484
transform -1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _498_
timestamp 1666464484
transform 1 0 13524 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11500 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_2  _500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 16008 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _501_
timestamp 1666464484
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _502_
timestamp 1666464484
transform 1 0 21252 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _503_
timestamp 1666464484
transform 1 0 19320 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _504_
timestamp 1666464484
transform 1 0 18492 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _505_
timestamp 1666464484
transform 1 0 16652 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _506_
timestamp 1666464484
transform 1 0 14996 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _507_
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _508_
timestamp 1666464484
transform 1 0 23828 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _509_
timestamp 1666464484
transform -1 0 25760 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _510_
timestamp 1666464484
transform -1 0 25760 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _511_
timestamp 1666464484
transform -1 0 24012 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _512_
timestamp 1666464484
transform 1 0 23092 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _513_
timestamp 1666464484
transform 1 0 24564 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _514_
timestamp 1666464484
transform 1 0 24196 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _515_
timestamp 1666464484
transform 1 0 23184 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _516_
timestamp 1666464484
transform -1 0 25116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _517_
timestamp 1666464484
transform 1 0 19596 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _518_
timestamp 1666464484
transform 1 0 20424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _519_
timestamp 1666464484
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _520_
timestamp 1666464484
transform 1 0 19320 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _521_
timestamp 1666464484
transform 1 0 17480 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _522_
timestamp 1666464484
transform 1 0 20056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _523_
timestamp 1666464484
transform 1 0 18308 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _524_
timestamp 1666464484
transform 1 0 21896 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _525_
timestamp 1666464484
transform 1 0 20608 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _526_
timestamp 1666464484
transform 1 0 21896 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _527_
timestamp 1666464484
transform 1 0 23368 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _528_
timestamp 1666464484
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _529_
timestamp 1666464484
transform -1 0 14904 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _530_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 14260 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _531_
timestamp 1666464484
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _532_
timestamp 1666464484
transform -1 0 18768 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _533_
timestamp 1666464484
transform 1 0 18492 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _534_
timestamp 1666464484
transform 1 0 21988 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _535_
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _536_
timestamp 1666464484
transform 1 0 22172 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _537_
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _538_
timestamp 1666464484
transform 1 0 25208 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _539_
timestamp 1666464484
transform 1 0 25392 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _540_
timestamp 1666464484
transform 1 0 26128 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _541_
timestamp 1666464484
transform 1 0 25484 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _542_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26312 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _543_
timestamp 1666464484
transform -1 0 26496 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _544_
timestamp 1666464484
transform -1 0 27140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _545_
timestamp 1666464484
transform 1 0 24564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _546_
timestamp 1666464484
transform -1 0 24932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _547_
timestamp 1666464484
transform 1 0 26404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _548_
timestamp 1666464484
transform -1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _549_
timestamp 1666464484
transform 1 0 26312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _550_
timestamp 1666464484
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _551_
timestamp 1666464484
transform -1 0 20976 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _552_
timestamp 1666464484
transform -1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _553_
timestamp 1666464484
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _554_
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _555_
timestamp 1666464484
transform -1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _556_
timestamp 1666464484
transform -1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _557_
timestamp 1666464484
transform -1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _558_
timestamp 1666464484
transform 1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _559_
timestamp 1666464484
transform -1 0 23368 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _560_
timestamp 1666464484
transform 1 0 23736 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _561_
timestamp 1666464484
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _562_
timestamp 1666464484
transform -1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _563_
timestamp 1666464484
transform -1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _564_
timestamp 1666464484
transform -1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _565_
timestamp 1666464484
transform -1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _566_
timestamp 1666464484
transform -1 0 19780 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _567_
timestamp 1666464484
transform -1 0 20516 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _568_
timestamp 1666464484
transform -1 0 20424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _569_
timestamp 1666464484
transform -1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _570_
timestamp 1666464484
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _571_
timestamp 1666464484
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _572_
timestamp 1666464484
transform -1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1666464484
transform 1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _574_
timestamp 1666464484
transform 1 0 8280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _575_
timestamp 1666464484
transform 1 0 13984 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _576_
timestamp 1666464484
transform 1 0 11684 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _577_
timestamp 1666464484
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _578_
timestamp 1666464484
transform -1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _579_
timestamp 1666464484
transform -1 0 5888 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _580_
timestamp 1666464484
transform -1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _581_
timestamp 1666464484
transform 1 0 11040 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _582_
timestamp 1666464484
transform -1 0 18216 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _583_
timestamp 1666464484
transform -1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _584_
timestamp 1666464484
transform -1 0 20976 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _585_
timestamp 1666464484
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _586_
timestamp 1666464484
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _587_
timestamp 1666464484
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _588_
timestamp 1666464484
transform -1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _589_
timestamp 1666464484
transform -1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _590_
timestamp 1666464484
transform -1 0 14628 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _591_
timestamp 1666464484
transform -1 0 15272 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _592_
timestamp 1666464484
transform -1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _593_
timestamp 1666464484
transform -1 0 6808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _594_
timestamp 1666464484
transform 1 0 7728 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _595_
timestamp 1666464484
transform 1 0 6532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _596_
timestamp 1666464484
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _597_
timestamp 1666464484
transform -1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _598_
timestamp 1666464484
transform -1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _599_
timestamp 1666464484
transform 1 0 6532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _600_
timestamp 1666464484
transform 1 0 7544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _601_
timestamp 1666464484
transform -1 0 6072 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _602_
timestamp 1666464484
transform 1 0 4416 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7176 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _604_
timestamp 1666464484
transform -1 0 6808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5704 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _606_
timestamp 1666464484
transform 1 0 8832 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 8464 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _608_
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _609_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6440 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _610_
timestamp 1666464484
transform 1 0 8096 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _611_
timestamp 1666464484
transform 1 0 8280 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _612_
timestamp 1666464484
transform 1 0 8004 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 10396 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _614_
timestamp 1666464484
transform 1 0 6992 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _616_
timestamp 1666464484
transform 1 0 9568 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _617_
timestamp 1666464484
transform 1 0 9844 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _618_
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _619_
timestamp 1666464484
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 9752 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _621_
timestamp 1666464484
transform 1 0 10580 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 11132 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _623_
timestamp 1666464484
transform 1 0 4784 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _624_
timestamp 1666464484
transform 1 0 4416 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _625_
timestamp 1666464484
transform -1 0 4600 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _626_
timestamp 1666464484
transform -1 0 2852 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _627_
timestamp 1666464484
transform -1 0 2392 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _628_
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _629_
timestamp 1666464484
transform -1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _630_
timestamp 1666464484
transform 1 0 20608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _631_
timestamp 1666464484
transform -1 0 21344 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _632_
timestamp 1666464484
transform 1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _633_
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _634_
timestamp 1666464484
transform -1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _635_
timestamp 1666464484
transform 1 0 21712 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _636_
timestamp 1666464484
transform -1 0 21988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _637_
timestamp 1666464484
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _638_
timestamp 1666464484
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _639_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _640_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2024 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _641_
timestamp 1666464484
transform -1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 5428 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _643_
timestamp 1666464484
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _644_
timestamp 1666464484
transform -1 0 4600 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _645_
timestamp 1666464484
transform -1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _646_
timestamp 1666464484
transform 1 0 2944 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _647_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3864 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _648_
timestamp 1666464484
transform -1 0 2208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _649_
timestamp 1666464484
transform 1 0 2944 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _650_
timestamp 1666464484
transform 1 0 3956 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _651_
timestamp 1666464484
transform 1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _652_
timestamp 1666464484
transform -1 0 5336 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _653_
timestamp 1666464484
transform 1 0 3956 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _654_
timestamp 1666464484
transform 1 0 4784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _655_
timestamp 1666464484
transform 1 0 2668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _656_
timestamp 1666464484
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _657_
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _658_
timestamp 1666464484
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _659_
timestamp 1666464484
transform -1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _660_
timestamp 1666464484
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _661_
timestamp 1666464484
transform -1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _662_
timestamp 1666464484
transform 1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _663_
timestamp 1666464484
transform -1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _664_
timestamp 1666464484
transform 1 0 7360 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _665_
timestamp 1666464484
transform 1 0 2668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _666_
timestamp 1666464484
transform -1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _667_
timestamp 1666464484
transform -1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _668_
timestamp 1666464484
transform -1 0 17020 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _669_
timestamp 1666464484
transform 1 0 21988 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 1666464484
transform 1 0 21252 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _671_
timestamp 1666464484
transform -1 0 21344 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp 1666464484
transform 1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _673_
timestamp 1666464484
transform -1 0 17848 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _674_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _675_
timestamp 1666464484
transform -1 0 16376 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _676_
timestamp 1666464484
transform 1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_2  _677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 13248 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _678_
timestamp 1666464484
transform 1 0 18032 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _679_
timestamp 1666464484
transform -1 0 18952 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _680_
timestamp 1666464484
transform 1 0 20056 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _681_
timestamp 1666464484
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _682_
timestamp 1666464484
transform -1 0 21528 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _683_
timestamp 1666464484
transform -1 0 23736 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _684_
timestamp 1666464484
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _685_
timestamp 1666464484
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _686_
timestamp 1666464484
transform -1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _688_
timestamp 1666464484
transform 1 0 11684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _689_
timestamp 1666464484
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _690_
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _691_
timestamp 1666464484
transform -1 0 11224 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _692_
timestamp 1666464484
transform 1 0 9384 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1666464484
transform -1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _694_
timestamp 1666464484
transform 1 0 9384 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _695_
timestamp 1666464484
transform -1 0 8280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _696_
timestamp 1666464484
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _697_
timestamp 1666464484
transform -1 0 26588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _698_
timestamp 1666464484
transform -1 0 25668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _699_
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _700_
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _701_
timestamp 1666464484
transform 1 0 21160 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _702_
timestamp 1666464484
transform 1 0 14720 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _703_
timestamp 1666464484
transform 1 0 23368 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _704_
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _705_
timestamp 1666464484
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _706_
timestamp 1666464484
transform -1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _707_
timestamp 1666464484
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _708_
timestamp 1666464484
transform -1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _709_
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _710_
timestamp 1666464484
transform 1 0 24564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _711_
timestamp 1666464484
transform 1 0 14260 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _712_
timestamp 1666464484
transform -1 0 15548 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _713_
timestamp 1666464484
transform -1 0 13800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _714_
timestamp 1666464484
transform -1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _715_
timestamp 1666464484
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _716_
timestamp 1666464484
transform 1 0 18584 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _717_
timestamp 1666464484
transform -1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _718_
timestamp 1666464484
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _719_
timestamp 1666464484
transform 1 0 6532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _720_
timestamp 1666464484
transform -1 0 6072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _721_
timestamp 1666464484
transform 1 0 15272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _722_
timestamp 1666464484
transform -1 0 16376 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _723_
timestamp 1666464484
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _724_
timestamp 1666464484
transform 1 0 19780 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _725_
timestamp 1666464484
transform -1 0 19136 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _726_
timestamp 1666464484
transform -1 0 20608 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _727_
timestamp 1666464484
transform 1 0 21344 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _728_
timestamp 1666464484
transform -1 0 15916 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _729_
timestamp 1666464484
transform 1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _730_
timestamp 1666464484
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _731_
timestamp 1666464484
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _732_
timestamp 1666464484
transform -1 0 16376 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _733_
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _734_
timestamp 1666464484
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _735_
timestamp 1666464484
transform 1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _736_
timestamp 1666464484
transform -1 0 20240 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _737_
timestamp 1666464484
transform 1 0 17940 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _738_
timestamp 1666464484
transform -1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _739_
timestamp 1666464484
transform -1 0 19320 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _740_
timestamp 1666464484
transform 1 0 20976 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _741_
timestamp 1666464484
transform 1 0 19412 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _742_
timestamp 1666464484
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _743_
timestamp 1666464484
transform 1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _744_
timestamp 1666464484
transform 1 0 17848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _745_
timestamp 1666464484
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _746_
timestamp 1666464484
transform 1 0 5612 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _747_
timestamp 1666464484
transform 1 0 5704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _748_
timestamp 1666464484
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _749_
timestamp 1666464484
transform 1 0 9292 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _750_
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _751_
timestamp 1666464484
transform -1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _752_
timestamp 1666464484
transform -1 0 11224 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _753_
timestamp 1666464484
transform 1 0 8096 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _754_
timestamp 1666464484
transform -1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _755_
timestamp 1666464484
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _756_
timestamp 1666464484
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _757_
timestamp 1666464484
transform 1 0 19044 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _758_
timestamp 1666464484
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _759_
timestamp 1666464484
transform -1 0 22816 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _760_
timestamp 1666464484
transform 1 0 23368 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _761_
timestamp 1666464484
transform -1 0 23092 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _762_
timestamp 1666464484
transform 1 0 23460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _763_
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _764_
timestamp 1666464484
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _765_
timestamp 1666464484
transform -1 0 6072 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _766_
timestamp 1666464484
transform -1 0 13432 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _767_
timestamp 1666464484
transform 1 0 13524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _768_
timestamp 1666464484
transform 1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _769_
timestamp 1666464484
transform -1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _770_
timestamp 1666464484
transform -1 0 10856 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _771_
timestamp 1666464484
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _772_
timestamp 1666464484
transform -1 0 10396 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _773_
timestamp 1666464484
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _774_
timestamp 1666464484
transform 1 0 12328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _775_
timestamp 1666464484
transform 1 0 4508 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _776_
timestamp 1666464484
transform -1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _777_
timestamp 1666464484
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _778_
timestamp 1666464484
transform -1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _779_
timestamp 1666464484
transform -1 0 4784 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _780_
timestamp 1666464484
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _781_
timestamp 1666464484
transform 1 0 16928 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _782_
timestamp 1666464484
transform -1 0 18952 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _783_
timestamp 1666464484
transform -1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _784_
timestamp 1666464484
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _785_
timestamp 1666464484
transform 1 0 12604 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _786_
timestamp 1666464484
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _787_
timestamp 1666464484
transform -1 0 11960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _788_
timestamp 1666464484
transform -1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _789_
timestamp 1666464484
transform 1 0 12512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _790_
timestamp 1666464484
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _791_
timestamp 1666464484
transform 1 0 16836 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _792_
timestamp 1666464484
transform -1 0 11224 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _793_
timestamp 1666464484
transform 1 0 6532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _794_
timestamp 1666464484
transform -1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _795_
timestamp 1666464484
transform 1 0 6992 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _796_
timestamp 1666464484
transform -1 0 3496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _797_
timestamp 1666464484
transform 1 0 11592 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _798_
timestamp 1666464484
transform -1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _799_
timestamp 1666464484
transform -1 0 11960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _800_
timestamp 1666464484
transform 1 0 11776 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _801_
timestamp 1666464484
transform -1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _802_
timestamp 1666464484
transform 1 0 10764 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _803_
timestamp 1666464484
transform 1 0 10120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _804_
timestamp 1666464484
transform 1 0 10672 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _805_
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _806_
timestamp 1666464484
transform 1 0 11868 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _807_
timestamp 1666464484
transform -1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _808_
timestamp 1666464484
transform 1 0 14260 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _809_
timestamp 1666464484
transform 1 0 14536 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _810_
timestamp 1666464484
transform -1 0 13800 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _811_
timestamp 1666464484
transform 1 0 14260 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _812_
timestamp 1666464484
transform -1 0 13156 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _813_
timestamp 1666464484
transform 1 0 14260 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _814_
timestamp 1666464484
transform -1 0 13800 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _815_
timestamp 1666464484
transform 1 0 16928 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _816_
timestamp 1666464484
transform -1 0 16468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _817_
timestamp 1666464484
transform 1 0 18216 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _818_
timestamp 1666464484
transform -1 0 21344 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _819_
timestamp 1666464484
transform 1 0 20240 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _820_
timestamp 1666464484
transform -1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _821_
timestamp 1666464484
transform 1 0 7360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _822_
timestamp 1666464484
transform 1 0 7360 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _823_
timestamp 1666464484
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _824_
timestamp 1666464484
transform 1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _825_
timestamp 1666464484
transform -1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _826_
timestamp 1666464484
transform -1 0 4508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _827_
timestamp 1666464484
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _828_
timestamp 1666464484
transform -1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _829_
timestamp 1666464484
transform -1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _830_
timestamp 1666464484
transform -1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _831_
timestamp 1666464484
transform -1 0 3036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _832_
timestamp 1666464484
transform -1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _833_
timestamp 1666464484
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _834_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20700 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp 1666464484
transform 1 0 21988 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _836_
timestamp 1666464484
transform 1 0 21988 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp 1666464484
transform 1 0 2576 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _838_
timestamp 1666464484
transform 1 0 2024 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp 1666464484
transform 1 0 3772 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp 1666464484
transform 1 0 2852 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _841_
timestamp 1666464484
transform 1 0 2024 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _842_
timestamp 1666464484
transform 1 0 2024 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _843_
timestamp 1666464484
transform 1 0 1840 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _844_
timestamp 1666464484
transform 1 0 2024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _845_
timestamp 1666464484
transform -1 0 3128 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _846_
timestamp 1666464484
transform 1 0 4416 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _847_
timestamp 1666464484
transform 1 0 4232 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _848_
timestamp 1666464484
transform 1 0 6900 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _849_
timestamp 1666464484
transform 1 0 6348 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _850_
timestamp 1666464484
transform 1 0 2024 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _851_
timestamp 1666464484
transform -1 0 3680 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _852_
timestamp 1666464484
transform 1 0 1932 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _853_
timestamp 1666464484
transform -1 0 3404 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _854_
timestamp 1666464484
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _855_
timestamp 1666464484
transform -1 0 3036 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 3772 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1656 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _858_
timestamp 1666464484
transform 1 0 3956 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _859_
timestamp 1666464484
transform 1 0 3956 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _860_
timestamp 1666464484
transform 1 0 5060 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _861_
timestamp 1666464484
transform 1 0 6532 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _862_
timestamp 1666464484
transform -1 0 3496 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _863_
timestamp 1666464484
transform 1 0 2300 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp 1666464484
transform 1 0 21068 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1666464484
transform -1 0 21528 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp 1666464484
transform -1 0 18952 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp 1666464484
transform 1 0 16192 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp 1666464484
transform 1 0 17480 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp 1666464484
transform 1 0 21988 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp 1666464484
transform 1 0 21988 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp 1666464484
transform 1 0 19320 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp 1666464484
transform 1 0 9844 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11684 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp 1666464484
transform 1 0 9108 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp 1666464484
transform 1 0 8648 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp 1666464484
transform -1 0 8004 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _878_
timestamp 1666464484
transform -1 0 27416 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _879_
timestamp 1666464484
transform 1 0 25484 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _880_
timestamp 1666464484
transform 1 0 25300 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _881_
timestamp 1666464484
transform 1 0 24748 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _882_
timestamp 1666464484
transform 1 0 23920 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _883_
timestamp 1666464484
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _884_
timestamp 1666464484
transform 1 0 14168 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _885_
timestamp 1666464484
transform 1 0 24104 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _886_
timestamp 1666464484
transform 1 0 21528 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _887_
timestamp 1666464484
transform 1 0 18400 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _888_
timestamp 1666464484
transform 1 0 15916 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _889_
timestamp 1666464484
transform -1 0 24472 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _890_
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _891_
timestamp 1666464484
transform -1 0 25576 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _892_
timestamp 1666464484
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _893_
timestamp 1666464484
transform 1 0 14260 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _894_
timestamp 1666464484
transform 1 0 14536 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _895_
timestamp 1666464484
transform 1 0 14812 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _896_
timestamp 1666464484
transform 1 0 16836 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _897_
timestamp 1666464484
transform 1 0 19044 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _898_
timestamp 1666464484
transform 1 0 19412 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _899_
timestamp 1666464484
transform 1 0 20884 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 1666464484
transform -1 0 8648 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1666464484
transform 1 0 9108 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1666464484
transform 1 0 6992 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 1666464484
transform 1 0 5336 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 1666464484
transform -1 0 17020 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 1666464484
transform 1 0 19504 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 1666464484
transform -1 0 20976 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 1666464484
transform -1 0 16100 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 1666464484
transform 1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 1666464484
transform 1 0 15824 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 1666464484
transform -1 0 20884 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 1666464484
transform 1 0 19136 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 1666464484
transform 1 0 17572 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _915_
timestamp 1666464484
transform -1 0 7176 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _916_
timestamp 1666464484
transform 1 0 5612 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _917_
timestamp 1666464484
transform 1 0 6992 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _918_
timestamp 1666464484
transform 1 0 9292 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _919_
timestamp 1666464484
transform 1 0 9108 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _920_
timestamp 1666464484
transform 1 0 11040 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _921_
timestamp 1666464484
transform 1 0 11684 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _922_
timestamp 1666464484
transform -1 0 10580 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _923_
timestamp 1666464484
transform 1 0 8832 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _924_
timestamp 1666464484
transform 1 0 5152 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _925_
timestamp 1666464484
transform 1 0 5520 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 1666464484
transform 1 0 9568 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 1666464484
transform 1 0 19412 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 1666464484
transform -1 0 23000 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 1666464484
transform 1 0 22172 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 1666464484
transform -1 0 10580 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 1666464484
transform 1 0 12144 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _932_
timestamp 1666464484
transform 1 0 12052 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 1666464484
transform -1 0 10580 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 1666464484
transform 1 0 2024 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 1666464484
transform 1 0 2668 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 1666464484
transform 1 0 2576 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _938_
timestamp 1666464484
transform 1 0 17112 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _939_
timestamp 1666464484
transform 1 0 18308 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _940_
timestamp 1666464484
transform 1 0 19412 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _941_
timestamp 1666464484
transform -1 0 21528 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _942_
timestamp 1666464484
transform 1 0 12512 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _943_
timestamp 1666464484
transform -1 0 18676 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _944_
timestamp 1666464484
transform 1 0 11592 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _945_
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _946_
timestamp 1666464484
transform 1 0 13248 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _947_
timestamp 1666464484
transform 1 0 14536 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _948_
timestamp 1666464484
transform -1 0 17480 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _949_
timestamp 1666464484
transform -1 0 11316 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _950_
timestamp 1666464484
transform 1 0 5152 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _951_
timestamp 1666464484
transform 1 0 4600 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _952_
timestamp 1666464484
transform 1 0 11684 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _953_
timestamp 1666464484
transform 1 0 11684 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _954_
timestamp 1666464484
transform 1 0 9752 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _955_
timestamp 1666464484
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _956_
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _957_
timestamp 1666464484
transform 1 0 14260 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _958_
timestamp 1666464484
transform 1 0 13524 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _959_
timestamp 1666464484
transform 1 0 14260 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _960_
timestamp 1666464484
transform 1 0 16836 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _961_
timestamp 1666464484
transform 1 0 21988 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _962_
timestamp 1666464484
transform 1 0 21712 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _963_
timestamp 1666464484
transform 1 0 7360 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _964_
timestamp 1666464484
transform 1 0 7820 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _965_
timestamp 1666464484
transform -1 0 6808 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _966_
timestamp 1666464484
transform -1 0 6072 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _967_
timestamp 1666464484
transform 1 0 5520 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _968_
timestamp 1666464484
transform 1 0 4232 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _969_
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _970_
timestamp 1666464484
transform 1 0 2208 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _971_
timestamp 1666464484
transform -1 0 3496 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _972_
timestamp 1666464484
transform 1 0 1656 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _973_
timestamp 1666464484
transform 1 0 1840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _974_
timestamp 1666464484
transform -1 0 6072 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _975_
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__195_
timestamp 1666464484
transform 1 0 11224 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__212_
timestamp 1666464484
transform 1 0 13156 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__213_
timestamp 1666464484
transform 1 0 16836 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__235_
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__236_
timestamp 1666464484
transform -1 0 10396 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__262_
timestamp 1666464484
transform -1 0 16376 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__263_
timestamp 1666464484
transform 1 0 19688 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__281_
timestamp 1666464484
transform 1 0 15364 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__282_
timestamp 1666464484
transform 1 0 21160 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1666464484
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__195_
timestamp 1666464484
transform -1 0 9660 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__212_
timestamp 1666464484
transform -1 0 13800 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__213_
timestamp 1666464484
transform -1 0 14812 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__235_
timestamp 1666464484
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__236_
timestamp 1666464484
transform -1 0 7084 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__262_
timestamp 1666464484
transform 1 0 12972 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__263_
timestamp 1666464484
transform -1 0 20056 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__281_
timestamp 1666464484
transform -1 0 14812 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__282_
timestamp 1666464484
transform -1 0 20056 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1666464484
transform -1 0 3404 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__195_
timestamp 1666464484
transform 1 0 11960 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__212_
timestamp 1666464484
transform 1 0 12972 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__213_
timestamp 1666464484
transform 1 0 19044 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__235_
timestamp 1666464484
transform -1 0 9660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__236_
timestamp 1666464484
transform 1 0 10396 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__262_
timestamp 1666464484
transform 1 0 12972 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__263_
timestamp 1666464484
transform 1 0 20792 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__281_
timestamp 1666464484
transform 1 0 15640 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__282_
timestamp 1666464484
transform 1 0 24196 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1666464484
transform -1 0 3404 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1666464484
transform -1 0 4968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1666464484
transform -1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1666464484
transform -1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1666464484
transform 1 0 8280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1666464484
transform 1 0 3956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1666464484
transform -1 0 4324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1666464484
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1666464484
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1666464484
transform -1 0 13800 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20148 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 4692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1666464484
transform -1 0 2116 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1666464484
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1666464484
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform 1 0 1564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1666464484
transform 1 0 3496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1666464484
transform 1 0 1564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1666464484
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 2852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform 1 0 4968 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform 1 0 9108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform 1 0 14260 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform 1 0 20148 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform 1 0 26312 0 1 26112
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 io_in[0]
port 1 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[1]
port 2 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 io_in[2]
port 3 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 io_in[3]
port 4 nsew signal input
flabel metal3 s 0 23264 800 23384 0 FreeSans 480 0 0 0 io_in[4]
port 5 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 io_in[5]
port 6 nsew signal input
flabel metal2 s 1858 28200 1914 29000 0 FreeSans 224 90 0 0 io_out[0]
port 7 nsew signal tristate
flabel metal2 s 5446 28200 5502 29000 0 FreeSans 224 90 0 0 io_out[1]
port 8 nsew signal tristate
flabel metal2 s 9034 28200 9090 29000 0 FreeSans 224 90 0 0 io_out[2]
port 9 nsew signal tristate
flabel metal2 s 12622 28200 12678 29000 0 FreeSans 224 90 0 0 io_out[3]
port 10 nsew signal tristate
flabel metal2 s 16210 28200 16266 29000 0 FreeSans 224 90 0 0 io_out[4]
port 11 nsew signal tristate
flabel metal2 s 19798 28200 19854 29000 0 FreeSans 224 90 0 0 io_out[5]
port 12 nsew signal tristate
flabel metal2 s 23386 28200 23442 29000 0 FreeSans 224 90 0 0 io_out[6]
port 13 nsew signal tristate
flabel metal2 s 26974 28200 27030 29000 0 FreeSans 224 90 0 0 io_out[7]
port 14 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 rst
port 15 nsew signal input
flabel metal4 s 4290 2128 4610 26704 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 10982 2128 11302 26704 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 17674 2128 17994 26704 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 24366 2128 24686 26704 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 7636 2128 7956 26704 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 14328 2128 14648 26704 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 21020 2128 21340 26704 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
flabel metal4 s 27712 2128 28032 26704 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 14490 26656 14490 26656 0 vccd1
rlabel via1 14568 26112 14568 26112 0 vssd1
rlabel metal1 3818 2618 3818 2618 0 CIRCUIT_2223.CLK
rlabel metal1 13340 13226 13340 13226 0 CIRCUIT_2223.GATES_1.input1\[0\]
rlabel metal1 15410 14348 15410 14348 0 CIRCUIT_2223.GATES_1.input1\[1\]
rlabel metal1 10810 16150 10810 16150 0 CIRCUIT_2223.GATES_1.input1\[2\]
rlabel metal1 11086 16082 11086 16082 0 CIRCUIT_2223.GATES_1.input1\[3\]
rlabel metal1 2944 12206 2944 12206 0 CIRCUIT_2223.GATES_11.input2
rlabel metal1 9936 19686 9936 19686 0 CIRCUIT_2223.GATES_2.input2
rlabel metal1 10074 19414 10074 19414 0 CIRCUIT_2223.GATES_3.input2
rlabel metal2 5658 24310 5658 24310 0 CIRCUIT_2223.GATES_4.input1\[0\]
rlabel metal1 5704 23290 5704 23290 0 CIRCUIT_2223.GATES_4.input1\[1\]
rlabel metal1 8280 25194 8280 25194 0 CIRCUIT_2223.GATES_4.input1\[2\]
rlabel metal2 8234 23698 8234 23698 0 CIRCUIT_2223.GATES_4.input1\[3\]
rlabel metal1 6072 18938 6072 18938 0 CIRCUIT_2223.GATES_5.input2
rlabel metal1 6256 15130 6256 15130 0 CIRCUIT_2223.MEMORY_18.clock
rlabel metal1 7682 13974 7682 13974 0 CIRCUIT_2223.MEMORY_18.d
rlabel metal1 9108 12138 9108 12138 0 CIRCUIT_2223.MEMORY_18.s_currentState
rlabel metal1 5842 16014 5842 16014 0 CIRCUIT_2223.MEMORY_19.d
rlabel metal1 5428 16218 5428 16218 0 CIRCUIT_2223.MEMORY_19.s_currentState
rlabel metal1 2116 16150 2116 16150 0 CIRCUIT_2223.MEMORY_20.d
rlabel metal2 2254 16388 2254 16388 0 CIRCUIT_2223.MEMORY_20.s_currentState
rlabel metal1 1978 15368 1978 15368 0 CIRCUIT_2223.MEMORY_21.d
rlabel metal1 3312 14994 3312 14994 0 CIRCUIT_2223.MEMORY_21.s_currentState
rlabel metal2 3082 14178 3082 14178 0 CIRCUIT_2223.MEMORY_22.d
rlabel metal2 2162 14110 2162 14110 0 CIRCUIT_2223.MEMORY_22.s_currentState
rlabel metal2 1978 13124 1978 13124 0 CIRCUIT_2223.MEMORY_23.s_currentState
rlabel metal2 6302 13532 6302 13532 0 CIRCUIT_2223.MEMORY_24.d
rlabel metal1 8648 13158 8648 13158 0 CIRCUIT_2223.MEMORY_24.s_currentState
rlabel metal1 5704 14926 5704 14926 0 CIRCUIT_2223.MEMORY_25.d
rlabel metal1 6578 14858 6578 14858 0 CIRCUIT_2223.MEMORY_25.s_currentState
rlabel metal2 7314 15164 7314 15164 0 CIRCUIT_2223.MEMORY_26.s_currentState
rlabel metal1 6486 19754 6486 19754 0 CIRCUIT_2223.s_logisimNet48
rlabel metal2 4002 24582 4002 24582 0 CIRCUIT_2223.tone_generator_1.GATES_1.result
rlabel via1 2249 24174 2249 24174 0 CIRCUIT_2223.tone_generator_1.GATES_2.result
rlabel via1 1881 19822 1881 19822 0 CIRCUIT_2223.tone_generator_1.GATES_3.result
rlabel metal2 2990 19550 2990 19550 0 CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState
rlabel metal2 3358 18870 3358 18870 0 CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState
rlabel metal2 1978 17884 1978 17884 0 CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState
rlabel metal1 3910 17714 3910 17714 0 CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState
rlabel metal1 4922 20366 4922 20366 0 CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState
rlabel metal1 5658 20570 5658 20570 0 CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState
rlabel via1 6877 21114 6877 21114 0 CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState
rlabel metal1 8280 21318 8280 21318 0 CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState
rlabel metal1 2185 21114 2185 21114 0 CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState
rlabel metal1 4462 22066 4462 22066 0 CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState
rlabel via1 4733 23698 4733 23698 0 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState
rlabel metal2 1702 24514 1702 24514 0 CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState
rlabel metal1 4232 24242 4232 24242 0 CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState
rlabel metal1 2392 24922 2392 24922 0 CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState
rlabel metal1 3184 23086 3184 23086 0 CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState
rlabel metal2 2070 22746 2070 22746 0 CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState
rlabel metal1 23644 20774 23644 20774 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2
rlabel metal1 19412 14382 19412 14382 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
rlabel metal2 23414 13328 23414 13328 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2
rlabel metal2 23230 13872 23230 13872 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
rlabel metal1 20746 13328 20746 13328 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
rlabel metal1 23414 15062 23414 15062 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
rlabel metal2 20838 15844 20838 15844 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2
rlabel metal2 17342 16660 17342 16660 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
rlabel metal1 15114 15470 15114 15470 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
rlabel via1 17618 15062 17618 15062 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2
rlabel metal2 20838 19176 20838 19176 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
rlabel metal2 22310 19584 22310 19584 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2
rlabel metal2 27094 18428 27094 18428 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock
rlabel metal1 16238 17544 16238 17544 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d
rlabel metal1 17618 17510 17618 17510 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
rlabel metal1 19688 18190 19688 18190 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d
rlabel metal2 20930 18802 20930 18802 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
rlabel metal1 23782 18836 23782 18836 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d
rlabel metal1 22724 18598 22724 18598 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
rlabel metal2 25438 19482 25438 19482 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d
rlabel metal2 25898 19652 25898 19652 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState
rlabel metal1 14628 16150 14628 16150 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d
rlabel metal2 15962 17238 15962 17238 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
rlabel metal1 24265 16014 24265 16014 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d
rlabel metal1 23644 17646 23644 17646 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
rlabel metal2 24242 17374 24242 17374 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d
rlabel metal1 24242 17646 24242 17646 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState
rlabel metal2 24794 13600 24794 13600 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d
rlabel metal1 24610 13328 24610 13328 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
rlabel metal2 26818 13838 26818 13838 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d
rlabel metal1 24426 15062 24426 15062 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
rlabel metal1 25990 18666 25990 18666 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d
rlabel metal1 24702 15368 24702 15368 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
rlabel metal1 25622 17680 25622 17680 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
rlabel metal2 6762 16966 6762 16966 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d
rlabel metal1 6624 17306 6624 17306 0 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState
rlabel metal1 11960 12138 11960 12138 0 CIRCUIT_2223.tone_generator_2_1.GATES_10.input2
rlabel metal1 8464 11118 8464 11118 0 CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
rlabel metal1 13248 7514 13248 7514 0 CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
rlabel metal1 13662 8806 13662 8806 0 CIRCUIT_2223.tone_generator_2_1.GATES_13.input2
rlabel metal1 9476 9146 9476 9146 0 CIRCUIT_2223.tone_generator_2_1.GATES_14.input2
rlabel metal1 12006 10132 12006 10132 0 CIRCUIT_2223.tone_generator_2_1.GATES_15.input2
rlabel metal2 5014 11492 5014 11492 0 CIRCUIT_2223.tone_generator_2_1.GATES_16.input2
rlabel metal1 5842 11696 5842 11696 0 CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
rlabel metal1 9936 12750 9936 12750 0 CIRCUIT_2223.tone_generator_2_1.GATES_27.result
rlabel metal1 4324 10438 4324 10438 0 CIRCUIT_2223.tone_generator_2_1.GATES_7.input2
rlabel metal1 6854 11730 6854 11730 0 CIRCUIT_2223.tone_generator_2_1.GATES_8.input2
rlabel metal2 6670 11356 6670 11356 0 CIRCUIT_2223.tone_generator_2_1.GATES_9.input2
rlabel metal1 5934 8058 5934 8058 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock
rlabel metal1 6124 6970 6124 6970 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d
rlabel metal2 5382 5916 5382 5916 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState
rlabel metal1 5520 8398 5520 8398 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d
rlabel metal1 5106 8500 5106 8500 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState
rlabel metal2 8050 6052 8050 6052 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d
rlabel metal1 8464 6426 8464 6426 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState
rlabel metal1 11914 6936 11914 6936 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d
rlabel metal1 11500 6630 11500 6630 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState
rlabel metal1 9016 13226 9016 13226 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d
rlabel metal1 10856 12070 10856 12070 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState
rlabel metal2 14030 5984 14030 5984 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d
rlabel metal2 13478 7616 13478 7616 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState
rlabel metal2 12006 5746 12006 5746 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d
rlabel metal1 11316 6290 11316 6290 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState
rlabel metal1 10074 8058 10074 8058 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d
rlabel metal2 8786 8092 8786 8092 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState
rlabel metal1 9936 9486 9936 9486 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d
rlabel metal1 5106 8976 5106 8976 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState
rlabel metal1 5520 10098 5520 10098 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d
rlabel metal1 6118 11118 6118 11118 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState
rlabel metal1 6486 5202 6486 5202 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState
rlabel metal1 9552 18326 9552 18326 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d
rlabel metal1 9568 18734 9568 18734 0 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState
rlabel metal1 19964 21658 19964 21658 0 CIRCUIT_2223.tone_generator_2_2.GATES_10.input2
rlabel metal2 13110 19652 13110 19652 0 CIRCUIT_2223.tone_generator_2_2.GATES_11.input2
rlabel metal1 11178 21420 11178 21420 0 CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
rlabel metal1 11592 23086 11592 23086 0 CIRCUIT_2223.tone_generator_2_2.GATES_13.input2
rlabel metal2 12466 22236 12466 22236 0 CIRCUIT_2223.tone_generator_2_2.GATES_14.input2
rlabel metal1 15134 22746 15134 22746 0 CIRCUIT_2223.tone_generator_2_2.GATES_15.input2
rlabel metal1 15410 21658 15410 21658 0 CIRCUIT_2223.tone_generator_2_2.GATES_16.input2
rlabel metal1 15640 20026 15640 20026 0 CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
rlabel metal2 16146 19958 16146 19958 0 CIRCUIT_2223.tone_generator_2_2.GATES_27.result
rlabel metal1 17480 21658 17480 21658 0 CIRCUIT_2223.tone_generator_2_2.GATES_7.input2
rlabel metal1 17894 19754 17894 19754 0 CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
rlabel metal1 20884 21114 20884 21114 0 CIRCUIT_2223.tone_generator_2_2.GATES_9.input2
rlabel metal2 17618 25024 17618 25024 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock
rlabel metal1 17756 24242 17756 24242 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d
rlabel metal2 18906 23324 18906 23324 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState
rlabel metal2 18630 25262 18630 25262 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d
rlabel metal1 19734 24582 19734 24582 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState
rlabel metal2 20746 25126 20746 25126 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d
rlabel metal1 20976 24174 20976 24174 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState
rlabel metal1 21583 23290 21583 23290 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d
rlabel metal1 20838 22950 20838 22950 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState
rlabel metal1 13340 17102 13340 17102 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d
rlabel metal2 13570 20128 13570 20128 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState
rlabel metal2 18354 21148 18354 21148 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d
rlabel metal1 15548 21114 15548 21114 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState
rlabel metal2 11914 24412 11914 24412 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d
rlabel metal2 12098 25330 12098 25330 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState
rlabel metal2 12466 23936 12466 23936 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d
rlabel metal1 13202 25466 13202 25466 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState
rlabel metal1 14306 24378 14306 24378 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d
rlabel metal1 15042 25840 15042 25840 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState
rlabel metal1 14904 24854 14904 24854 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d
rlabel metal1 15962 24718 15962 24718 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState
rlabel metal1 17618 19822 17618 19822 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState
rlabel metal1 11193 18666 11193 18666 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d
rlabel metal1 10396 19822 10396 19822 0 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState
rlabel metal1 22816 11526 22816 11526 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2
rlabel metal2 14858 10540 14858 10540 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2
rlabel via1 16974 9146 16974 9146 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
rlabel metal1 16100 9690 16100 9690 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
rlabel metal1 18124 12614 18124 12614 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
rlabel metal1 17894 8432 17894 8432 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
rlabel metal2 19458 8602 19458 8602 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2
rlabel metal2 20562 9792 20562 9792 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2
rlabel via2 17526 13243 17526 13243 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result
rlabel metal2 18998 11968 18998 11968 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2
rlabel metal2 22126 10642 22126 10642 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2
rlabel metal1 23184 9894 23184 9894 0 CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2
rlabel metal1 20690 6970 20690 6970 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock
rlabel metal1 25024 7446 25024 7446 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d
rlabel metal1 22632 7514 22632 7514 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState
rlabel metal2 23598 8942 23598 8942 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d
rlabel metal2 23230 9248 23230 9248 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState
rlabel metal2 25254 9792 25254 9792 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d
rlabel metal2 23782 8602 23782 8602 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState
rlabel metal2 24886 11356 24886 11356 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d
rlabel metal2 23230 11968 23230 11968 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState
rlabel metal1 14904 13362 14904 13362 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d
rlabel metal1 15732 11730 15732 11730 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState
rlabel metal2 14858 7582 14858 7582 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d
rlabel metal1 15686 7174 15686 7174 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState
rlabel metal1 16100 6834 16100 6834 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d
rlabel metal2 17250 7854 17250 7854 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState
rlabel metal1 17204 6358 17204 6358 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d
rlabel metal1 19136 13226 19136 13226 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState
rlabel metal2 19366 6494 19366 6494 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d
rlabel metal1 19872 6766 19872 6766 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState
rlabel metal2 19734 6188 19734 6188 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d
rlabel metal1 21298 7378 21298 7378 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState
rlabel metal1 23138 6800 23138 6800 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState
rlabel via1 8330 21998 8330 21998 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d
rlabel metal1 7038 22202 7038 22202 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
rlabel metal1 7038 23834 7038 23834 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock
rlabel via1 9425 24106 9425 24106 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d
rlabel metal2 9614 23868 9614 23868 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
rlabel viali 5653 24106 5653 24106 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock
rlabel metal1 7360 23698 7360 23698 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
rlabel metal1 4830 24854 4830 24854 0 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState
rlabel metal1 2622 18183 2622 18183 0 _000_
rlabel metal2 3082 17476 3082 17476 0 _001_
rlabel metal2 4094 17408 4094 17408 0 _002_
rlabel metal2 4738 20638 4738 20638 0 _003_
rlabel metal1 6532 20570 6532 20570 0 _004_
rlabel metal2 7498 21352 7498 21352 0 _005_
rlabel metal2 2806 20672 2806 20672 0 _006_
rlabel metal2 3450 21080 3450 21080 0 _007_
rlabel metal2 5382 21828 5382 21828 0 _008_
rlabel metal2 26542 17884 26542 17884 0 _009_
rlabel metal2 27370 18190 27370 18190 0 _010_
rlabel metal1 26963 15470 26963 15470 0 _011_
rlabel metal1 25530 15606 25530 15606 0 _012_
rlabel metal2 26634 14076 26634 14076 0 _013_
rlabel metal2 25346 13124 25346 13124 0 _014_
rlabel metal1 26319 13974 26319 13974 0 _015_
rlabel metal1 24564 13838 24564 13838 0 _016_
rlabel metal1 25438 17136 25438 17136 0 _017_
rlabel metal2 23966 17340 23966 17340 0 _018_
rlabel metal2 23322 16626 23322 16626 0 _019_
rlabel metal2 22034 16796 22034 16796 0 _020_
rlabel metal2 15778 16626 15778 16626 0 _021_
rlabel metal1 25576 18802 25576 18802 0 _022_
rlabel metal1 23920 19346 23920 19346 0 _023_
rlabel metal2 22862 18496 22862 18496 0 _024_
rlabel metal2 21574 18972 21574 18972 0 _025_
rlabel metal2 19366 17782 19366 17782 0 _026_
rlabel metal2 18446 18428 18446 18428 0 _027_
rlabel metal1 17533 17578 17533 17578 0 _028_
rlabel metal1 16468 17714 16468 17714 0 _029_
rlabel metal1 22901 7446 22901 7446 0 _030_
rlabel metal1 23460 6834 23460 6834 0 _031_
rlabel metal1 24748 7922 24748 7922 0 _032_
rlabel metal1 23644 8398 23644 8398 0 _033_
rlabel metal1 24748 9010 24748 9010 0 _034_
rlabel metal2 25530 9044 25530 9044 0 _035_
rlabel metal2 24978 10914 24978 10914 0 _036_
rlabel metal2 24794 10642 24794 10642 0 _037_
rlabel metal2 15318 12750 15318 12750 0 _038_
rlabel metal2 15962 6902 15962 6902 0 _039_
rlabel metal1 14950 7310 14950 7310 0 _040_
rlabel metal2 16146 6222 16146 6222 0 _041_
rlabel metal2 13754 6290 13754 6290 0 _042_
rlabel metal1 17664 5746 17664 5746 0 _043_
rlabel metal2 16882 5746 16882 5746 0 _044_
rlabel metal2 19642 5236 19642 5236 0 _045_
rlabel metal2 18446 6052 18446 6052 0 _046_
rlabel metal1 20608 7310 20608 7310 0 _047_
rlabel metal1 19136 5746 19136 5746 0 _048_
rlabel metal1 22356 8806 22356 8806 0 _049_
rlabel metal2 20930 7004 20930 7004 0 _050_
rlabel metal1 7958 23834 7958 23834 0 _051_
rlabel metal2 7038 25228 7038 25228 0 _052_
rlabel metal2 5382 25262 5382 25262 0 _053_
rlabel metal1 6493 6698 6493 6698 0 _054_
rlabel metal2 7222 6052 7222 6052 0 _055_
rlabel metal2 6026 5916 6026 5916 0 _056_
rlabel metal2 5658 5508 5658 5508 0 _057_
rlabel metal2 8326 5848 8326 5848 0 _058_
rlabel metal1 6992 6290 6992 6290 0 _059_
rlabel metal2 10626 6222 10626 6222 0 _060_
rlabel metal2 9154 6018 9154 6018 0 _061_
rlabel metal2 10442 12002 10442 12002 0 _062_
rlabel metal1 11500 5338 11500 5338 0 _063_
rlabel metal1 11224 5746 11224 5746 0 _064_
rlabel metal2 12650 6494 12650 6494 0 _065_
rlabel metal1 11684 6290 11684 6290 0 _066_
rlabel metal1 9292 6426 9292 6426 0 _067_
rlabel metal1 10718 6358 10718 6358 0 _068_
rlabel metal2 10258 9724 10258 9724 0 _069_
rlabel metal1 8648 9486 8648 9486 0 _070_
rlabel metal2 6578 9826 6578 9826 0 _071_
rlabel metal1 5152 9146 5152 9146 0 _072_
rlabel metal2 6578 8738 6578 8738 0 _073_
rlabel metal2 5566 8772 5566 8772 0 _074_
rlabel metal2 18538 23664 18538 23664 0 _075_
rlabel metal2 17158 24956 17158 24956 0 _076_
rlabel metal2 19734 24446 19734 24446 0 _077_
rlabel metal2 18354 24990 18354 24990 0 _078_
rlabel metal1 20746 25806 20746 25806 0 _079_
rlabel metal2 19458 25806 19458 25806 0 _080_
rlabel metal1 20792 22678 20792 22678 0 _081_
rlabel metal2 21482 23630 21482 23630 0 _082_
rlabel metal2 13478 17408 13478 17408 0 _083_
rlabel metal2 17342 20672 17342 20672 0 _084_
rlabel metal2 13662 20128 13662 20128 0 _085_
rlabel metal2 13202 23630 13202 23630 0 _086_
rlabel metal1 11730 22746 11730 22746 0 _087_
rlabel metal2 13294 25772 13294 25772 0 _088_
rlabel metal2 11914 25500 11914 25500 0 _089_
rlabel metal2 14122 25364 14122 25364 0 _090_
rlabel metal1 13064 25806 13064 25806 0 _091_
rlabel metal2 16146 25568 16146 25568 0 _092_
rlabel metal1 15042 24718 15042 24718 0 _093_
rlabel metal2 16606 24718 16606 24718 0 _094_
rlabel metal1 17296 24854 17296 24854 0 _095_
rlabel metal1 21344 21862 21344 21862 0 _096_
rlabel metal1 21482 20298 21482 20298 0 _097_
rlabel metal1 7912 17850 7912 17850 0 _098_
rlabel metal1 8089 19414 8089 19414 0 _099_
rlabel metal1 4823 18666 4823 18666 0 _100_
rlabel metal2 4646 17782 4646 17782 0 _101_
rlabel metal1 5474 15334 5474 15334 0 _102_
rlabel metal1 5612 14586 5612 14586 0 _103_
rlabel metal2 5014 14824 5014 14824 0 _104_
rlabel metal1 4232 14586 4232 14586 0 _105_
rlabel metal1 6026 13838 6026 13838 0 _106_
rlabel metal1 4278 13838 4278 13838 0 _107_
rlabel metal2 2254 12988 2254 12988 0 _108_
rlabel metal1 1794 12954 1794 12954 0 _109_
rlabel metal2 2254 14144 2254 14144 0 _110_
rlabel metal1 3542 14042 3542 14042 0 _111_
rlabel metal2 1702 15266 1702 15266 0 _112_
rlabel metal2 3726 15640 3726 15640 0 _113_
rlabel metal2 2806 16218 2806 16218 0 _114_
rlabel metal1 5527 16150 5527 16150 0 _115_
rlabel metal2 6026 16252 6026 16252 0 _116_
rlabel metal1 15410 13906 15410 13906 0 _117_
rlabel metal2 7498 14348 7498 14348 0 _118_
rlabel via1 21017 10030 21017 10030 0 _119_
rlabel metal1 20470 10744 20470 10744 0 _120_
rlabel metal2 21942 11934 21942 11934 0 _121_
rlabel metal2 2898 4556 2898 4556 0 _122_
rlabel via1 2341 3434 2341 3434 0 _123_
rlabel metal1 4135 3094 4135 3094 0 _124_
rlabel metal1 3066 4182 3066 4182 0 _125_
rlabel metal1 2944 5882 2944 5882 0 _126_
rlabel metal2 5290 6970 5290 6970 0 _127_
rlabel metal2 2714 8738 2714 8738 0 _128_
rlabel metal1 2433 9622 2433 9622 0 _129_
rlabel metal1 21344 12954 21344 12954 0 _130_
rlabel metal2 22954 16422 22954 16422 0 _131_
rlabel metal1 19059 15062 19059 15062 0 _132_
rlabel metal1 16693 14382 16693 14382 0 _133_
rlabel metal1 18395 13974 18395 13974 0 _134_
rlabel metal1 22179 13974 22179 13974 0 _135_
rlabel metal1 23087 13226 23087 13226 0 _136_
rlabel metal1 19596 12954 19596 12954 0 _137_
rlabel metal1 10064 14382 10064 14382 0 _138_
rlabel metal1 11904 14382 11904 14382 0 _139_
rlabel metal1 9236 14994 9236 14994 0 _140_
rlabel metal1 8586 16150 8586 16150 0 _141_
rlabel metal1 16800 18734 16800 18734 0 _142_
rlabel metal1 19724 20910 19724 20910 0 _143_
rlabel metal1 21344 21114 21344 21114 0 _144_
rlabel metal1 15880 11118 15880 11118 0 _145_
rlabel metal1 15118 8874 15118 8874 0 _146_
rlabel metal2 15962 9078 15962 9078 0 _147_
rlabel metal1 16100 11866 16100 11866 0 _148_
rlabel metal1 17326 9962 17326 9962 0 _149_
rlabel metal1 20664 8942 20664 8942 0 _150_
rlabel via1 19453 9554 19453 9554 0 _151_
rlabel metal1 17756 11322 17756 11322 0 _152_
rlabel metal1 19304 18666 19304 18666 0 _153_
rlabel metal1 23061 19754 23061 19754 0 _154_
rlabel metal2 23506 20706 23506 20706 0 _155_
rlabel metal1 9342 13294 9342 13294 0 _156_
rlabel metal1 13013 7378 13013 7378 0 _157_
rlabel metal1 12272 8942 12272 8942 0 _158_
rlabel metal2 10994 8738 10994 8738 0 _159_
rlabel metal2 12466 10880 12466 10880 0 _160_
rlabel metal2 2162 10914 2162 10914 0 _161_
rlabel metal1 2859 11798 2859 11798 0 _162_
rlabel metal1 3859 10710 3859 10710 0 _163_
rlabel via1 5469 12138 5469 12138 0 _164_
rlabel metal1 4538 12886 4538 12886 0 _165_
rlabel metal1 11960 10778 11960 10778 0 _166_
rlabel metal1 11270 17850 11270 17850 0 _167_
rlabel metal1 10120 21114 10120 21114 0 _168_
rlabel via1 10069 22678 10069 22678 0 _169_
rlabel metal1 9614 21896 9614 21896 0 _170_
rlabel metal1 14480 21998 14480 21998 0 _171_
rlabel metal2 13110 21318 13110 21318 0 _172_
rlabel metal1 14336 19754 14336 19754 0 _173_
rlabel metal1 16422 21896 16422 21896 0 _174_
rlabel metal1 7544 18326 7544 18326 0 _175_
rlabel metal1 8648 19278 8648 19278 0 _176_
rlabel metal2 6578 18530 6578 18530 0 _177_
rlabel metal2 5750 18734 5750 18734 0 _178_
rlabel metal2 1794 13294 1794 13294 0 _179_
rlabel metal2 13110 17544 13110 17544 0 _180_
rlabel metal1 14168 17578 14168 17578 0 _181_
rlabel metal1 11086 19278 11086 19278 0 _182_
rlabel metal2 5290 19652 5290 19652 0 _183_
rlabel metal1 22448 20434 22448 20434 0 _184_
rlabel metal2 6762 18700 6762 18700 0 _185_
rlabel metal2 23598 18870 23598 18870 0 _186_
rlabel metal1 10028 19482 10028 19482 0 _187_
rlabel metal1 22540 14994 22540 14994 0 _188_
rlabel metal1 7544 18734 7544 18734 0 _189_
rlabel metal1 5566 7786 5566 7786 0 _190_
rlabel metal1 22908 6290 22908 6290 0 _191_
rlabel metal2 12650 16898 12650 16898 0 _192_
rlabel metal1 18722 17578 18722 17578 0 _193_
rlabel metal1 13202 18258 13202 18258 0 _194_
rlabel metal1 5290 12172 5290 12172 0 _195_
rlabel metal1 12788 21454 12788 21454 0 _196_
rlabel metal1 13938 23494 13938 23494 0 _197_
rlabel metal1 15272 23154 15272 23154 0 _198_
rlabel metal1 20102 22032 20102 22032 0 _199_
rlabel metal2 15870 21148 15870 21148 0 _200_
rlabel metal1 16100 20026 16100 20026 0 _201_
rlabel metal1 17756 20026 17756 20026 0 _202_
rlabel metal2 16974 20264 16974 20264 0 _203_
rlabel metal1 15852 20434 15852 20434 0 _204_
rlabel metal1 14766 20298 14766 20298 0 _205_
rlabel metal1 16192 20570 16192 20570 0 _206_
rlabel metal2 17250 22814 17250 22814 0 _207_
rlabel metal2 18722 22882 18722 22882 0 _208_
rlabel metal1 13984 22542 13984 22542 0 _209_
rlabel metal2 16330 22780 16330 22780 0 _210_
rlabel metal1 16606 20910 16606 20910 0 _211_
rlabel metal1 12604 18326 12604 18326 0 _212_
rlabel metal1 14720 19482 14720 19482 0 _213_
rlabel metal1 22494 17068 22494 17068 0 _214_
rlabel metal1 25438 18190 25438 18190 0 _215_
rlabel metal2 13110 8432 13110 8432 0 _216_
rlabel metal2 12834 9690 12834 9690 0 _217_
rlabel metal1 12650 10098 12650 10098 0 _218_
rlabel metal1 14260 8058 14260 8058 0 _219_
rlabel metal1 10925 11050 10925 11050 0 _220_
rlabel metal1 7544 11322 7544 11322 0 _221_
rlabel viali 8144 11730 8144 11730 0 _222_
rlabel metal1 7958 11696 7958 11696 0 _223_
rlabel viali 7774 11730 7774 11730 0 _224_
rlabel metal1 7130 11696 7130 11696 0 _225_
rlabel metal2 9246 11390 9246 11390 0 _226_
rlabel metal2 7682 10234 7682 10234 0 _227_
rlabel metal2 5566 10336 5566 10336 0 _228_
rlabel metal2 7498 9758 7498 9758 0 _229_
rlabel metal1 7728 9146 7728 9146 0 _230_
rlabel metal1 8510 10234 8510 10234 0 _231_
rlabel metal1 9890 14314 9890 14314 0 _232_
rlabel metal1 10948 11730 10948 11730 0 _233_
rlabel metal1 11224 12750 11224 12750 0 _234_
rlabel metal1 10212 11118 10212 11118 0 _235_
rlabel metal2 13018 8942 13018 8942 0 _236_
rlabel metal1 5382 6324 5382 6324 0 _237_
rlabel metal2 18538 13022 18538 13022 0 _238_
rlabel metal1 18489 12818 18489 12818 0 _239_
rlabel metal1 19182 12886 19182 12886 0 _240_
rlabel via1 18740 12818 18740 12818 0 _241_
rlabel metal1 22678 12410 22678 12410 0 _242_
rlabel metal1 17618 13328 17618 13328 0 _243_
rlabel metal2 18262 8058 18262 8058 0 _244_
rlabel metal2 18446 7684 18446 7684 0 _245_
rlabel metal1 17664 7514 17664 7514 0 _246_
rlabel metal1 17664 7854 17664 7854 0 _247_
rlabel metal1 18584 8058 18584 8058 0 _248_
rlabel metal1 20010 9146 20010 9146 0 _249_
rlabel metal1 20378 8330 20378 8330 0 _250_
rlabel metal2 23046 8840 23046 8840 0 _251_
rlabel metal2 22862 9282 22862 9282 0 _252_
rlabel metal2 18354 9860 18354 9860 0 _253_
rlabel metal2 17618 9350 17618 9350 0 _254_
rlabel metal2 18906 9146 18906 9146 0 _255_
rlabel metal2 17434 13532 17434 13532 0 _256_
rlabel metal1 15364 12954 15364 12954 0 _257_
rlabel metal1 14766 11798 14766 11798 0 _258_
rlabel metal1 14904 13770 14904 13770 0 _259_
rlabel metal1 13202 13396 13202 13396 0 _260_
rlabel via2 12466 13515 12466 13515 0 _261_
rlabel metal1 16100 12886 16100 12886 0 _262_
rlabel metal2 19734 10064 19734 10064 0 _263_
rlabel metal1 24242 15470 24242 15470 0 _264_
rlabel metal1 25024 20026 25024 20026 0 _265_
rlabel metal1 24840 14926 24840 14926 0 _266_
rlabel metal1 24426 14858 24426 14858 0 _267_
rlabel metal1 23368 15606 23368 15606 0 _268_
rlabel metal1 20240 17238 20240 17238 0 _269_
rlabel via1 20564 17170 20564 17170 0 _270_
rlabel metal1 19964 14586 19964 14586 0 _271_
rlabel metal1 19964 15130 19964 15130 0 _272_
rlabel metal1 18354 17102 18354 17102 0 _273_
rlabel metal1 21252 17034 21252 17034 0 _274_
rlabel metal1 22885 16558 22885 16558 0 _275_
rlabel metal2 22494 17238 22494 17238 0 _276_
rlabel metal1 22954 13464 22954 13464 0 _277_
rlabel metal1 22954 15674 22954 15674 0 _278_
rlabel metal1 23460 16422 23460 16422 0 _279_
rlabel metal1 14306 15402 14306 15402 0 _280_
rlabel metal2 15410 16082 15410 16082 0 _281_
rlabel metal1 21160 16558 21160 16558 0 _282_
rlabel metal1 5060 25874 5060 25874 0 _283_
rlabel metal1 6256 25262 6256 25262 0 _284_
rlabel metal2 6394 24752 6394 24752 0 _285_
rlabel metal1 5658 25806 5658 25806 0 _286_
rlabel metal1 10166 24854 10166 24854 0 _287_
rlabel metal1 8924 25330 8924 25330 0 _288_
rlabel metal1 8326 25772 8326 25772 0 _289_
rlabel metal2 7406 25602 7406 25602 0 _290_
rlabel metal1 10350 24650 10350 24650 0 _291_
rlabel metal1 9752 24650 9752 24650 0 _292_
rlabel metal1 9844 24922 9844 24922 0 _293_
rlabel metal1 8464 25398 8464 25398 0 _294_
rlabel metal2 9890 26010 9890 26010 0 _295_
rlabel metal1 9982 20434 9982 20434 0 _296_
rlabel metal1 10810 24174 10810 24174 0 _297_
rlabel metal2 10718 24752 10718 24752 0 _298_
rlabel metal1 10166 25262 10166 25262 0 _299_
rlabel metal1 4462 25840 4462 25840 0 _300_
rlabel metal1 20562 12818 20562 12818 0 _301_
rlabel metal1 22770 11186 22770 11186 0 _302_
rlabel metal1 21252 10642 21252 10642 0 _303_
rlabel metal2 20286 10438 20286 10438 0 _304_
rlabel metal2 21758 11764 21758 11764 0 _305_
rlabel metal1 6670 3706 6670 3706 0 _306_
rlabel metal2 2806 5236 2806 5236 0 _307_
rlabel metal1 4600 5066 4600 5066 0 _308_
rlabel metal1 4738 5202 4738 5202 0 _309_
rlabel metal1 3450 5678 3450 5678 0 _310_
rlabel metal1 3174 4624 3174 4624 0 _311_
rlabel metal1 4232 6086 4232 6086 0 _312_
rlabel metal2 3174 5508 3174 5508 0 _313_
rlabel metal1 4370 6664 4370 6664 0 _314_
rlabel metal2 5658 7854 5658 7854 0 _315_
rlabel metal1 4738 5678 4738 5678 0 _316_
rlabel metal1 4784 5882 4784 5882 0 _317_
rlabel metal1 2070 8330 2070 8330 0 _318_
rlabel metal1 2714 20468 2714 20468 0 _319_
rlabel metal1 7544 19822 7544 19822 0 _320_
rlabel metal1 20654 15980 20654 15980 0 _321_
rlabel metal2 21482 13804 21482 13804 0 _322_
rlabel metal1 22724 17646 22724 17646 0 _323_
rlabel metal2 19642 15674 19642 15674 0 _324_
rlabel metal1 16698 14994 16698 14994 0 _325_
rlabel metal1 11178 11764 11178 11764 0 _326_
rlabel metal2 18354 13974 18354 13974 0 _327_
rlabel metal1 20286 14416 20286 14416 0 _328_
rlabel metal1 21988 12954 21988 12954 0 _329_
rlabel metal2 24058 13770 24058 13770 0 _330_
rlabel metal2 19366 12988 19366 12988 0 _331_
rlabel metal1 9660 15334 9660 15334 0 _332_
rlabel metal1 8464 14382 8464 14382 0 _333_
rlabel metal1 10948 14994 10948 14994 0 _334_
rlabel metal1 7406 16048 7406 16048 0 _335_
rlabel metal2 8050 16252 8050 16252 0 _336_
rlabel metal1 15548 19278 15548 19278 0 _337_
rlabel metal1 16698 19346 16698 19346 0 _338_
rlabel metal2 19826 20774 19826 20774 0 _339_
rlabel metal1 21068 20570 21068 20570 0 _340_
rlabel metal1 16284 10778 16284 10778 0 _341_
rlabel metal2 14582 9146 14582 9146 0 _342_
rlabel metal2 16146 9180 16146 9180 0 _343_
rlabel metal1 16790 12614 16790 12614 0 _344_
rlabel metal1 19550 12614 19550 12614 0 _345_
rlabel metal2 16790 10268 16790 10268 0 _346_
rlabel metal1 19550 8602 19550 8602 0 _347_
rlabel metal1 19504 10234 19504 10234 0 _348_
rlabel metal2 18078 11594 18078 11594 0 _349_
rlabel metal1 22264 20366 22264 20366 0 _350_
rlabel metal2 18722 18938 18722 18938 0 _351_
rlabel metal1 23184 19482 23184 19482 0 _352_
rlabel metal1 23368 20434 23368 20434 0 _353_
rlabel metal2 10166 10132 10166 10132 0 _354_
rlabel metal1 7636 11254 7636 11254 0 _355_
rlabel metal1 13570 8058 13570 8058 0 _356_
rlabel metal1 12052 9554 12052 9554 0 _357_
rlabel metal1 11270 8466 11270 8466 0 _358_
rlabel metal1 5244 11662 5244 11662 0 _359_
rlabel metal2 12558 11356 12558 11356 0 _360_
rlabel metal2 4186 11084 4186 11084 0 _361_
rlabel metal2 4002 11900 4002 11900 0 _362_
rlabel metal1 6486 11152 6486 11152 0 _363_
rlabel metal1 9706 11594 9706 11594 0 _364_
rlabel metal1 5658 12954 5658 12954 0 _365_
rlabel metal1 7084 12410 7084 12410 0 _366_
rlabel metal2 11730 11356 11730 11356 0 _367_
rlabel metal1 12466 22100 12466 22100 0 _368_
rlabel metal2 10534 18666 10534 18666 0 _369_
rlabel metal1 10580 20910 10580 20910 0 _370_
rlabel metal1 10488 23086 10488 23086 0 _371_
rlabel metal1 11914 21930 11914 21930 0 _372_
rlabel metal2 14950 21182 14950 21182 0 _373_
rlabel metal1 13708 21998 13708 21998 0 _374_
rlabel metal1 12926 20944 12926 20944 0 _375_
rlabel metal1 14260 20570 14260 20570 0 _376_
rlabel metal1 16606 21658 16606 21658 0 _377_
rlabel metal1 18676 19482 18676 19482 0 _378_
rlabel metal2 20654 19958 20654 19958 0 _379_
rlabel metal2 3266 2193 3266 2193 0 clk
rlabel metal1 11914 15402 11914 15402 0 clknet_0__195_
rlabel metal1 14352 18394 14352 18394 0 clknet_0__212_
rlabel metal1 18170 23800 18170 23800 0 clknet_0__213_
rlabel metal1 10488 10710 10488 10710 0 clknet_0__235_
rlabel metal1 9384 4590 9384 4590 0 clknet_0__236_
rlabel metal3 13754 12580 13754 12580 0 clknet_0__262_
rlabel metal2 20838 6528 20838 6528 0 clknet_0__263_
rlabel metal2 15686 15946 15686 15946 0 clknet_0__281_
rlabel metal1 22448 16422 22448 16422 0 clknet_0__282_
rlabel metal2 3358 7650 3358 7650 0 clknet_0_clk
rlabel metal1 6578 12886 6578 12886 0 clknet_1_0__leaf__195_
rlabel metal1 12650 16218 12650 16218 0 clknet_1_0__leaf__212_
rlabel metal2 15778 25262 15778 25262 0 clknet_1_0__leaf__213_
rlabel metal2 12190 9248 12190 9248 0 clknet_1_0__leaf__235_
rlabel metal2 5566 5508 5566 5508 0 clknet_1_0__leaf__236_
rlabel metal1 15824 8534 15824 8534 0 clknet_1_0__leaf__262_
rlabel metal1 18814 5338 18814 5338 0 clknet_1_0__leaf__263_
rlabel metal1 14352 15130 14352 15130 0 clknet_1_0__leaf__281_
rlabel metal2 22402 17714 22402 17714 0 clknet_1_0__leaf__282_
rlabel metal2 2070 6528 2070 6528 0 clknet_1_0__leaf_clk
rlabel metal1 12926 15674 12926 15674 0 clknet_1_1__leaf__195_
rlabel metal1 12374 19278 12374 19278 0 clknet_1_1__leaf__212_
rlabel metal2 19918 25024 19918 25024 0 clknet_1_1__leaf__213_
rlabel metal1 9016 10778 9016 10778 0 clknet_1_1__leaf__235_
rlabel metal2 10810 4998 10810 4998 0 clknet_1_1__leaf__236_
rlabel metal2 14766 13056 14766 13056 0 clknet_1_1__leaf__262_
rlabel metal1 24518 6290 24518 6290 0 clknet_1_1__leaf__263_
rlabel metal2 16882 16422 16882 16422 0 clknet_1_1__leaf__281_
rlabel metal1 25523 18258 25523 18258 0 clknet_1_1__leaf__282_
rlabel metal1 3266 12172 3266 12172 0 clknet_1_1__leaf_clk
rlabel metal1 2668 2618 2668 2618 0 io_in[0]
rlabel metal3 1142 12716 1142 12716 0 io_in[1]
rlabel metal2 1610 19244 1610 19244 0 io_in[2]
rlabel metal2 1702 20111 1702 20111 0 io_in[3]
rlabel metal2 3542 23511 3542 23511 0 io_in[4]
rlabel metal3 1188 26860 1188 26860 0 io_in[5]
rlabel metal1 2254 26554 2254 26554 0 io_out[0]
rlabel metal1 5336 26554 5336 26554 0 io_out[1]
rlabel metal1 9200 26554 9200 26554 0 io_out[2]
rlabel metal1 13570 26214 13570 26214 0 io_out[3]
rlabel metal1 16652 26214 16652 26214 0 io_out[4]
rlabel metal1 20102 26554 20102 26554 0 io_out[5]
rlabel metal1 23598 26554 23598 26554 0 io_out[6]
rlabel metal1 26772 26554 26772 26554 0 io_out[7]
rlabel metal2 1702 14620 1702 14620 0 net1
rlabel metal1 8924 26010 8924 26010 0 net10
rlabel metal2 13846 26146 13846 26146 0 net11
rlabel metal1 14582 25704 14582 25704 0 net12
rlabel metal1 16146 25398 16146 25398 0 net13
rlabel metal1 23322 21862 23322 21862 0 net14
rlabel metal1 24886 21658 24886 21658 0 net15
rlabel metal1 1932 21454 1932 21454 0 net16
rlabel metal1 1702 17782 1702 17782 0 net17
rlabel metal2 5198 11764 5198 11764 0 net18
rlabel metal2 12098 8160 12098 8160 0 net19
rlabel metal1 6118 12376 6118 12376 0 net2
rlabel metal2 10442 14586 10442 14586 0 net20
rlabel metal1 4186 2550 4186 2550 0 net21
rlabel metal1 21022 14382 21022 14382 0 net22
rlabel metal1 17572 13906 17572 13906 0 net23
rlabel metal1 16284 14382 16284 14382 0 net24
rlabel metal2 21482 15232 21482 15232 0 net25
rlabel metal1 6026 13396 6026 13396 0 net26
rlabel metal1 13248 12954 13248 12954 0 net27
rlabel metal2 4186 9758 4186 9758 0 net28
rlabel metal1 1748 14042 1748 14042 0 net3
rlabel metal2 4830 5168 4830 5168 0 net4
rlabel metal1 5428 3706 5428 3706 0 net5
rlabel metal1 4738 11118 4738 11118 0 net6
rlabel metal1 2208 5678 2208 5678 0 net7
rlabel metal2 4554 26180 4554 26180 0 net8
rlabel metal1 5060 26010 5060 26010 0 net9
rlabel metal2 2806 3502 2806 3502 0 rst
rlabel metal1 2806 4556 2806 4556 0 slow_clock\[0\]
rlabel metal2 3450 4216 3450 4216 0 slow_clock\[1\]
rlabel via1 5190 4182 5190 4182 0 slow_clock\[2\]
rlabel metal1 3818 4590 3818 4590 0 slow_clock\[3\]
rlabel metal2 4002 6494 4002 6494 0 slow_clock\[4\]
rlabel metal1 3818 6834 3818 6834 0 slow_clock\[5\]
rlabel metal1 3266 9044 3266 9044 0 slow_clock\[6\]
<< properties >>
string FIXED_BBOX 0 0 29000 29000
<< end >>
